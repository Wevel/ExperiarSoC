magic
tech sky130A
magscale 1 2
timestamp 1683759936
<< obsli1 >>
rect 1104 2159 118864 187697
<< obsm1 >>
rect 934 892 119126 189100
<< metal2 >>
rect 1306 189200 1362 190000
rect 2870 189200 2926 190000
rect 4434 189200 4490 190000
rect 5998 189200 6054 190000
rect 7562 189200 7618 190000
rect 9126 189200 9182 190000
rect 10690 189200 10746 190000
rect 12254 189200 12310 190000
rect 13818 189200 13874 190000
rect 15382 189200 15438 190000
rect 16946 189200 17002 190000
rect 18510 189200 18566 190000
rect 20074 189200 20130 190000
rect 21638 189200 21694 190000
rect 23202 189200 23258 190000
rect 24766 189200 24822 190000
rect 26330 189200 26386 190000
rect 27894 189200 27950 190000
rect 29458 189200 29514 190000
rect 31022 189200 31078 190000
rect 32586 189200 32642 190000
rect 34150 189200 34206 190000
rect 35714 189200 35770 190000
rect 37278 189200 37334 190000
rect 38842 189200 38898 190000
rect 40406 189200 40462 190000
rect 41970 189200 42026 190000
rect 43534 189200 43590 190000
rect 45098 189200 45154 190000
rect 46662 189200 46718 190000
rect 48226 189200 48282 190000
rect 49790 189200 49846 190000
rect 51354 189200 51410 190000
rect 52918 189200 52974 190000
rect 54482 189200 54538 190000
rect 56046 189200 56102 190000
rect 57610 189200 57666 190000
rect 59174 189200 59230 190000
rect 60738 189200 60794 190000
rect 62302 189200 62358 190000
rect 63866 189200 63922 190000
rect 65430 189200 65486 190000
rect 66994 189200 67050 190000
rect 68558 189200 68614 190000
rect 70122 189200 70178 190000
rect 71686 189200 71742 190000
rect 73250 189200 73306 190000
rect 74814 189200 74870 190000
rect 76378 189200 76434 190000
rect 77942 189200 77998 190000
rect 79506 189200 79562 190000
rect 81070 189200 81126 190000
rect 82634 189200 82690 190000
rect 84198 189200 84254 190000
rect 85762 189200 85818 190000
rect 87326 189200 87382 190000
rect 88890 189200 88946 190000
rect 90454 189200 90510 190000
rect 92018 189200 92074 190000
rect 93582 189200 93638 190000
rect 95146 189200 95202 190000
rect 96710 189200 96766 190000
rect 98274 189200 98330 190000
rect 99838 189200 99894 190000
rect 101402 189200 101458 190000
rect 102966 189200 103022 190000
rect 104530 189200 104586 190000
rect 106094 189200 106150 190000
rect 107658 189200 107714 190000
rect 109222 189200 109278 190000
rect 110786 189200 110842 190000
rect 112350 189200 112406 190000
rect 113914 189200 113970 190000
rect 115478 189200 115534 190000
rect 117042 189200 117098 190000
rect 118606 189200 118662 190000
rect 3146 0 3202 800
rect 4894 0 4950 800
rect 6642 0 6698 800
rect 8390 0 8446 800
rect 10138 0 10194 800
rect 11886 0 11942 800
rect 13634 0 13690 800
rect 15382 0 15438 800
rect 17130 0 17186 800
rect 18878 0 18934 800
rect 20626 0 20682 800
rect 22374 0 22430 800
rect 24122 0 24178 800
rect 25870 0 25926 800
rect 27618 0 27674 800
rect 29366 0 29422 800
rect 31114 0 31170 800
rect 32862 0 32918 800
rect 34610 0 34666 800
rect 36358 0 36414 800
rect 38106 0 38162 800
rect 39854 0 39910 800
rect 41602 0 41658 800
rect 43350 0 43406 800
rect 45098 0 45154 800
rect 46846 0 46902 800
rect 48594 0 48650 800
rect 50342 0 50398 800
rect 52090 0 52146 800
rect 53838 0 53894 800
rect 55586 0 55642 800
rect 57334 0 57390 800
rect 59082 0 59138 800
rect 60830 0 60886 800
rect 62578 0 62634 800
rect 64326 0 64382 800
rect 66074 0 66130 800
rect 67822 0 67878 800
rect 69570 0 69626 800
rect 71318 0 71374 800
rect 73066 0 73122 800
rect 74814 0 74870 800
rect 76562 0 76618 800
rect 78310 0 78366 800
rect 80058 0 80114 800
rect 81806 0 81862 800
rect 83554 0 83610 800
rect 85302 0 85358 800
rect 87050 0 87106 800
rect 88798 0 88854 800
rect 90546 0 90602 800
rect 92294 0 92350 800
rect 94042 0 94098 800
rect 95790 0 95846 800
rect 97538 0 97594 800
rect 99286 0 99342 800
rect 101034 0 101090 800
rect 102782 0 102838 800
rect 104530 0 104586 800
rect 106278 0 106334 800
rect 108026 0 108082 800
rect 109774 0 109830 800
rect 111522 0 111578 800
rect 113270 0 113326 800
rect 115018 0 115074 800
rect 116766 0 116822 800
<< obsm2 >>
rect 938 189144 1250 189200
rect 1418 189144 2814 189200
rect 2982 189144 4378 189200
rect 4546 189144 5942 189200
rect 6110 189144 7506 189200
rect 7674 189144 9070 189200
rect 9238 189144 10634 189200
rect 10802 189144 12198 189200
rect 12366 189144 13762 189200
rect 13930 189144 15326 189200
rect 15494 189144 16890 189200
rect 17058 189144 18454 189200
rect 18622 189144 20018 189200
rect 20186 189144 21582 189200
rect 21750 189144 23146 189200
rect 23314 189144 24710 189200
rect 24878 189144 26274 189200
rect 26442 189144 27838 189200
rect 28006 189144 29402 189200
rect 29570 189144 30966 189200
rect 31134 189144 32530 189200
rect 32698 189144 34094 189200
rect 34262 189144 35658 189200
rect 35826 189144 37222 189200
rect 37390 189144 38786 189200
rect 38954 189144 40350 189200
rect 40518 189144 41914 189200
rect 42082 189144 43478 189200
rect 43646 189144 45042 189200
rect 45210 189144 46606 189200
rect 46774 189144 48170 189200
rect 48338 189144 49734 189200
rect 49902 189144 51298 189200
rect 51466 189144 52862 189200
rect 53030 189144 54426 189200
rect 54594 189144 55990 189200
rect 56158 189144 57554 189200
rect 57722 189144 59118 189200
rect 59286 189144 60682 189200
rect 60850 189144 62246 189200
rect 62414 189144 63810 189200
rect 63978 189144 65374 189200
rect 65542 189144 66938 189200
rect 67106 189144 68502 189200
rect 68670 189144 70066 189200
rect 70234 189144 71630 189200
rect 71798 189144 73194 189200
rect 73362 189144 74758 189200
rect 74926 189144 76322 189200
rect 76490 189144 77886 189200
rect 78054 189144 79450 189200
rect 79618 189144 81014 189200
rect 81182 189144 82578 189200
rect 82746 189144 84142 189200
rect 84310 189144 85706 189200
rect 85874 189144 87270 189200
rect 87438 189144 88834 189200
rect 89002 189144 90398 189200
rect 90566 189144 91962 189200
rect 92130 189144 93526 189200
rect 93694 189144 95090 189200
rect 95258 189144 96654 189200
rect 96822 189144 98218 189200
rect 98386 189144 99782 189200
rect 99950 189144 101346 189200
rect 101514 189144 102910 189200
rect 103078 189144 104474 189200
rect 104642 189144 106038 189200
rect 106206 189144 107602 189200
rect 107770 189144 109166 189200
rect 109334 189144 110730 189200
rect 110898 189144 112294 189200
rect 112462 189144 113858 189200
rect 114026 189144 115422 189200
rect 115590 189144 116986 189200
rect 117154 189144 118550 189200
rect 118718 189144 119122 189200
rect 938 856 119122 189144
rect 938 734 3090 856
rect 3258 734 4838 856
rect 5006 734 6586 856
rect 6754 734 8334 856
rect 8502 734 10082 856
rect 10250 734 11830 856
rect 11998 734 13578 856
rect 13746 734 15326 856
rect 15494 734 17074 856
rect 17242 734 18822 856
rect 18990 734 20570 856
rect 20738 734 22318 856
rect 22486 734 24066 856
rect 24234 734 25814 856
rect 25982 734 27562 856
rect 27730 734 29310 856
rect 29478 734 31058 856
rect 31226 734 32806 856
rect 32974 734 34554 856
rect 34722 734 36302 856
rect 36470 734 38050 856
rect 38218 734 39798 856
rect 39966 734 41546 856
rect 41714 734 43294 856
rect 43462 734 45042 856
rect 45210 734 46790 856
rect 46958 734 48538 856
rect 48706 734 50286 856
rect 50454 734 52034 856
rect 52202 734 53782 856
rect 53950 734 55530 856
rect 55698 734 57278 856
rect 57446 734 59026 856
rect 59194 734 60774 856
rect 60942 734 62522 856
rect 62690 734 64270 856
rect 64438 734 66018 856
rect 66186 734 67766 856
rect 67934 734 69514 856
rect 69682 734 71262 856
rect 71430 734 73010 856
rect 73178 734 74758 856
rect 74926 734 76506 856
rect 76674 734 78254 856
rect 78422 734 80002 856
rect 80170 734 81750 856
rect 81918 734 83498 856
rect 83666 734 85246 856
rect 85414 734 86994 856
rect 87162 734 88742 856
rect 88910 734 90490 856
rect 90658 734 92238 856
rect 92406 734 93986 856
rect 94154 734 95734 856
rect 95902 734 97482 856
rect 97650 734 99230 856
rect 99398 734 100978 856
rect 101146 734 102726 856
rect 102894 734 104474 856
rect 104642 734 106222 856
rect 106390 734 107970 856
rect 108138 734 109718 856
rect 109886 734 111466 856
rect 111634 734 113214 856
rect 113382 734 114962 856
rect 115130 734 116710 856
rect 116878 734 119122 856
<< metal3 >>
rect 0 182384 800 182504
rect 0 180616 800 180736
rect 0 178848 800 178968
rect 0 177080 800 177200
rect 0 175312 800 175432
rect 119200 173816 120000 173936
rect 0 173544 800 173664
rect 0 171776 800 171896
rect 0 170008 800 170128
rect 0 168240 800 168360
rect 0 166472 800 166592
rect 0 164704 800 164824
rect 0 162936 800 163056
rect 0 161168 800 161288
rect 0 159400 800 159520
rect 0 157632 800 157752
rect 0 155864 800 155984
rect 0 154096 800 154216
rect 0 152328 800 152448
rect 0 150560 800 150680
rect 0 148792 800 148912
rect 0 147024 800 147144
rect 0 145256 800 145376
rect 0 143488 800 143608
rect 119200 142264 120000 142384
rect 0 141720 800 141840
rect 0 139952 800 140072
rect 0 138184 800 138304
rect 0 136416 800 136536
rect 0 134648 800 134768
rect 0 132880 800 133000
rect 0 131112 800 131232
rect 0 129344 800 129464
rect 0 127576 800 127696
rect 0 125808 800 125928
rect 0 124040 800 124160
rect 0 122272 800 122392
rect 0 120504 800 120624
rect 0 118736 800 118856
rect 0 116968 800 117088
rect 0 115200 800 115320
rect 0 113432 800 113552
rect 0 111664 800 111784
rect 119200 110712 120000 110832
rect 0 109896 800 110016
rect 0 108128 800 108248
rect 0 106360 800 106480
rect 0 104592 800 104712
rect 0 102824 800 102944
rect 0 101056 800 101176
rect 0 99288 800 99408
rect 0 97520 800 97640
rect 0 95752 800 95872
rect 0 93984 800 94104
rect 0 92216 800 92336
rect 0 90448 800 90568
rect 0 88680 800 88800
rect 0 86912 800 87032
rect 0 85144 800 85264
rect 0 83376 800 83496
rect 0 81608 800 81728
rect 0 79840 800 79960
rect 119200 79160 120000 79280
rect 0 78072 800 78192
rect 0 76304 800 76424
rect 0 74536 800 74656
rect 0 72768 800 72888
rect 0 71000 800 71120
rect 0 69232 800 69352
rect 0 67464 800 67584
rect 0 65696 800 65816
rect 0 63928 800 64048
rect 0 62160 800 62280
rect 0 60392 800 60512
rect 0 58624 800 58744
rect 0 56856 800 56976
rect 0 55088 800 55208
rect 0 53320 800 53440
rect 0 51552 800 51672
rect 0 49784 800 49904
rect 0 48016 800 48136
rect 119200 47608 120000 47728
rect 0 46248 800 46368
rect 0 44480 800 44600
rect 0 42712 800 42832
rect 0 40944 800 41064
rect 0 39176 800 39296
rect 0 37408 800 37528
rect 0 35640 800 35760
rect 0 33872 800 33992
rect 0 32104 800 32224
rect 0 30336 800 30456
rect 0 28568 800 28688
rect 0 26800 800 26920
rect 0 25032 800 25152
rect 0 23264 800 23384
rect 0 21496 800 21616
rect 0 19728 800 19848
rect 0 17960 800 18080
rect 0 16192 800 16312
rect 119200 16056 120000 16176
rect 0 14424 800 14544
rect 0 12656 800 12776
rect 0 10888 800 11008
rect 0 9120 800 9240
rect 0 7352 800 7472
<< obsm3 >>
rect 800 182584 119200 187713
rect 880 182304 119200 182584
rect 800 180816 119200 182304
rect 880 180536 119200 180816
rect 800 179048 119200 180536
rect 880 178768 119200 179048
rect 800 177280 119200 178768
rect 880 177000 119200 177280
rect 800 175512 119200 177000
rect 880 175232 119200 175512
rect 800 174016 119200 175232
rect 800 173744 119120 174016
rect 880 173736 119120 173744
rect 880 173464 119200 173736
rect 800 171976 119200 173464
rect 880 171696 119200 171976
rect 800 170208 119200 171696
rect 880 169928 119200 170208
rect 800 168440 119200 169928
rect 880 168160 119200 168440
rect 800 166672 119200 168160
rect 880 166392 119200 166672
rect 800 164904 119200 166392
rect 880 164624 119200 164904
rect 800 163136 119200 164624
rect 880 162856 119200 163136
rect 800 161368 119200 162856
rect 880 161088 119200 161368
rect 800 159600 119200 161088
rect 880 159320 119200 159600
rect 800 157832 119200 159320
rect 880 157552 119200 157832
rect 800 156064 119200 157552
rect 880 155784 119200 156064
rect 800 154296 119200 155784
rect 880 154016 119200 154296
rect 800 152528 119200 154016
rect 880 152248 119200 152528
rect 800 150760 119200 152248
rect 880 150480 119200 150760
rect 800 148992 119200 150480
rect 880 148712 119200 148992
rect 800 147224 119200 148712
rect 880 146944 119200 147224
rect 800 145456 119200 146944
rect 880 145176 119200 145456
rect 800 143688 119200 145176
rect 880 143408 119200 143688
rect 800 142464 119200 143408
rect 800 142184 119120 142464
rect 800 141920 119200 142184
rect 880 141640 119200 141920
rect 800 140152 119200 141640
rect 880 139872 119200 140152
rect 800 138384 119200 139872
rect 880 138104 119200 138384
rect 800 136616 119200 138104
rect 880 136336 119200 136616
rect 800 134848 119200 136336
rect 880 134568 119200 134848
rect 800 133080 119200 134568
rect 880 132800 119200 133080
rect 800 131312 119200 132800
rect 880 131032 119200 131312
rect 800 129544 119200 131032
rect 880 129264 119200 129544
rect 800 127776 119200 129264
rect 880 127496 119200 127776
rect 800 126008 119200 127496
rect 880 125728 119200 126008
rect 800 124240 119200 125728
rect 880 123960 119200 124240
rect 800 122472 119200 123960
rect 880 122192 119200 122472
rect 800 120704 119200 122192
rect 880 120424 119200 120704
rect 800 118936 119200 120424
rect 880 118656 119200 118936
rect 800 117168 119200 118656
rect 880 116888 119200 117168
rect 800 115400 119200 116888
rect 880 115120 119200 115400
rect 800 113632 119200 115120
rect 880 113352 119200 113632
rect 800 111864 119200 113352
rect 880 111584 119200 111864
rect 800 110912 119200 111584
rect 800 110632 119120 110912
rect 800 110096 119200 110632
rect 880 109816 119200 110096
rect 800 108328 119200 109816
rect 880 108048 119200 108328
rect 800 106560 119200 108048
rect 880 106280 119200 106560
rect 800 104792 119200 106280
rect 880 104512 119200 104792
rect 800 103024 119200 104512
rect 880 102744 119200 103024
rect 800 101256 119200 102744
rect 880 100976 119200 101256
rect 800 99488 119200 100976
rect 880 99208 119200 99488
rect 800 97720 119200 99208
rect 880 97440 119200 97720
rect 800 95952 119200 97440
rect 880 95672 119200 95952
rect 800 94184 119200 95672
rect 880 93904 119200 94184
rect 800 92416 119200 93904
rect 880 92136 119200 92416
rect 800 90648 119200 92136
rect 880 90368 119200 90648
rect 800 88880 119200 90368
rect 880 88600 119200 88880
rect 800 87112 119200 88600
rect 880 86832 119200 87112
rect 800 85344 119200 86832
rect 880 85064 119200 85344
rect 800 83576 119200 85064
rect 880 83296 119200 83576
rect 800 81808 119200 83296
rect 880 81528 119200 81808
rect 800 80040 119200 81528
rect 880 79760 119200 80040
rect 800 79360 119200 79760
rect 800 79080 119120 79360
rect 800 78272 119200 79080
rect 880 77992 119200 78272
rect 800 76504 119200 77992
rect 880 76224 119200 76504
rect 800 74736 119200 76224
rect 880 74456 119200 74736
rect 800 72968 119200 74456
rect 880 72688 119200 72968
rect 800 71200 119200 72688
rect 880 70920 119200 71200
rect 800 69432 119200 70920
rect 880 69152 119200 69432
rect 800 67664 119200 69152
rect 880 67384 119200 67664
rect 800 65896 119200 67384
rect 880 65616 119200 65896
rect 800 64128 119200 65616
rect 880 63848 119200 64128
rect 800 62360 119200 63848
rect 880 62080 119200 62360
rect 800 60592 119200 62080
rect 880 60312 119200 60592
rect 800 58824 119200 60312
rect 880 58544 119200 58824
rect 800 57056 119200 58544
rect 880 56776 119200 57056
rect 800 55288 119200 56776
rect 880 55008 119200 55288
rect 800 53520 119200 55008
rect 880 53240 119200 53520
rect 800 51752 119200 53240
rect 880 51472 119200 51752
rect 800 49984 119200 51472
rect 880 49704 119200 49984
rect 800 48216 119200 49704
rect 880 47936 119200 48216
rect 800 47808 119200 47936
rect 800 47528 119120 47808
rect 800 46448 119200 47528
rect 880 46168 119200 46448
rect 800 44680 119200 46168
rect 880 44400 119200 44680
rect 800 42912 119200 44400
rect 880 42632 119200 42912
rect 800 41144 119200 42632
rect 880 40864 119200 41144
rect 800 39376 119200 40864
rect 880 39096 119200 39376
rect 800 37608 119200 39096
rect 880 37328 119200 37608
rect 800 35840 119200 37328
rect 880 35560 119200 35840
rect 800 34072 119200 35560
rect 880 33792 119200 34072
rect 800 32304 119200 33792
rect 880 32024 119200 32304
rect 800 30536 119200 32024
rect 880 30256 119200 30536
rect 800 28768 119200 30256
rect 880 28488 119200 28768
rect 800 27000 119200 28488
rect 880 26720 119200 27000
rect 800 25232 119200 26720
rect 880 24952 119200 25232
rect 800 23464 119200 24952
rect 880 23184 119200 23464
rect 800 21696 119200 23184
rect 880 21416 119200 21696
rect 800 19928 119200 21416
rect 880 19648 119200 19928
rect 800 18160 119200 19648
rect 880 17880 119200 18160
rect 800 16392 119200 17880
rect 880 16256 119200 16392
rect 880 16112 119120 16256
rect 800 15976 119120 16112
rect 800 14624 119200 15976
rect 880 14344 119200 14624
rect 800 12856 119200 14344
rect 880 12576 119200 12856
rect 800 11088 119200 12576
rect 880 10808 119200 11088
rect 800 9320 119200 10808
rect 880 9040 119200 9320
rect 800 7552 119200 9040
rect 880 7272 119200 7552
rect 800 2143 119200 7272
<< metal4 >>
rect 4208 2128 4528 187728
rect 19568 2128 19888 187728
rect 34928 2128 35248 187728
rect 50288 2128 50608 187728
rect 65648 2128 65968 187728
rect 81008 2128 81328 187728
rect 96368 2128 96688 187728
rect 111728 2128 112048 187728
<< obsm4 >>
rect 1715 2211 4128 187509
rect 4608 2211 19488 187509
rect 19968 2211 34848 187509
rect 35328 2211 50208 187509
rect 50688 2211 65568 187509
rect 66048 2211 80928 187509
rect 81408 2211 96288 187509
rect 96768 2211 108685 187509
<< labels >>
rlabel metal2 s 73066 0 73122 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 1306 189200 1362 190000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 16946 189200 17002 190000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 18510 189200 18566 190000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 20074 189200 20130 190000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 21638 189200 21694 190000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 23202 189200 23258 190000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 24766 189200 24822 190000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 26330 189200 26386 190000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 27894 189200 27950 190000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 29458 189200 29514 190000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 31022 189200 31078 190000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 2870 189200 2926 190000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 32586 189200 32642 190000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 34150 189200 34206 190000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 35714 189200 35770 190000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 37278 189200 37334 190000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 38842 189200 38898 190000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 40406 189200 40462 190000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 41970 189200 42026 190000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 43534 189200 43590 190000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 45098 189200 45154 190000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 46662 189200 46718 190000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 4434 189200 4490 190000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 48226 189200 48282 190000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 49790 189200 49846 190000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 51354 189200 51410 190000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 52918 189200 52974 190000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 54482 189200 54538 190000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 56046 189200 56102 190000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 57610 189200 57666 190000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 59174 189200 59230 190000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 5998 189200 6054 190000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 7562 189200 7618 190000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 9126 189200 9182 190000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 10690 189200 10746 190000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 12254 189200 12310 190000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 13818 189200 13874 190000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 15382 189200 15438 190000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 60738 189200 60794 190000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 76378 189200 76434 190000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 77942 189200 77998 190000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 79506 189200 79562 190000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 81070 189200 81126 190000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 82634 189200 82690 190000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 84198 189200 84254 190000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 85762 189200 85818 190000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 87326 189200 87382 190000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 88890 189200 88946 190000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 90454 189200 90510 190000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 62302 189200 62358 190000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 92018 189200 92074 190000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 93582 189200 93638 190000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 95146 189200 95202 190000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 96710 189200 96766 190000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 98274 189200 98330 190000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 99838 189200 99894 190000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 101402 189200 101458 190000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 102966 189200 103022 190000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 104530 189200 104586 190000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 106094 189200 106150 190000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 63866 189200 63922 190000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 107658 189200 107714 190000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 109222 189200 109278 190000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 110786 189200 110842 190000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 112350 189200 112406 190000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 113914 189200 113970 190000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 115478 189200 115534 190000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 117042 189200 117098 190000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 118606 189200 118662 190000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 65430 189200 65486 190000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 66994 189200 67050 190000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 68558 189200 68614 190000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 70122 189200 70178 190000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 71686 189200 71742 190000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 73250 189200 73306 190000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 74814 189200 74870 190000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 119200 79160 120000 79280 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 119200 110712 120000 110832 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 119200 142264 120000 142384 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 119200 173816 120000 173936 6 jtag_tms
port 128 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 peripheral_irq[0]
port 129 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 peripheral_irq[1]
port 130 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 peripheral_irq[2]
port 131 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 peripheral_irq[3]
port 132 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 peripheral_irq[4]
port 133 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 peripheral_irq[5]
port 134 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 peripheral_irq[6]
port 135 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 peripheral_irq[7]
port 136 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 peripheral_irq[8]
port 137 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 peripheral_irq[9]
port 138 nsew signal output
rlabel metal3 s 119200 16056 120000 16176 6 probe_blink[0]
port 139 nsew signal output
rlabel metal3 s 119200 47608 120000 47728 6 probe_blink[1]
port 140 nsew signal output
rlabel metal4 s 4208 2128 4528 187728 6 vccd1
port 141 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 187728 6 vccd1
port 141 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 187728 6 vccd1
port 141 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 187728 6 vccd1
port 141 nsew power bidirectional
rlabel metal2 s 108026 0 108082 800 6 vga_b[0]
port 142 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 vga_b[1]
port 143 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 vga_g[0]
port 144 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 vga_g[1]
port 145 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 vga_hsync
port 146 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 vga_r[0]
port 147 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 vga_r[1]
port 148 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 vga_vsync
port 149 nsew signal input
rlabel metal4 s 19568 2128 19888 187728 6 vssd1
port 150 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 187728 6 vssd1
port 150 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 187728 6 vssd1
port 150 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 187728 6 vssd1
port 150 nsew ground bidirectional
rlabel metal3 s 0 7352 800 7472 6 wb_ack_o
port 151 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[0]
port 152 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 wb_adr_i[10]
port 153 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 wb_adr_i[11]
port 154 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 wb_adr_i[12]
port 155 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 wb_adr_i[13]
port 156 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 wb_adr_i[14]
port 157 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 wb_adr_i[15]
port 158 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 wb_adr_i[16]
port 159 nsew signal input
rlabel metal3 s 0 118736 800 118856 6 wb_adr_i[17]
port 160 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 wb_adr_i[18]
port 161 nsew signal input
rlabel metal3 s 0 129344 800 129464 6 wb_adr_i[19]
port 162 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wb_adr_i[1]
port 163 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 wb_adr_i[20]
port 164 nsew signal input
rlabel metal3 s 0 139952 800 140072 6 wb_adr_i[21]
port 165 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 wb_adr_i[22]
port 166 nsew signal input
rlabel metal3 s 0 150560 800 150680 6 wb_adr_i[23]
port 167 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 wb_adr_i[2]
port 168 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 wb_adr_i[3]
port 169 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 wb_adr_i[4]
port 170 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 wb_adr_i[5]
port 171 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 wb_adr_i[6]
port 172 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 wb_adr_i[7]
port 173 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 wb_adr_i[8]
port 174 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 wb_adr_i[9]
port 175 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wb_clk_i
port 176 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wb_cyc_i
port 177 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 wb_data_i[0]
port 178 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 wb_data_i[10]
port 179 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 wb_data_i[11]
port 180 nsew signal input
rlabel metal3 s 0 93984 800 94104 6 wb_data_i[12]
port 181 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 wb_data_i[13]
port 182 nsew signal input
rlabel metal3 s 0 104592 800 104712 6 wb_data_i[14]
port 183 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 wb_data_i[15]
port 184 nsew signal input
rlabel metal3 s 0 115200 800 115320 6 wb_data_i[16]
port 185 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 wb_data_i[17]
port 186 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 wb_data_i[18]
port 187 nsew signal input
rlabel metal3 s 0 131112 800 131232 6 wb_data_i[19]
port 188 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_data_i[1]
port 189 nsew signal input
rlabel metal3 s 0 136416 800 136536 6 wb_data_i[20]
port 190 nsew signal input
rlabel metal3 s 0 141720 800 141840 6 wb_data_i[21]
port 191 nsew signal input
rlabel metal3 s 0 147024 800 147144 6 wb_data_i[22]
port 192 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 wb_data_i[23]
port 193 nsew signal input
rlabel metal3 s 0 155864 800 155984 6 wb_data_i[24]
port 194 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 wb_data_i[25]
port 195 nsew signal input
rlabel metal3 s 0 162936 800 163056 6 wb_data_i[26]
port 196 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 wb_data_i[27]
port 197 nsew signal input
rlabel metal3 s 0 170008 800 170128 6 wb_data_i[28]
port 198 nsew signal input
rlabel metal3 s 0 173544 800 173664 6 wb_data_i[29]
port 199 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 wb_data_i[2]
port 200 nsew signal input
rlabel metal3 s 0 177080 800 177200 6 wb_data_i[30]
port 201 nsew signal input
rlabel metal3 s 0 180616 800 180736 6 wb_data_i[31]
port 202 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 wb_data_i[3]
port 203 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 wb_data_i[4]
port 204 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 wb_data_i[5]
port 205 nsew signal input
rlabel metal3 s 0 62160 800 62280 6 wb_data_i[6]
port 206 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 wb_data_i[7]
port 207 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 wb_data_i[8]
port 208 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 wb_data_i[9]
port 209 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 wb_data_o[0]
port 210 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 wb_data_o[10]
port 211 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 wb_data_o[11]
port 212 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 wb_data_o[12]
port 213 nsew signal output
rlabel metal3 s 0 101056 800 101176 6 wb_data_o[13]
port 214 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 wb_data_o[14]
port 215 nsew signal output
rlabel metal3 s 0 111664 800 111784 6 wb_data_o[15]
port 216 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 wb_data_o[16]
port 217 nsew signal output
rlabel metal3 s 0 122272 800 122392 6 wb_data_o[17]
port 218 nsew signal output
rlabel metal3 s 0 127576 800 127696 6 wb_data_o[18]
port 219 nsew signal output
rlabel metal3 s 0 132880 800 133000 6 wb_data_o[19]
port 220 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 wb_data_o[1]
port 221 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 wb_data_o[20]
port 222 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 wb_data_o[21]
port 223 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 wb_data_o[22]
port 224 nsew signal output
rlabel metal3 s 0 154096 800 154216 6 wb_data_o[23]
port 225 nsew signal output
rlabel metal3 s 0 157632 800 157752 6 wb_data_o[24]
port 226 nsew signal output
rlabel metal3 s 0 161168 800 161288 6 wb_data_o[25]
port 227 nsew signal output
rlabel metal3 s 0 164704 800 164824 6 wb_data_o[26]
port 228 nsew signal output
rlabel metal3 s 0 168240 800 168360 6 wb_data_o[27]
port 229 nsew signal output
rlabel metal3 s 0 171776 800 171896 6 wb_data_o[28]
port 230 nsew signal output
rlabel metal3 s 0 175312 800 175432 6 wb_data_o[29]
port 231 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 wb_data_o[2]
port 232 nsew signal output
rlabel metal3 s 0 178848 800 178968 6 wb_data_o[30]
port 233 nsew signal output
rlabel metal3 s 0 182384 800 182504 6 wb_data_o[31]
port 234 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 wb_data_o[3]
port 235 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 wb_data_o[4]
port 236 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 wb_data_o[5]
port 237 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 wb_data_o[6]
port 238 nsew signal output
rlabel metal3 s 0 69232 800 69352 6 wb_data_o[7]
port 239 nsew signal output
rlabel metal3 s 0 74536 800 74656 6 wb_data_o[8]
port 240 nsew signal output
rlabel metal3 s 0 79840 800 79960 6 wb_data_o[9]
port 241 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 wb_error_o
port 242 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 wb_rst_i
port 243 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 wb_sel_i[0]
port 244 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 wb_sel_i[1]
port 245 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 wb_sel_i[2]
port 246 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 wb_sel_i[3]
port 247 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 wb_stall_o
port 248 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 wb_stb_i
port 249 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 wb_we_i
port 250 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 190000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 51541376
string GDS_FILE /mnt/f/WSL/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/23_05_10_23_54/results/signoff/Peripherals.magic.gds
string GDS_START 1351076
<< end >>

