magic
tech sky130A
magscale 1 2
timestamp 1651278901
<< obsli1 >>
rect 1104 2159 78844 92497
<< obsm1 >>
rect 566 2128 78844 92528
<< metal2 >>
rect 40038 94200 40094 95000
rect 19982 0 20038 800
rect 60002 0 60058 800
<< obsm2 >>
rect 478 94144 39982 94489
rect 40150 94144 78090 94489
rect 478 856 78090 94144
rect 478 439 19926 856
rect 20094 439 59946 856
rect 60114 439 78090 856
<< metal3 >>
rect 0 94392 800 94512
rect 0 93304 800 93424
rect 79200 93440 80000 93560
rect 0 92216 800 92336
rect 0 91264 800 91384
rect 79200 90448 80000 90568
rect 0 90176 800 90296
rect 0 89088 800 89208
rect 0 88136 800 88256
rect 79200 87456 80000 87576
rect 0 87048 800 87168
rect 0 85960 800 86080
rect 0 85008 800 85128
rect 79200 84464 80000 84584
rect 0 83920 800 84040
rect 0 82832 800 82952
rect 0 81880 800 82000
rect 79200 81472 80000 81592
rect 0 80792 800 80912
rect 0 79704 800 79824
rect 0 78752 800 78872
rect 79200 78480 80000 78600
rect 0 77664 800 77784
rect 0 76576 800 76696
rect 0 75624 800 75744
rect 79200 75624 80000 75744
rect 0 74536 800 74656
rect 0 73448 800 73568
rect 0 72496 800 72616
rect 79200 72632 80000 72752
rect 0 71408 800 71528
rect 0 70320 800 70440
rect 79200 69640 80000 69760
rect 0 69232 800 69352
rect 0 68280 800 68400
rect 0 67192 800 67312
rect 79200 66648 80000 66768
rect 0 66104 800 66224
rect 0 65152 800 65272
rect 0 64064 800 64184
rect 79200 63656 80000 63776
rect 0 62976 800 63096
rect 0 62024 800 62144
rect 0 60936 800 61056
rect 79200 60664 80000 60784
rect 0 59848 800 59968
rect 0 58896 800 59016
rect 0 57808 800 57928
rect 79200 57808 80000 57928
rect 0 56720 800 56840
rect 0 55768 800 55888
rect 0 54680 800 54800
rect 79200 54816 80000 54936
rect 0 53592 800 53712
rect 0 52640 800 52760
rect 79200 51824 80000 51944
rect 0 51552 800 51672
rect 0 50464 800 50584
rect 0 49512 800 49632
rect 79200 48832 80000 48952
rect 0 48424 800 48544
rect 0 47336 800 47456
rect 0 46248 800 46368
rect 79200 45840 80000 45960
rect 0 45296 800 45416
rect 0 44208 800 44328
rect 0 43120 800 43240
rect 79200 42848 80000 42968
rect 0 42168 800 42288
rect 0 41080 800 41200
rect 0 39992 800 40112
rect 79200 39856 80000 39976
rect 0 39040 800 39160
rect 0 37952 800 38072
rect 0 36864 800 36984
rect 79200 37000 80000 37120
rect 0 35912 800 36032
rect 0 34824 800 34944
rect 79200 34008 80000 34128
rect 0 33736 800 33856
rect 0 32784 800 32904
rect 0 31696 800 31816
rect 79200 31016 80000 31136
rect 0 30608 800 30728
rect 0 29656 800 29776
rect 0 28568 800 28688
rect 79200 28024 80000 28144
rect 0 27480 800 27600
rect 0 26528 800 26648
rect 0 25440 800 25560
rect 79200 25032 80000 25152
rect 0 24352 800 24472
rect 0 23264 800 23384
rect 0 22312 800 22432
rect 79200 22040 80000 22160
rect 0 21224 800 21344
rect 0 20136 800 20256
rect 0 19184 800 19304
rect 79200 19184 80000 19304
rect 0 18096 800 18216
rect 0 17008 800 17128
rect 0 16056 800 16176
rect 79200 16192 80000 16312
rect 0 14968 800 15088
rect 0 13880 800 14000
rect 79200 13200 80000 13320
rect 0 12928 800 13048
rect 0 11840 800 11960
rect 0 10752 800 10872
rect 79200 10208 80000 10328
rect 0 9800 800 9920
rect 0 8712 800 8832
rect 0 7624 800 7744
rect 79200 7216 80000 7336
rect 0 6672 800 6792
rect 0 5584 800 5704
rect 0 4496 800 4616
rect 79200 4224 80000 4344
rect 0 3544 800 3664
rect 0 2456 800 2576
rect 0 1368 800 1488
rect 79200 1368 80000 1488
rect 0 416 800 536
<< obsm3 >>
rect 880 94312 79200 94485
rect 473 93640 79200 94312
rect 473 93504 79120 93640
rect 880 93360 79120 93504
rect 880 93224 79200 93360
rect 473 92416 79200 93224
rect 880 92136 79200 92416
rect 473 91464 79200 92136
rect 880 91184 79200 91464
rect 473 90648 79200 91184
rect 473 90376 79120 90648
rect 880 90368 79120 90376
rect 880 90096 79200 90368
rect 473 89288 79200 90096
rect 880 89008 79200 89288
rect 473 88336 79200 89008
rect 880 88056 79200 88336
rect 473 87656 79200 88056
rect 473 87376 79120 87656
rect 473 87248 79200 87376
rect 880 86968 79200 87248
rect 473 86160 79200 86968
rect 880 85880 79200 86160
rect 473 85208 79200 85880
rect 880 84928 79200 85208
rect 473 84664 79200 84928
rect 473 84384 79120 84664
rect 473 84120 79200 84384
rect 880 83840 79200 84120
rect 473 83032 79200 83840
rect 880 82752 79200 83032
rect 473 82080 79200 82752
rect 880 81800 79200 82080
rect 473 81672 79200 81800
rect 473 81392 79120 81672
rect 473 80992 79200 81392
rect 880 80712 79200 80992
rect 473 79904 79200 80712
rect 880 79624 79200 79904
rect 473 78952 79200 79624
rect 880 78680 79200 78952
rect 880 78672 79120 78680
rect 473 78400 79120 78672
rect 473 77864 79200 78400
rect 880 77584 79200 77864
rect 473 76776 79200 77584
rect 880 76496 79200 76776
rect 473 75824 79200 76496
rect 880 75544 79120 75824
rect 473 74736 79200 75544
rect 880 74456 79200 74736
rect 473 73648 79200 74456
rect 880 73368 79200 73648
rect 473 72832 79200 73368
rect 473 72696 79120 72832
rect 880 72552 79120 72696
rect 880 72416 79200 72552
rect 473 71608 79200 72416
rect 880 71328 79200 71608
rect 473 70520 79200 71328
rect 880 70240 79200 70520
rect 473 69840 79200 70240
rect 473 69560 79120 69840
rect 473 69432 79200 69560
rect 880 69152 79200 69432
rect 473 68480 79200 69152
rect 880 68200 79200 68480
rect 473 67392 79200 68200
rect 880 67112 79200 67392
rect 473 66848 79200 67112
rect 473 66568 79120 66848
rect 473 66304 79200 66568
rect 880 66024 79200 66304
rect 473 65352 79200 66024
rect 880 65072 79200 65352
rect 473 64264 79200 65072
rect 880 63984 79200 64264
rect 473 63856 79200 63984
rect 473 63576 79120 63856
rect 473 63176 79200 63576
rect 880 62896 79200 63176
rect 473 62224 79200 62896
rect 880 61944 79200 62224
rect 473 61136 79200 61944
rect 880 60864 79200 61136
rect 880 60856 79120 60864
rect 473 60584 79120 60856
rect 473 60048 79200 60584
rect 880 59768 79200 60048
rect 473 59096 79200 59768
rect 880 58816 79200 59096
rect 473 58008 79200 58816
rect 880 57728 79120 58008
rect 473 56920 79200 57728
rect 880 56640 79200 56920
rect 473 55968 79200 56640
rect 880 55688 79200 55968
rect 473 55016 79200 55688
rect 473 54880 79120 55016
rect 880 54736 79120 54880
rect 880 54600 79200 54736
rect 473 53792 79200 54600
rect 880 53512 79200 53792
rect 473 52840 79200 53512
rect 880 52560 79200 52840
rect 473 52024 79200 52560
rect 473 51752 79120 52024
rect 880 51744 79120 51752
rect 880 51472 79200 51744
rect 473 50664 79200 51472
rect 880 50384 79200 50664
rect 473 49712 79200 50384
rect 880 49432 79200 49712
rect 473 49032 79200 49432
rect 473 48752 79120 49032
rect 473 48624 79200 48752
rect 880 48344 79200 48624
rect 473 47536 79200 48344
rect 880 47256 79200 47536
rect 473 46448 79200 47256
rect 880 46168 79200 46448
rect 473 46040 79200 46168
rect 473 45760 79120 46040
rect 473 45496 79200 45760
rect 880 45216 79200 45496
rect 473 44408 79200 45216
rect 880 44128 79200 44408
rect 473 43320 79200 44128
rect 880 43048 79200 43320
rect 880 43040 79120 43048
rect 473 42768 79120 43040
rect 473 42368 79200 42768
rect 880 42088 79200 42368
rect 473 41280 79200 42088
rect 880 41000 79200 41280
rect 473 40192 79200 41000
rect 880 40056 79200 40192
rect 880 39912 79120 40056
rect 473 39776 79120 39912
rect 473 39240 79200 39776
rect 880 38960 79200 39240
rect 473 38152 79200 38960
rect 880 37872 79200 38152
rect 473 37200 79200 37872
rect 473 37064 79120 37200
rect 880 36920 79120 37064
rect 880 36784 79200 36920
rect 473 36112 79200 36784
rect 880 35832 79200 36112
rect 473 35024 79200 35832
rect 880 34744 79200 35024
rect 473 34208 79200 34744
rect 473 33936 79120 34208
rect 880 33928 79120 33936
rect 880 33656 79200 33928
rect 473 32984 79200 33656
rect 880 32704 79200 32984
rect 473 31896 79200 32704
rect 880 31616 79200 31896
rect 473 31216 79200 31616
rect 473 30936 79120 31216
rect 473 30808 79200 30936
rect 880 30528 79200 30808
rect 473 29856 79200 30528
rect 880 29576 79200 29856
rect 473 28768 79200 29576
rect 880 28488 79200 28768
rect 473 28224 79200 28488
rect 473 27944 79120 28224
rect 473 27680 79200 27944
rect 880 27400 79200 27680
rect 473 26728 79200 27400
rect 880 26448 79200 26728
rect 473 25640 79200 26448
rect 880 25360 79200 25640
rect 473 25232 79200 25360
rect 473 24952 79120 25232
rect 473 24552 79200 24952
rect 880 24272 79200 24552
rect 473 23464 79200 24272
rect 880 23184 79200 23464
rect 473 22512 79200 23184
rect 880 22240 79200 22512
rect 880 22232 79120 22240
rect 473 21960 79120 22232
rect 473 21424 79200 21960
rect 880 21144 79200 21424
rect 473 20336 79200 21144
rect 880 20056 79200 20336
rect 473 19384 79200 20056
rect 880 19104 79120 19384
rect 473 18296 79200 19104
rect 880 18016 79200 18296
rect 473 17208 79200 18016
rect 880 16928 79200 17208
rect 473 16392 79200 16928
rect 473 16256 79120 16392
rect 880 16112 79120 16256
rect 880 15976 79200 16112
rect 473 15168 79200 15976
rect 880 14888 79200 15168
rect 473 14080 79200 14888
rect 880 13800 79200 14080
rect 473 13400 79200 13800
rect 473 13128 79120 13400
rect 880 13120 79120 13128
rect 880 12848 79200 13120
rect 473 12040 79200 12848
rect 880 11760 79200 12040
rect 473 10952 79200 11760
rect 880 10672 79200 10952
rect 473 10408 79200 10672
rect 473 10128 79120 10408
rect 473 10000 79200 10128
rect 880 9720 79200 10000
rect 473 8912 79200 9720
rect 880 8632 79200 8912
rect 473 7824 79200 8632
rect 880 7544 79200 7824
rect 473 7416 79200 7544
rect 473 7136 79120 7416
rect 473 6872 79200 7136
rect 880 6592 79200 6872
rect 473 5784 79200 6592
rect 880 5504 79200 5784
rect 473 4696 79200 5504
rect 880 4424 79200 4696
rect 880 4416 79120 4424
rect 473 4144 79120 4416
rect 473 3744 79200 4144
rect 880 3464 79200 3744
rect 473 2656 79200 3464
rect 880 2376 79200 2656
rect 473 1568 79200 2376
rect 880 1288 79120 1568
rect 473 616 79200 1288
rect 880 443 79200 616
<< metal4 >>
rect 4208 2128 4528 92528
rect 19568 2128 19888 92528
rect 34928 2128 35248 92528
rect 50288 2128 50608 92528
rect 65648 2128 65968 92528
<< labels >>
rlabel metal2 s 19982 0 20038 800 6 clk
port 1 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 peripheralBus_address[0]
port 2 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 peripheralBus_address[10]
port 3 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 peripheralBus_address[11]
port 4 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 peripheralBus_address[12]
port 5 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 peripheralBus_address[13]
port 6 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 peripheralBus_address[14]
port 7 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 peripheralBus_address[15]
port 8 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 peripheralBus_address[16]
port 9 nsew signal input
rlabel metal3 s 0 56720 800 56840 6 peripheralBus_address[17]
port 10 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 peripheralBus_address[18]
port 11 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 peripheralBus_address[19]
port 12 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 peripheralBus_address[1]
port 13 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 peripheralBus_address[20]
port 14 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 peripheralBus_address[21]
port 15 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 peripheralBus_address[22]
port 16 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 peripheralBus_address[23]
port 17 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 peripheralBus_address[2]
port 18 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 peripheralBus_address[3]
port 19 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 peripheralBus_address[4]
port 20 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 peripheralBus_address[5]
port 21 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 peripheralBus_address[6]
port 22 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 peripheralBus_address[7]
port 23 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 peripheralBus_address[8]
port 24 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 peripheralBus_address[9]
port 25 nsew signal input
rlabel metal3 s 0 416 800 536 6 peripheralBus_busy
port 26 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 peripheralBus_dataIn[0]
port 27 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 peripheralBus_dataIn[10]
port 28 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 peripheralBus_dataIn[11]
port 29 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 peripheralBus_dataIn[12]
port 30 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 peripheralBus_dataIn[13]
port 31 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 peripheralBus_dataIn[14]
port 32 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 peripheralBus_dataIn[15]
port 33 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 peripheralBus_dataIn[16]
port 34 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 peripheralBus_dataIn[17]
port 35 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 peripheralBus_dataIn[18]
port 36 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 peripheralBus_dataIn[19]
port 37 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 peripheralBus_dataIn[1]
port 38 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 peripheralBus_dataIn[20]
port 39 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 peripheralBus_dataIn[21]
port 40 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 peripheralBus_dataIn[22]
port 41 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 peripheralBus_dataIn[23]
port 42 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 peripheralBus_dataIn[24]
port 43 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 peripheralBus_dataIn[25]
port 44 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 peripheralBus_dataIn[26]
port 45 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 peripheralBus_dataIn[27]
port 46 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 peripheralBus_dataIn[28]
port 47 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 peripheralBus_dataIn[29]
port 48 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 peripheralBus_dataIn[2]
port 49 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 peripheralBus_dataIn[30]
port 50 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 peripheralBus_dataIn[31]
port 51 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 peripheralBus_dataIn[3]
port 52 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 peripheralBus_dataIn[4]
port 53 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 peripheralBus_dataIn[5]
port 54 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 peripheralBus_dataIn[6]
port 55 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 peripheralBus_dataIn[7]
port 56 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 peripheralBus_dataIn[8]
port 57 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 peripheralBus_dataIn[9]
port 58 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 peripheralBus_dataOut[0]
port 59 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 peripheralBus_dataOut[10]
port 60 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 peripheralBus_dataOut[11]
port 61 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 peripheralBus_dataOut[12]
port 62 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 peripheralBus_dataOut[13]
port 63 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 peripheralBus_dataOut[14]
port 64 nsew signal output
rlabel metal3 s 0 52640 800 52760 6 peripheralBus_dataOut[15]
port 65 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 peripheralBus_dataOut[16]
port 66 nsew signal output
rlabel metal3 s 0 58896 800 59016 6 peripheralBus_dataOut[17]
port 67 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 peripheralBus_dataOut[18]
port 68 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 peripheralBus_dataOut[19]
port 69 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 peripheralBus_dataOut[1]
port 70 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 peripheralBus_dataOut[20]
port 71 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 peripheralBus_dataOut[21]
port 72 nsew signal output
rlabel metal3 s 0 74536 800 74656 6 peripheralBus_dataOut[22]
port 73 nsew signal output
rlabel metal3 s 0 77664 800 77784 6 peripheralBus_dataOut[23]
port 74 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 peripheralBus_dataOut[24]
port 75 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 peripheralBus_dataOut[25]
port 76 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 peripheralBus_dataOut[26]
port 77 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 peripheralBus_dataOut[27]
port 78 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 peripheralBus_dataOut[28]
port 79 nsew signal output
rlabel metal3 s 0 90176 800 90296 6 peripheralBus_dataOut[29]
port 80 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 peripheralBus_dataOut[2]
port 81 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 peripheralBus_dataOut[30]
port 82 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 peripheralBus_dataOut[31]
port 83 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 peripheralBus_dataOut[3]
port 84 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 peripheralBus_dataOut[4]
port 85 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 peripheralBus_dataOut[5]
port 86 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 peripheralBus_dataOut[6]
port 87 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 peripheralBus_dataOut[7]
port 88 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 peripheralBus_dataOut[8]
port 89 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 peripheralBus_dataOut[9]
port 90 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 peripheralBus_oe
port 91 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 peripheralBus_we
port 92 nsew signal input
rlabel metal3 s 79200 1368 80000 1488 6 pwm_en[0]
port 93 nsew signal output
rlabel metal3 s 79200 60664 80000 60784 6 pwm_en[10]
port 94 nsew signal output
rlabel metal3 s 79200 66648 80000 66768 6 pwm_en[11]
port 95 nsew signal output
rlabel metal3 s 79200 72632 80000 72752 6 pwm_en[12]
port 96 nsew signal output
rlabel metal3 s 79200 78480 80000 78600 6 pwm_en[13]
port 97 nsew signal output
rlabel metal3 s 79200 84464 80000 84584 6 pwm_en[14]
port 98 nsew signal output
rlabel metal3 s 79200 90448 80000 90568 6 pwm_en[15]
port 99 nsew signal output
rlabel metal3 s 79200 7216 80000 7336 6 pwm_en[1]
port 100 nsew signal output
rlabel metal3 s 79200 13200 80000 13320 6 pwm_en[2]
port 101 nsew signal output
rlabel metal3 s 79200 19184 80000 19304 6 pwm_en[3]
port 102 nsew signal output
rlabel metal3 s 79200 25032 80000 25152 6 pwm_en[4]
port 103 nsew signal output
rlabel metal3 s 79200 31016 80000 31136 6 pwm_en[5]
port 104 nsew signal output
rlabel metal3 s 79200 37000 80000 37120 6 pwm_en[6]
port 105 nsew signal output
rlabel metal3 s 79200 42848 80000 42968 6 pwm_en[7]
port 106 nsew signal output
rlabel metal3 s 79200 48832 80000 48952 6 pwm_en[8]
port 107 nsew signal output
rlabel metal3 s 79200 54816 80000 54936 6 pwm_en[9]
port 108 nsew signal output
rlabel metal3 s 79200 4224 80000 4344 6 pwm_out[0]
port 109 nsew signal output
rlabel metal3 s 79200 63656 80000 63776 6 pwm_out[10]
port 110 nsew signal output
rlabel metal3 s 79200 69640 80000 69760 6 pwm_out[11]
port 111 nsew signal output
rlabel metal3 s 79200 75624 80000 75744 6 pwm_out[12]
port 112 nsew signal output
rlabel metal3 s 79200 81472 80000 81592 6 pwm_out[13]
port 113 nsew signal output
rlabel metal3 s 79200 87456 80000 87576 6 pwm_out[14]
port 114 nsew signal output
rlabel metal3 s 79200 93440 80000 93560 6 pwm_out[15]
port 115 nsew signal output
rlabel metal3 s 79200 10208 80000 10328 6 pwm_out[1]
port 116 nsew signal output
rlabel metal3 s 79200 16192 80000 16312 6 pwm_out[2]
port 117 nsew signal output
rlabel metal3 s 79200 22040 80000 22160 6 pwm_out[3]
port 118 nsew signal output
rlabel metal3 s 79200 28024 80000 28144 6 pwm_out[4]
port 119 nsew signal output
rlabel metal3 s 79200 34008 80000 34128 6 pwm_out[5]
port 120 nsew signal output
rlabel metal3 s 79200 39856 80000 39976 6 pwm_out[6]
port 121 nsew signal output
rlabel metal3 s 79200 45840 80000 45960 6 pwm_out[7]
port 122 nsew signal output
rlabel metal3 s 79200 51824 80000 51944 6 pwm_out[8]
port 123 nsew signal output
rlabel metal3 s 79200 57808 80000 57928 6 pwm_out[9]
port 124 nsew signal output
rlabel metal2 s 40038 94200 40094 95000 6 requestOutput
port 125 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 rst
port 126 nsew signal input
rlabel metal4 s 4208 2128 4528 92528 6 vccd1
port 127 nsew power input
rlabel metal4 s 34928 2128 35248 92528 6 vccd1
port 127 nsew power input
rlabel metal4 s 65648 2128 65968 92528 6 vccd1
port 127 nsew power input
rlabel metal4 s 19568 2128 19888 92528 6 vssd1
port 128 nsew ground input
rlabel metal4 s 50288 2128 50608 92528 6 vssd1
port 128 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 95000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17534950
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripheral_PWM/runs/Peripheral_PWM/results/finishing/PWM.magic.gds
string GDS_START 765714
<< end >>

