magic
tech sky130A
magscale 1 2
timestamp 1653084718
<< obsli1 >>
rect 1104 2159 68816 97393
<< obsm1 >>
rect 14 1504 69998 98116
<< metal2 >>
rect 202 99200 258 100000
rect 662 99200 718 100000
rect 1122 99200 1178 100000
rect 1674 99200 1730 100000
rect 2134 99200 2190 100000
rect 2594 99200 2650 100000
rect 3146 99200 3202 100000
rect 3606 99200 3662 100000
rect 4066 99200 4122 100000
rect 4618 99200 4674 100000
rect 5078 99200 5134 100000
rect 5538 99200 5594 100000
rect 6090 99200 6146 100000
rect 6550 99200 6606 100000
rect 7102 99200 7158 100000
rect 7562 99200 7618 100000
rect 8022 99200 8078 100000
rect 8574 99200 8630 100000
rect 9034 99200 9090 100000
rect 9494 99200 9550 100000
rect 10046 99200 10102 100000
rect 10506 99200 10562 100000
rect 10966 99200 11022 100000
rect 11518 99200 11574 100000
rect 11978 99200 12034 100000
rect 12438 99200 12494 100000
rect 12990 99200 13046 100000
rect 13450 99200 13506 100000
rect 14002 99200 14058 100000
rect 14462 99200 14518 100000
rect 14922 99200 14978 100000
rect 15474 99200 15530 100000
rect 15934 99200 15990 100000
rect 16394 99200 16450 100000
rect 16946 99200 17002 100000
rect 17406 99200 17462 100000
rect 17866 99200 17922 100000
rect 18418 99200 18474 100000
rect 18878 99200 18934 100000
rect 19430 99200 19486 100000
rect 19890 99200 19946 100000
rect 20350 99200 20406 100000
rect 20902 99200 20958 100000
rect 21362 99200 21418 100000
rect 21822 99200 21878 100000
rect 22374 99200 22430 100000
rect 22834 99200 22890 100000
rect 23294 99200 23350 100000
rect 23846 99200 23902 100000
rect 24306 99200 24362 100000
rect 24766 99200 24822 100000
rect 25318 99200 25374 100000
rect 25778 99200 25834 100000
rect 26330 99200 26386 100000
rect 26790 99200 26846 100000
rect 27250 99200 27306 100000
rect 27802 99200 27858 100000
rect 28262 99200 28318 100000
rect 28722 99200 28778 100000
rect 29274 99200 29330 100000
rect 29734 99200 29790 100000
rect 30194 99200 30250 100000
rect 30746 99200 30802 100000
rect 31206 99200 31262 100000
rect 31666 99200 31722 100000
rect 32218 99200 32274 100000
rect 32678 99200 32734 100000
rect 33230 99200 33286 100000
rect 33690 99200 33746 100000
rect 34150 99200 34206 100000
rect 34702 99200 34758 100000
rect 35162 99200 35218 100000
rect 35622 99200 35678 100000
rect 36174 99200 36230 100000
rect 36634 99200 36690 100000
rect 37094 99200 37150 100000
rect 37646 99200 37702 100000
rect 38106 99200 38162 100000
rect 38658 99200 38714 100000
rect 39118 99200 39174 100000
rect 39578 99200 39634 100000
rect 40130 99200 40186 100000
rect 40590 99200 40646 100000
rect 41050 99200 41106 100000
rect 41602 99200 41658 100000
rect 42062 99200 42118 100000
rect 42522 99200 42578 100000
rect 43074 99200 43130 100000
rect 43534 99200 43590 100000
rect 43994 99200 44050 100000
rect 44546 99200 44602 100000
rect 45006 99200 45062 100000
rect 45558 99200 45614 100000
rect 46018 99200 46074 100000
rect 46478 99200 46534 100000
rect 47030 99200 47086 100000
rect 47490 99200 47546 100000
rect 47950 99200 48006 100000
rect 48502 99200 48558 100000
rect 48962 99200 49018 100000
rect 49422 99200 49478 100000
rect 49974 99200 50030 100000
rect 50434 99200 50490 100000
rect 50894 99200 50950 100000
rect 51446 99200 51502 100000
rect 51906 99200 51962 100000
rect 52458 99200 52514 100000
rect 52918 99200 52974 100000
rect 53378 99200 53434 100000
rect 53930 99200 53986 100000
rect 54390 99200 54446 100000
rect 54850 99200 54906 100000
rect 55402 99200 55458 100000
rect 55862 99200 55918 100000
rect 56322 99200 56378 100000
rect 56874 99200 56930 100000
rect 57334 99200 57390 100000
rect 57886 99200 57942 100000
rect 58346 99200 58402 100000
rect 58806 99200 58862 100000
rect 59358 99200 59414 100000
rect 59818 99200 59874 100000
rect 60278 99200 60334 100000
rect 60830 99200 60886 100000
rect 61290 99200 61346 100000
rect 61750 99200 61806 100000
rect 62302 99200 62358 100000
rect 62762 99200 62818 100000
rect 63222 99200 63278 100000
rect 63774 99200 63830 100000
rect 64234 99200 64290 100000
rect 64786 99200 64842 100000
rect 65246 99200 65302 100000
rect 65706 99200 65762 100000
rect 66258 99200 66314 100000
rect 66718 99200 66774 100000
rect 67178 99200 67234 100000
rect 67730 99200 67786 100000
rect 68190 99200 68246 100000
rect 68650 99200 68706 100000
rect 69202 99200 69258 100000
rect 69662 99200 69718 100000
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2226 0 2282 800
rect 2870 0 2926 800
rect 3514 0 3570 800
rect 4158 0 4214 800
rect 4802 0 4858 800
rect 5446 0 5502 800
rect 6090 0 6146 800
rect 6734 0 6790 800
rect 7378 0 7434 800
rect 8022 0 8078 800
rect 8666 0 8722 800
rect 9310 0 9366 800
rect 9954 0 10010 800
rect 10598 0 10654 800
rect 11242 0 11298 800
rect 11886 0 11942 800
rect 12530 0 12586 800
rect 13174 0 13230 800
rect 13818 0 13874 800
rect 14554 0 14610 800
rect 15198 0 15254 800
rect 15842 0 15898 800
rect 16486 0 16542 800
rect 17130 0 17186 800
rect 17774 0 17830 800
rect 18418 0 18474 800
rect 19062 0 19118 800
rect 19706 0 19762 800
rect 20350 0 20406 800
rect 20994 0 21050 800
rect 21638 0 21694 800
rect 22282 0 22338 800
rect 22926 0 22982 800
rect 23570 0 23626 800
rect 24214 0 24270 800
rect 24858 0 24914 800
rect 25502 0 25558 800
rect 26146 0 26202 800
rect 26790 0 26846 800
rect 27434 0 27490 800
rect 28078 0 28134 800
rect 28814 0 28870 800
rect 29458 0 29514 800
rect 30102 0 30158 800
rect 30746 0 30802 800
rect 31390 0 31446 800
rect 32034 0 32090 800
rect 32678 0 32734 800
rect 33322 0 33378 800
rect 33966 0 34022 800
rect 34610 0 34666 800
rect 35254 0 35310 800
rect 35898 0 35954 800
rect 36542 0 36598 800
rect 37186 0 37242 800
rect 37830 0 37886 800
rect 38474 0 38530 800
rect 39118 0 39174 800
rect 39762 0 39818 800
rect 40406 0 40462 800
rect 41050 0 41106 800
rect 41694 0 41750 800
rect 42430 0 42486 800
rect 43074 0 43130 800
rect 43718 0 43774 800
rect 44362 0 44418 800
rect 45006 0 45062 800
rect 45650 0 45706 800
rect 46294 0 46350 800
rect 46938 0 46994 800
rect 47582 0 47638 800
rect 48226 0 48282 800
rect 48870 0 48926 800
rect 49514 0 49570 800
rect 50158 0 50214 800
rect 50802 0 50858 800
rect 51446 0 51502 800
rect 52090 0 52146 800
rect 52734 0 52790 800
rect 53378 0 53434 800
rect 54022 0 54078 800
rect 54666 0 54722 800
rect 55310 0 55366 800
rect 55954 0 56010 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
<< obsm2 >>
rect 20 99144 146 99657
rect 314 99144 606 99657
rect 774 99144 1066 99657
rect 1234 99144 1618 99657
rect 1786 99144 2078 99657
rect 2246 99144 2538 99657
rect 2706 99144 3090 99657
rect 3258 99144 3550 99657
rect 3718 99144 4010 99657
rect 4178 99144 4562 99657
rect 4730 99144 5022 99657
rect 5190 99144 5482 99657
rect 5650 99144 6034 99657
rect 6202 99144 6494 99657
rect 6662 99144 7046 99657
rect 7214 99144 7506 99657
rect 7674 99144 7966 99657
rect 8134 99144 8518 99657
rect 8686 99144 8978 99657
rect 9146 99144 9438 99657
rect 9606 99144 9990 99657
rect 10158 99144 10450 99657
rect 10618 99144 10910 99657
rect 11078 99144 11462 99657
rect 11630 99144 11922 99657
rect 12090 99144 12382 99657
rect 12550 99144 12934 99657
rect 13102 99144 13394 99657
rect 13562 99144 13946 99657
rect 14114 99144 14406 99657
rect 14574 99144 14866 99657
rect 15034 99144 15418 99657
rect 15586 99144 15878 99657
rect 16046 99144 16338 99657
rect 16506 99144 16890 99657
rect 17058 99144 17350 99657
rect 17518 99144 17810 99657
rect 17978 99144 18362 99657
rect 18530 99144 18822 99657
rect 18990 99144 19374 99657
rect 19542 99144 19834 99657
rect 20002 99144 20294 99657
rect 20462 99144 20846 99657
rect 21014 99144 21306 99657
rect 21474 99144 21766 99657
rect 21934 99144 22318 99657
rect 22486 99144 22778 99657
rect 22946 99144 23238 99657
rect 23406 99144 23790 99657
rect 23958 99144 24250 99657
rect 24418 99144 24710 99657
rect 24878 99144 25262 99657
rect 25430 99144 25722 99657
rect 25890 99144 26274 99657
rect 26442 99144 26734 99657
rect 26902 99144 27194 99657
rect 27362 99144 27746 99657
rect 27914 99144 28206 99657
rect 28374 99144 28666 99657
rect 28834 99144 29218 99657
rect 29386 99144 29678 99657
rect 29846 99144 30138 99657
rect 30306 99144 30690 99657
rect 30858 99144 31150 99657
rect 31318 99144 31610 99657
rect 31778 99144 32162 99657
rect 32330 99144 32622 99657
rect 32790 99144 33174 99657
rect 33342 99144 33634 99657
rect 33802 99144 34094 99657
rect 34262 99144 34646 99657
rect 34814 99144 35106 99657
rect 35274 99144 35566 99657
rect 35734 99144 36118 99657
rect 36286 99144 36578 99657
rect 36746 99144 37038 99657
rect 37206 99144 37590 99657
rect 37758 99144 38050 99657
rect 38218 99144 38602 99657
rect 38770 99144 39062 99657
rect 39230 99144 39522 99657
rect 39690 99144 40074 99657
rect 40242 99144 40534 99657
rect 40702 99144 40994 99657
rect 41162 99144 41546 99657
rect 41714 99144 42006 99657
rect 42174 99144 42466 99657
rect 42634 99144 43018 99657
rect 43186 99144 43478 99657
rect 43646 99144 43938 99657
rect 44106 99144 44490 99657
rect 44658 99144 44950 99657
rect 45118 99144 45502 99657
rect 45670 99144 45962 99657
rect 46130 99144 46422 99657
rect 46590 99144 46974 99657
rect 47142 99144 47434 99657
rect 47602 99144 47894 99657
rect 48062 99144 48446 99657
rect 48614 99144 48906 99657
rect 49074 99144 49366 99657
rect 49534 99144 49918 99657
rect 50086 99144 50378 99657
rect 50546 99144 50838 99657
rect 51006 99144 51390 99657
rect 51558 99144 51850 99657
rect 52018 99144 52402 99657
rect 52570 99144 52862 99657
rect 53030 99144 53322 99657
rect 53490 99144 53874 99657
rect 54042 99144 54334 99657
rect 54502 99144 54794 99657
rect 54962 99144 55346 99657
rect 55514 99144 55806 99657
rect 55974 99144 56266 99657
rect 56434 99144 56818 99657
rect 56986 99144 57278 99657
rect 57446 99144 57830 99657
rect 57998 99144 58290 99657
rect 58458 99144 58750 99657
rect 58918 99144 59302 99657
rect 59470 99144 59762 99657
rect 59930 99144 60222 99657
rect 60390 99144 60774 99657
rect 60942 99144 61234 99657
rect 61402 99144 61694 99657
rect 61862 99144 62246 99657
rect 62414 99144 62706 99657
rect 62874 99144 63166 99657
rect 63334 99144 63718 99657
rect 63886 99144 64178 99657
rect 64346 99144 64730 99657
rect 64898 99144 65190 99657
rect 65358 99144 65650 99657
rect 65818 99144 66202 99657
rect 66370 99144 66662 99657
rect 66830 99144 67122 99657
rect 67290 99144 67674 99657
rect 67842 99144 68134 99657
rect 68302 99144 68594 99657
rect 68762 99144 69146 99657
rect 69314 99144 69606 99657
rect 69774 99144 69994 99657
rect 20 856 69994 99144
rect 20 31 238 856
rect 406 31 882 856
rect 1050 31 1526 856
rect 1694 31 2170 856
rect 2338 31 2814 856
rect 2982 31 3458 856
rect 3626 31 4102 856
rect 4270 31 4746 856
rect 4914 31 5390 856
rect 5558 31 6034 856
rect 6202 31 6678 856
rect 6846 31 7322 856
rect 7490 31 7966 856
rect 8134 31 8610 856
rect 8778 31 9254 856
rect 9422 31 9898 856
rect 10066 31 10542 856
rect 10710 31 11186 856
rect 11354 31 11830 856
rect 11998 31 12474 856
rect 12642 31 13118 856
rect 13286 31 13762 856
rect 13930 31 14498 856
rect 14666 31 15142 856
rect 15310 31 15786 856
rect 15954 31 16430 856
rect 16598 31 17074 856
rect 17242 31 17718 856
rect 17886 31 18362 856
rect 18530 31 19006 856
rect 19174 31 19650 856
rect 19818 31 20294 856
rect 20462 31 20938 856
rect 21106 31 21582 856
rect 21750 31 22226 856
rect 22394 31 22870 856
rect 23038 31 23514 856
rect 23682 31 24158 856
rect 24326 31 24802 856
rect 24970 31 25446 856
rect 25614 31 26090 856
rect 26258 31 26734 856
rect 26902 31 27378 856
rect 27546 31 28022 856
rect 28190 31 28758 856
rect 28926 31 29402 856
rect 29570 31 30046 856
rect 30214 31 30690 856
rect 30858 31 31334 856
rect 31502 31 31978 856
rect 32146 31 32622 856
rect 32790 31 33266 856
rect 33434 31 33910 856
rect 34078 31 34554 856
rect 34722 31 35198 856
rect 35366 31 35842 856
rect 36010 31 36486 856
rect 36654 31 37130 856
rect 37298 31 37774 856
rect 37942 31 38418 856
rect 38586 31 39062 856
rect 39230 31 39706 856
rect 39874 31 40350 856
rect 40518 31 40994 856
rect 41162 31 41638 856
rect 41806 31 42374 856
rect 42542 31 43018 856
rect 43186 31 43662 856
rect 43830 31 44306 856
rect 44474 31 44950 856
rect 45118 31 45594 856
rect 45762 31 46238 856
rect 46406 31 46882 856
rect 47050 31 47526 856
rect 47694 31 48170 856
rect 48338 31 48814 856
rect 48982 31 49458 856
rect 49626 31 50102 856
rect 50270 31 50746 856
rect 50914 31 51390 856
rect 51558 31 52034 856
rect 52202 31 52678 856
rect 52846 31 53322 856
rect 53490 31 53966 856
rect 54134 31 54610 856
rect 54778 31 55254 856
rect 55422 31 55898 856
rect 56066 31 56634 856
rect 56802 31 57278 856
rect 57446 31 57922 856
rect 58090 31 58566 856
rect 58734 31 59210 856
rect 59378 31 59854 856
rect 60022 31 60498 856
rect 60666 31 61142 856
rect 61310 31 61786 856
rect 61954 31 62430 856
rect 62598 31 63074 856
rect 63242 31 63718 856
rect 63886 31 64362 856
rect 64530 31 65006 856
rect 65174 31 65650 856
rect 65818 31 66294 856
rect 66462 31 66938 856
rect 67106 31 67582 856
rect 67750 31 68226 856
rect 68394 31 68870 856
rect 69038 31 69514 856
rect 69682 31 69994 856
<< metal3 >>
rect 69200 99560 70000 99680
rect 69200 99016 70000 99136
rect 69200 98472 70000 98592
rect 69200 97928 70000 98048
rect 69200 97384 70000 97504
rect 69200 96840 70000 96960
rect 69200 96296 70000 96416
rect 69200 95752 70000 95872
rect 69200 95208 70000 95328
rect 69200 94528 70000 94648
rect 69200 93984 70000 94104
rect 69200 93440 70000 93560
rect 69200 92896 70000 93016
rect 69200 92352 70000 92472
rect 69200 91808 70000 91928
rect 69200 91264 70000 91384
rect 69200 90720 70000 90840
rect 69200 90176 70000 90296
rect 69200 89496 70000 89616
rect 69200 88952 70000 89072
rect 69200 88408 70000 88528
rect 69200 87864 70000 87984
rect 69200 87320 70000 87440
rect 69200 86776 70000 86896
rect 69200 86232 70000 86352
rect 69200 85688 70000 85808
rect 69200 85144 70000 85264
rect 69200 84600 70000 84720
rect 69200 83920 70000 84040
rect 69200 83376 70000 83496
rect 69200 82832 70000 82952
rect 69200 82288 70000 82408
rect 69200 81744 70000 81864
rect 69200 81200 70000 81320
rect 69200 80656 70000 80776
rect 69200 80112 70000 80232
rect 69200 79568 70000 79688
rect 69200 78888 70000 79008
rect 69200 78344 70000 78464
rect 69200 77800 70000 77920
rect 69200 77256 70000 77376
rect 69200 76712 70000 76832
rect 69200 76168 70000 76288
rect 69200 75624 70000 75744
rect 69200 75080 70000 75200
rect 69200 74536 70000 74656
rect 69200 73992 70000 74112
rect 69200 73312 70000 73432
rect 69200 72768 70000 72888
rect 69200 72224 70000 72344
rect 69200 71680 70000 71800
rect 69200 71136 70000 71256
rect 69200 70592 70000 70712
rect 69200 70048 70000 70168
rect 69200 69504 70000 69624
rect 69200 68960 70000 69080
rect 69200 68280 70000 68400
rect 69200 67736 70000 67856
rect 69200 67192 70000 67312
rect 69200 66648 70000 66768
rect 69200 66104 70000 66224
rect 69200 65560 70000 65680
rect 69200 65016 70000 65136
rect 69200 64472 70000 64592
rect 69200 63928 70000 64048
rect 69200 63248 70000 63368
rect 69200 62704 70000 62824
rect 69200 62160 70000 62280
rect 69200 61616 70000 61736
rect 69200 61072 70000 61192
rect 69200 60528 70000 60648
rect 69200 59984 70000 60104
rect 69200 59440 70000 59560
rect 69200 58896 70000 59016
rect 69200 58352 70000 58472
rect 69200 57672 70000 57792
rect 69200 57128 70000 57248
rect 69200 56584 70000 56704
rect 69200 56040 70000 56160
rect 69200 55496 70000 55616
rect 69200 54952 70000 55072
rect 69200 54408 70000 54528
rect 69200 53864 70000 53984
rect 69200 53320 70000 53440
rect 69200 52640 70000 52760
rect 69200 52096 70000 52216
rect 69200 51552 70000 51672
rect 69200 51008 70000 51128
rect 69200 50464 70000 50584
rect 69200 49920 70000 50040
rect 69200 49376 70000 49496
rect 69200 48832 70000 48952
rect 69200 48288 70000 48408
rect 69200 47744 70000 47864
rect 69200 47064 70000 47184
rect 69200 46520 70000 46640
rect 69200 45976 70000 46096
rect 69200 45432 70000 45552
rect 69200 44888 70000 45008
rect 69200 44344 70000 44464
rect 69200 43800 70000 43920
rect 69200 43256 70000 43376
rect 69200 42712 70000 42832
rect 69200 42032 70000 42152
rect 69200 41488 70000 41608
rect 69200 40944 70000 41064
rect 69200 40400 70000 40520
rect 69200 39856 70000 39976
rect 69200 39312 70000 39432
rect 69200 38768 70000 38888
rect 69200 38224 70000 38344
rect 69200 37680 70000 37800
rect 69200 37136 70000 37256
rect 69200 36456 70000 36576
rect 69200 35912 70000 36032
rect 69200 35368 70000 35488
rect 69200 34824 70000 34944
rect 69200 34280 70000 34400
rect 69200 33736 70000 33856
rect 69200 33192 70000 33312
rect 69200 32648 70000 32768
rect 69200 32104 70000 32224
rect 69200 31424 70000 31544
rect 69200 30880 70000 31000
rect 69200 30336 70000 30456
rect 69200 29792 70000 29912
rect 69200 29248 70000 29368
rect 69200 28704 70000 28824
rect 69200 28160 70000 28280
rect 69200 27616 70000 27736
rect 69200 27072 70000 27192
rect 69200 26392 70000 26512
rect 69200 25848 70000 25968
rect 69200 25304 70000 25424
rect 69200 24760 70000 24880
rect 69200 24216 70000 24336
rect 69200 23672 70000 23792
rect 69200 23128 70000 23248
rect 69200 22584 70000 22704
rect 69200 22040 70000 22160
rect 69200 21496 70000 21616
rect 69200 20816 70000 20936
rect 69200 20272 70000 20392
rect 69200 19728 70000 19848
rect 69200 19184 70000 19304
rect 69200 18640 70000 18760
rect 69200 18096 70000 18216
rect 69200 17552 70000 17672
rect 69200 17008 70000 17128
rect 69200 16464 70000 16584
rect 69200 15784 70000 15904
rect 69200 15240 70000 15360
rect 69200 14696 70000 14816
rect 69200 14152 70000 14272
rect 69200 13608 70000 13728
rect 69200 13064 70000 13184
rect 69200 12520 70000 12640
rect 69200 11976 70000 12096
rect 69200 11432 70000 11552
rect 69200 10888 70000 11008
rect 69200 10208 70000 10328
rect 69200 9664 70000 9784
rect 69200 9120 70000 9240
rect 69200 8576 70000 8696
rect 69200 8032 70000 8152
rect 69200 7488 70000 7608
rect 69200 6944 70000 7064
rect 69200 6400 70000 6520
rect 69200 5856 70000 5976
rect 69200 5176 70000 5296
rect 69200 4632 70000 4752
rect 69200 4088 70000 4208
rect 69200 3544 70000 3664
rect 69200 3000 70000 3120
rect 69200 2456 70000 2576
rect 69200 1912 70000 2032
rect 69200 1368 70000 1488
rect 69200 824 70000 944
rect 69200 280 70000 400
<< obsm3 >>
rect 4210 99480 69120 99653
rect 4210 99216 69999 99480
rect 4210 98936 69120 99216
rect 4210 98672 69999 98936
rect 4210 98392 69120 98672
rect 4210 98128 69999 98392
rect 4210 97848 69120 98128
rect 4210 97584 69999 97848
rect 4210 97304 69120 97584
rect 4210 97040 69999 97304
rect 4210 96760 69120 97040
rect 4210 96496 69999 96760
rect 4210 96216 69120 96496
rect 4210 95952 69999 96216
rect 4210 95672 69120 95952
rect 4210 95408 69999 95672
rect 4210 95128 69120 95408
rect 4210 94728 69999 95128
rect 4210 94448 69120 94728
rect 4210 94184 69999 94448
rect 4210 93904 69120 94184
rect 4210 93640 69999 93904
rect 4210 93360 69120 93640
rect 4210 93096 69999 93360
rect 4210 92816 69120 93096
rect 4210 92552 69999 92816
rect 4210 92272 69120 92552
rect 4210 92008 69999 92272
rect 4210 91728 69120 92008
rect 4210 91464 69999 91728
rect 4210 91184 69120 91464
rect 4210 90920 69999 91184
rect 4210 90640 69120 90920
rect 4210 90376 69999 90640
rect 4210 90096 69120 90376
rect 4210 89696 69999 90096
rect 4210 89416 69120 89696
rect 4210 89152 69999 89416
rect 4210 88872 69120 89152
rect 4210 88608 69999 88872
rect 4210 88328 69120 88608
rect 4210 88064 69999 88328
rect 4210 87784 69120 88064
rect 4210 87520 69999 87784
rect 4210 87240 69120 87520
rect 4210 86976 69999 87240
rect 4210 86696 69120 86976
rect 4210 86432 69999 86696
rect 4210 86152 69120 86432
rect 4210 85888 69999 86152
rect 4210 85608 69120 85888
rect 4210 85344 69999 85608
rect 4210 85064 69120 85344
rect 4210 84800 69999 85064
rect 4210 84520 69120 84800
rect 4210 84120 69999 84520
rect 4210 83840 69120 84120
rect 4210 83576 69999 83840
rect 4210 83296 69120 83576
rect 4210 83032 69999 83296
rect 4210 82752 69120 83032
rect 4210 82488 69999 82752
rect 4210 82208 69120 82488
rect 4210 81944 69999 82208
rect 4210 81664 69120 81944
rect 4210 81400 69999 81664
rect 4210 81120 69120 81400
rect 4210 80856 69999 81120
rect 4210 80576 69120 80856
rect 4210 80312 69999 80576
rect 4210 80032 69120 80312
rect 4210 79768 69999 80032
rect 4210 79488 69120 79768
rect 4210 79088 69999 79488
rect 4210 78808 69120 79088
rect 4210 78544 69999 78808
rect 4210 78264 69120 78544
rect 4210 78000 69999 78264
rect 4210 77720 69120 78000
rect 4210 77456 69999 77720
rect 4210 77176 69120 77456
rect 4210 76912 69999 77176
rect 4210 76632 69120 76912
rect 4210 76368 69999 76632
rect 4210 76088 69120 76368
rect 4210 75824 69999 76088
rect 4210 75544 69120 75824
rect 4210 75280 69999 75544
rect 4210 75000 69120 75280
rect 4210 74736 69999 75000
rect 4210 74456 69120 74736
rect 4210 74192 69999 74456
rect 4210 73912 69120 74192
rect 4210 73512 69999 73912
rect 4210 73232 69120 73512
rect 4210 72968 69999 73232
rect 4210 72688 69120 72968
rect 4210 72424 69999 72688
rect 4210 72144 69120 72424
rect 4210 71880 69999 72144
rect 4210 71600 69120 71880
rect 4210 71336 69999 71600
rect 4210 71056 69120 71336
rect 4210 70792 69999 71056
rect 4210 70512 69120 70792
rect 4210 70248 69999 70512
rect 4210 69968 69120 70248
rect 4210 69704 69999 69968
rect 4210 69424 69120 69704
rect 4210 69160 69999 69424
rect 4210 68880 69120 69160
rect 4210 68480 69999 68880
rect 4210 68200 69120 68480
rect 4210 67936 69999 68200
rect 4210 67656 69120 67936
rect 4210 67392 69999 67656
rect 4210 67112 69120 67392
rect 4210 66848 69999 67112
rect 4210 66568 69120 66848
rect 4210 66304 69999 66568
rect 4210 66024 69120 66304
rect 4210 65760 69999 66024
rect 4210 65480 69120 65760
rect 4210 65216 69999 65480
rect 4210 64936 69120 65216
rect 4210 64672 69999 64936
rect 4210 64392 69120 64672
rect 4210 64128 69999 64392
rect 4210 63848 69120 64128
rect 4210 63448 69999 63848
rect 4210 63168 69120 63448
rect 4210 62904 69999 63168
rect 4210 62624 69120 62904
rect 4210 62360 69999 62624
rect 4210 62080 69120 62360
rect 4210 61816 69999 62080
rect 4210 61536 69120 61816
rect 4210 61272 69999 61536
rect 4210 60992 69120 61272
rect 4210 60728 69999 60992
rect 4210 60448 69120 60728
rect 4210 60184 69999 60448
rect 4210 59904 69120 60184
rect 4210 59640 69999 59904
rect 4210 59360 69120 59640
rect 4210 59096 69999 59360
rect 4210 58816 69120 59096
rect 4210 58552 69999 58816
rect 4210 58272 69120 58552
rect 4210 57872 69999 58272
rect 4210 57592 69120 57872
rect 4210 57328 69999 57592
rect 4210 57048 69120 57328
rect 4210 56784 69999 57048
rect 4210 56504 69120 56784
rect 4210 56240 69999 56504
rect 4210 55960 69120 56240
rect 4210 55696 69999 55960
rect 4210 55416 69120 55696
rect 4210 55152 69999 55416
rect 4210 54872 69120 55152
rect 4210 54608 69999 54872
rect 4210 54328 69120 54608
rect 4210 54064 69999 54328
rect 4210 53784 69120 54064
rect 4210 53520 69999 53784
rect 4210 53240 69120 53520
rect 4210 52840 69999 53240
rect 4210 52560 69120 52840
rect 4210 52296 69999 52560
rect 4210 52016 69120 52296
rect 4210 51752 69999 52016
rect 4210 51472 69120 51752
rect 4210 51208 69999 51472
rect 4210 50928 69120 51208
rect 4210 50664 69999 50928
rect 4210 50384 69120 50664
rect 4210 50120 69999 50384
rect 4210 49840 69120 50120
rect 4210 49576 69999 49840
rect 4210 49296 69120 49576
rect 4210 49032 69999 49296
rect 4210 48752 69120 49032
rect 4210 48488 69999 48752
rect 4210 48208 69120 48488
rect 4210 47944 69999 48208
rect 4210 47664 69120 47944
rect 4210 47264 69999 47664
rect 4210 46984 69120 47264
rect 4210 46720 69999 46984
rect 4210 46440 69120 46720
rect 4210 46176 69999 46440
rect 4210 45896 69120 46176
rect 4210 45632 69999 45896
rect 4210 45352 69120 45632
rect 4210 45088 69999 45352
rect 4210 44808 69120 45088
rect 4210 44544 69999 44808
rect 4210 44264 69120 44544
rect 4210 44000 69999 44264
rect 4210 43720 69120 44000
rect 4210 43456 69999 43720
rect 4210 43176 69120 43456
rect 4210 42912 69999 43176
rect 4210 42632 69120 42912
rect 4210 42232 69999 42632
rect 4210 41952 69120 42232
rect 4210 41688 69999 41952
rect 4210 41408 69120 41688
rect 4210 41144 69999 41408
rect 4210 40864 69120 41144
rect 4210 40600 69999 40864
rect 4210 40320 69120 40600
rect 4210 40056 69999 40320
rect 4210 39776 69120 40056
rect 4210 39512 69999 39776
rect 4210 39232 69120 39512
rect 4210 38968 69999 39232
rect 4210 38688 69120 38968
rect 4210 38424 69999 38688
rect 4210 38144 69120 38424
rect 4210 37880 69999 38144
rect 4210 37600 69120 37880
rect 4210 37336 69999 37600
rect 4210 37056 69120 37336
rect 4210 36656 69999 37056
rect 4210 36376 69120 36656
rect 4210 36112 69999 36376
rect 4210 35832 69120 36112
rect 4210 35568 69999 35832
rect 4210 35288 69120 35568
rect 4210 35024 69999 35288
rect 4210 34744 69120 35024
rect 4210 34480 69999 34744
rect 4210 34200 69120 34480
rect 4210 33936 69999 34200
rect 4210 33656 69120 33936
rect 4210 33392 69999 33656
rect 4210 33112 69120 33392
rect 4210 32848 69999 33112
rect 4210 32568 69120 32848
rect 4210 32304 69999 32568
rect 4210 32024 69120 32304
rect 4210 31624 69999 32024
rect 4210 31344 69120 31624
rect 4210 31080 69999 31344
rect 4210 30800 69120 31080
rect 4210 30536 69999 30800
rect 4210 30256 69120 30536
rect 4210 29992 69999 30256
rect 4210 29712 69120 29992
rect 4210 29448 69999 29712
rect 4210 29168 69120 29448
rect 4210 28904 69999 29168
rect 4210 28624 69120 28904
rect 4210 28360 69999 28624
rect 4210 28080 69120 28360
rect 4210 27816 69999 28080
rect 4210 27536 69120 27816
rect 4210 27272 69999 27536
rect 4210 26992 69120 27272
rect 4210 26592 69999 26992
rect 4210 26312 69120 26592
rect 4210 26048 69999 26312
rect 4210 25768 69120 26048
rect 4210 25504 69999 25768
rect 4210 25224 69120 25504
rect 4210 24960 69999 25224
rect 4210 24680 69120 24960
rect 4210 24416 69999 24680
rect 4210 24136 69120 24416
rect 4210 23872 69999 24136
rect 4210 23592 69120 23872
rect 4210 23328 69999 23592
rect 4210 23048 69120 23328
rect 4210 22784 69999 23048
rect 4210 22504 69120 22784
rect 4210 22240 69999 22504
rect 4210 21960 69120 22240
rect 4210 21696 69999 21960
rect 4210 21416 69120 21696
rect 4210 21016 69999 21416
rect 4210 20736 69120 21016
rect 4210 20472 69999 20736
rect 4210 20192 69120 20472
rect 4210 19928 69999 20192
rect 4210 19648 69120 19928
rect 4210 19384 69999 19648
rect 4210 19104 69120 19384
rect 4210 18840 69999 19104
rect 4210 18560 69120 18840
rect 4210 18296 69999 18560
rect 4210 18016 69120 18296
rect 4210 17752 69999 18016
rect 4210 17472 69120 17752
rect 4210 17208 69999 17472
rect 4210 16928 69120 17208
rect 4210 16664 69999 16928
rect 4210 16384 69120 16664
rect 4210 15984 69999 16384
rect 4210 15704 69120 15984
rect 4210 15440 69999 15704
rect 4210 15160 69120 15440
rect 4210 14896 69999 15160
rect 4210 14616 69120 14896
rect 4210 14352 69999 14616
rect 4210 14072 69120 14352
rect 4210 13808 69999 14072
rect 4210 13528 69120 13808
rect 4210 13264 69999 13528
rect 4210 12984 69120 13264
rect 4210 12720 69999 12984
rect 4210 12440 69120 12720
rect 4210 12176 69999 12440
rect 4210 11896 69120 12176
rect 4210 11632 69999 11896
rect 4210 11352 69120 11632
rect 4210 11088 69999 11352
rect 4210 10808 69120 11088
rect 4210 10408 69999 10808
rect 4210 10128 69120 10408
rect 4210 9864 69999 10128
rect 4210 9584 69120 9864
rect 4210 9320 69999 9584
rect 4210 9040 69120 9320
rect 4210 8776 69999 9040
rect 4210 8496 69120 8776
rect 4210 8232 69999 8496
rect 4210 7952 69120 8232
rect 4210 7688 69999 7952
rect 4210 7408 69120 7688
rect 4210 7144 69999 7408
rect 4210 6864 69120 7144
rect 4210 6600 69999 6864
rect 4210 6320 69120 6600
rect 4210 6056 69999 6320
rect 4210 5776 69120 6056
rect 4210 5376 69999 5776
rect 4210 5096 69120 5376
rect 4210 4832 69999 5096
rect 4210 4552 69120 4832
rect 4210 4288 69999 4552
rect 4210 4008 69120 4288
rect 4210 3744 69999 4008
rect 4210 3464 69120 3744
rect 4210 3200 69999 3464
rect 4210 2920 69120 3200
rect 4210 2656 69999 2920
rect 4210 2376 69120 2656
rect 4210 2112 69999 2376
rect 4210 1832 69120 2112
rect 4210 1568 69999 1832
rect 4210 1288 69120 1568
rect 4210 1024 69999 1288
rect 4210 744 69120 1024
rect 4210 480 69999 744
rect 4210 200 69120 480
rect 4210 35 69999 200
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
<< obsm4 >>
rect 34651 2048 34848 96525
rect 35328 2048 50208 96525
rect 50688 2048 65568 96525
rect 66048 2048 69861 96525
rect 34651 1531 69861 2048
<< labels >>
rlabel metal3 s 69200 5856 70000 5976 6 sram_addr0[0]
port 1 nsew signal output
rlabel metal3 s 69200 6400 70000 6520 6 sram_addr0[1]
port 2 nsew signal output
rlabel metal3 s 69200 6944 70000 7064 6 sram_addr0[2]
port 3 nsew signal output
rlabel metal3 s 69200 7488 70000 7608 6 sram_addr0[3]
port 4 nsew signal output
rlabel metal3 s 69200 8032 70000 8152 6 sram_addr0[4]
port 5 nsew signal output
rlabel metal3 s 69200 8576 70000 8696 6 sram_addr0[5]
port 6 nsew signal output
rlabel metal3 s 69200 9120 70000 9240 6 sram_addr0[6]
port 7 nsew signal output
rlabel metal3 s 69200 9664 70000 9784 6 sram_addr0[7]
port 8 nsew signal output
rlabel metal3 s 69200 10208 70000 10328 6 sram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 2594 99200 2650 100000 6 sram_addr1[0]
port 10 nsew signal output
rlabel metal2 s 3146 99200 3202 100000 6 sram_addr1[1]
port 11 nsew signal output
rlabel metal2 s 3606 99200 3662 100000 6 sram_addr1[2]
port 12 nsew signal output
rlabel metal2 s 4066 99200 4122 100000 6 sram_addr1[3]
port 13 nsew signal output
rlabel metal2 s 4618 99200 4674 100000 6 sram_addr1[4]
port 14 nsew signal output
rlabel metal2 s 5078 99200 5134 100000 6 sram_addr1[5]
port 15 nsew signal output
rlabel metal2 s 5538 99200 5594 100000 6 sram_addr1[6]
port 16 nsew signal output
rlabel metal2 s 6090 99200 6146 100000 6 sram_addr1[7]
port 17 nsew signal output
rlabel metal2 s 6550 99200 6606 100000 6 sram_addr1[8]
port 18 nsew signal output
rlabel metal3 s 69200 280 70000 400 6 sram_clk0
port 19 nsew signal output
rlabel metal2 s 202 99200 258 100000 6 sram_clk1
port 20 nsew signal output
rlabel metal3 s 69200 824 70000 944 6 sram_csb0[0]
port 21 nsew signal output
rlabel metal3 s 69200 1368 70000 1488 6 sram_csb0[1]
port 22 nsew signal output
rlabel metal3 s 69200 1912 70000 2032 6 sram_csb0[2]
port 23 nsew signal output
rlabel metal3 s 69200 2456 70000 2576 6 sram_csb0[3]
port 24 nsew signal output
rlabel metal2 s 662 99200 718 100000 6 sram_csb1[0]
port 25 nsew signal output
rlabel metal2 s 1122 99200 1178 100000 6 sram_csb1[1]
port 26 nsew signal output
rlabel metal2 s 1674 99200 1730 100000 6 sram_csb1[2]
port 27 nsew signal output
rlabel metal2 s 2134 99200 2190 100000 6 sram_csb1[3]
port 28 nsew signal output
rlabel metal3 s 69200 10888 70000 11008 6 sram_din0[0]
port 29 nsew signal output
rlabel metal3 s 69200 16464 70000 16584 6 sram_din0[10]
port 30 nsew signal output
rlabel metal3 s 69200 17008 70000 17128 6 sram_din0[11]
port 31 nsew signal output
rlabel metal3 s 69200 17552 70000 17672 6 sram_din0[12]
port 32 nsew signal output
rlabel metal3 s 69200 18096 70000 18216 6 sram_din0[13]
port 33 nsew signal output
rlabel metal3 s 69200 18640 70000 18760 6 sram_din0[14]
port 34 nsew signal output
rlabel metal3 s 69200 19184 70000 19304 6 sram_din0[15]
port 35 nsew signal output
rlabel metal3 s 69200 19728 70000 19848 6 sram_din0[16]
port 36 nsew signal output
rlabel metal3 s 69200 20272 70000 20392 6 sram_din0[17]
port 37 nsew signal output
rlabel metal3 s 69200 20816 70000 20936 6 sram_din0[18]
port 38 nsew signal output
rlabel metal3 s 69200 21496 70000 21616 6 sram_din0[19]
port 39 nsew signal output
rlabel metal3 s 69200 11432 70000 11552 6 sram_din0[1]
port 40 nsew signal output
rlabel metal3 s 69200 22040 70000 22160 6 sram_din0[20]
port 41 nsew signal output
rlabel metal3 s 69200 22584 70000 22704 6 sram_din0[21]
port 42 nsew signal output
rlabel metal3 s 69200 23128 70000 23248 6 sram_din0[22]
port 43 nsew signal output
rlabel metal3 s 69200 23672 70000 23792 6 sram_din0[23]
port 44 nsew signal output
rlabel metal3 s 69200 24216 70000 24336 6 sram_din0[24]
port 45 nsew signal output
rlabel metal3 s 69200 24760 70000 24880 6 sram_din0[25]
port 46 nsew signal output
rlabel metal3 s 69200 25304 70000 25424 6 sram_din0[26]
port 47 nsew signal output
rlabel metal3 s 69200 25848 70000 25968 6 sram_din0[27]
port 48 nsew signal output
rlabel metal3 s 69200 26392 70000 26512 6 sram_din0[28]
port 49 nsew signal output
rlabel metal3 s 69200 27072 70000 27192 6 sram_din0[29]
port 50 nsew signal output
rlabel metal3 s 69200 11976 70000 12096 6 sram_din0[2]
port 51 nsew signal output
rlabel metal3 s 69200 27616 70000 27736 6 sram_din0[30]
port 52 nsew signal output
rlabel metal3 s 69200 28160 70000 28280 6 sram_din0[31]
port 53 nsew signal output
rlabel metal3 s 69200 12520 70000 12640 6 sram_din0[3]
port 54 nsew signal output
rlabel metal3 s 69200 13064 70000 13184 6 sram_din0[4]
port 55 nsew signal output
rlabel metal3 s 69200 13608 70000 13728 6 sram_din0[5]
port 56 nsew signal output
rlabel metal3 s 69200 14152 70000 14272 6 sram_din0[6]
port 57 nsew signal output
rlabel metal3 s 69200 14696 70000 14816 6 sram_din0[7]
port 58 nsew signal output
rlabel metal3 s 69200 15240 70000 15360 6 sram_din0[8]
port 59 nsew signal output
rlabel metal3 s 69200 15784 70000 15904 6 sram_din0[9]
port 60 nsew signal output
rlabel metal3 s 69200 28704 70000 28824 6 sram_dout0[0]
port 61 nsew signal input
rlabel metal3 s 69200 84600 70000 84720 6 sram_dout0[100]
port 62 nsew signal input
rlabel metal3 s 69200 85144 70000 85264 6 sram_dout0[101]
port 63 nsew signal input
rlabel metal3 s 69200 85688 70000 85808 6 sram_dout0[102]
port 64 nsew signal input
rlabel metal3 s 69200 86232 70000 86352 6 sram_dout0[103]
port 65 nsew signal input
rlabel metal3 s 69200 86776 70000 86896 6 sram_dout0[104]
port 66 nsew signal input
rlabel metal3 s 69200 87320 70000 87440 6 sram_dout0[105]
port 67 nsew signal input
rlabel metal3 s 69200 87864 70000 87984 6 sram_dout0[106]
port 68 nsew signal input
rlabel metal3 s 69200 88408 70000 88528 6 sram_dout0[107]
port 69 nsew signal input
rlabel metal3 s 69200 88952 70000 89072 6 sram_dout0[108]
port 70 nsew signal input
rlabel metal3 s 69200 89496 70000 89616 6 sram_dout0[109]
port 71 nsew signal input
rlabel metal3 s 69200 34280 70000 34400 6 sram_dout0[10]
port 72 nsew signal input
rlabel metal3 s 69200 90176 70000 90296 6 sram_dout0[110]
port 73 nsew signal input
rlabel metal3 s 69200 90720 70000 90840 6 sram_dout0[111]
port 74 nsew signal input
rlabel metal3 s 69200 91264 70000 91384 6 sram_dout0[112]
port 75 nsew signal input
rlabel metal3 s 69200 91808 70000 91928 6 sram_dout0[113]
port 76 nsew signal input
rlabel metal3 s 69200 92352 70000 92472 6 sram_dout0[114]
port 77 nsew signal input
rlabel metal3 s 69200 92896 70000 93016 6 sram_dout0[115]
port 78 nsew signal input
rlabel metal3 s 69200 93440 70000 93560 6 sram_dout0[116]
port 79 nsew signal input
rlabel metal3 s 69200 93984 70000 94104 6 sram_dout0[117]
port 80 nsew signal input
rlabel metal3 s 69200 94528 70000 94648 6 sram_dout0[118]
port 81 nsew signal input
rlabel metal3 s 69200 95208 70000 95328 6 sram_dout0[119]
port 82 nsew signal input
rlabel metal3 s 69200 34824 70000 34944 6 sram_dout0[11]
port 83 nsew signal input
rlabel metal3 s 69200 95752 70000 95872 6 sram_dout0[120]
port 84 nsew signal input
rlabel metal3 s 69200 96296 70000 96416 6 sram_dout0[121]
port 85 nsew signal input
rlabel metal3 s 69200 96840 70000 96960 6 sram_dout0[122]
port 86 nsew signal input
rlabel metal3 s 69200 97384 70000 97504 6 sram_dout0[123]
port 87 nsew signal input
rlabel metal3 s 69200 97928 70000 98048 6 sram_dout0[124]
port 88 nsew signal input
rlabel metal3 s 69200 98472 70000 98592 6 sram_dout0[125]
port 89 nsew signal input
rlabel metal3 s 69200 99016 70000 99136 6 sram_dout0[126]
port 90 nsew signal input
rlabel metal3 s 69200 99560 70000 99680 6 sram_dout0[127]
port 91 nsew signal input
rlabel metal3 s 69200 35368 70000 35488 6 sram_dout0[12]
port 92 nsew signal input
rlabel metal3 s 69200 35912 70000 36032 6 sram_dout0[13]
port 93 nsew signal input
rlabel metal3 s 69200 36456 70000 36576 6 sram_dout0[14]
port 94 nsew signal input
rlabel metal3 s 69200 37136 70000 37256 6 sram_dout0[15]
port 95 nsew signal input
rlabel metal3 s 69200 37680 70000 37800 6 sram_dout0[16]
port 96 nsew signal input
rlabel metal3 s 69200 38224 70000 38344 6 sram_dout0[17]
port 97 nsew signal input
rlabel metal3 s 69200 38768 70000 38888 6 sram_dout0[18]
port 98 nsew signal input
rlabel metal3 s 69200 39312 70000 39432 6 sram_dout0[19]
port 99 nsew signal input
rlabel metal3 s 69200 29248 70000 29368 6 sram_dout0[1]
port 100 nsew signal input
rlabel metal3 s 69200 39856 70000 39976 6 sram_dout0[20]
port 101 nsew signal input
rlabel metal3 s 69200 40400 70000 40520 6 sram_dout0[21]
port 102 nsew signal input
rlabel metal3 s 69200 40944 70000 41064 6 sram_dout0[22]
port 103 nsew signal input
rlabel metal3 s 69200 41488 70000 41608 6 sram_dout0[23]
port 104 nsew signal input
rlabel metal3 s 69200 42032 70000 42152 6 sram_dout0[24]
port 105 nsew signal input
rlabel metal3 s 69200 42712 70000 42832 6 sram_dout0[25]
port 106 nsew signal input
rlabel metal3 s 69200 43256 70000 43376 6 sram_dout0[26]
port 107 nsew signal input
rlabel metal3 s 69200 43800 70000 43920 6 sram_dout0[27]
port 108 nsew signal input
rlabel metal3 s 69200 44344 70000 44464 6 sram_dout0[28]
port 109 nsew signal input
rlabel metal3 s 69200 44888 70000 45008 6 sram_dout0[29]
port 110 nsew signal input
rlabel metal3 s 69200 29792 70000 29912 6 sram_dout0[2]
port 111 nsew signal input
rlabel metal3 s 69200 45432 70000 45552 6 sram_dout0[30]
port 112 nsew signal input
rlabel metal3 s 69200 45976 70000 46096 6 sram_dout0[31]
port 113 nsew signal input
rlabel metal3 s 69200 46520 70000 46640 6 sram_dout0[32]
port 114 nsew signal input
rlabel metal3 s 69200 47064 70000 47184 6 sram_dout0[33]
port 115 nsew signal input
rlabel metal3 s 69200 47744 70000 47864 6 sram_dout0[34]
port 116 nsew signal input
rlabel metal3 s 69200 48288 70000 48408 6 sram_dout0[35]
port 117 nsew signal input
rlabel metal3 s 69200 48832 70000 48952 6 sram_dout0[36]
port 118 nsew signal input
rlabel metal3 s 69200 49376 70000 49496 6 sram_dout0[37]
port 119 nsew signal input
rlabel metal3 s 69200 49920 70000 50040 6 sram_dout0[38]
port 120 nsew signal input
rlabel metal3 s 69200 50464 70000 50584 6 sram_dout0[39]
port 121 nsew signal input
rlabel metal3 s 69200 30336 70000 30456 6 sram_dout0[3]
port 122 nsew signal input
rlabel metal3 s 69200 51008 70000 51128 6 sram_dout0[40]
port 123 nsew signal input
rlabel metal3 s 69200 51552 70000 51672 6 sram_dout0[41]
port 124 nsew signal input
rlabel metal3 s 69200 52096 70000 52216 6 sram_dout0[42]
port 125 nsew signal input
rlabel metal3 s 69200 52640 70000 52760 6 sram_dout0[43]
port 126 nsew signal input
rlabel metal3 s 69200 53320 70000 53440 6 sram_dout0[44]
port 127 nsew signal input
rlabel metal3 s 69200 53864 70000 53984 6 sram_dout0[45]
port 128 nsew signal input
rlabel metal3 s 69200 54408 70000 54528 6 sram_dout0[46]
port 129 nsew signal input
rlabel metal3 s 69200 54952 70000 55072 6 sram_dout0[47]
port 130 nsew signal input
rlabel metal3 s 69200 55496 70000 55616 6 sram_dout0[48]
port 131 nsew signal input
rlabel metal3 s 69200 56040 70000 56160 6 sram_dout0[49]
port 132 nsew signal input
rlabel metal3 s 69200 30880 70000 31000 6 sram_dout0[4]
port 133 nsew signal input
rlabel metal3 s 69200 56584 70000 56704 6 sram_dout0[50]
port 134 nsew signal input
rlabel metal3 s 69200 57128 70000 57248 6 sram_dout0[51]
port 135 nsew signal input
rlabel metal3 s 69200 57672 70000 57792 6 sram_dout0[52]
port 136 nsew signal input
rlabel metal3 s 69200 58352 70000 58472 6 sram_dout0[53]
port 137 nsew signal input
rlabel metal3 s 69200 58896 70000 59016 6 sram_dout0[54]
port 138 nsew signal input
rlabel metal3 s 69200 59440 70000 59560 6 sram_dout0[55]
port 139 nsew signal input
rlabel metal3 s 69200 59984 70000 60104 6 sram_dout0[56]
port 140 nsew signal input
rlabel metal3 s 69200 60528 70000 60648 6 sram_dout0[57]
port 141 nsew signal input
rlabel metal3 s 69200 61072 70000 61192 6 sram_dout0[58]
port 142 nsew signal input
rlabel metal3 s 69200 61616 70000 61736 6 sram_dout0[59]
port 143 nsew signal input
rlabel metal3 s 69200 31424 70000 31544 6 sram_dout0[5]
port 144 nsew signal input
rlabel metal3 s 69200 62160 70000 62280 6 sram_dout0[60]
port 145 nsew signal input
rlabel metal3 s 69200 62704 70000 62824 6 sram_dout0[61]
port 146 nsew signal input
rlabel metal3 s 69200 63248 70000 63368 6 sram_dout0[62]
port 147 nsew signal input
rlabel metal3 s 69200 63928 70000 64048 6 sram_dout0[63]
port 148 nsew signal input
rlabel metal3 s 69200 64472 70000 64592 6 sram_dout0[64]
port 149 nsew signal input
rlabel metal3 s 69200 65016 70000 65136 6 sram_dout0[65]
port 150 nsew signal input
rlabel metal3 s 69200 65560 70000 65680 6 sram_dout0[66]
port 151 nsew signal input
rlabel metal3 s 69200 66104 70000 66224 6 sram_dout0[67]
port 152 nsew signal input
rlabel metal3 s 69200 66648 70000 66768 6 sram_dout0[68]
port 153 nsew signal input
rlabel metal3 s 69200 67192 70000 67312 6 sram_dout0[69]
port 154 nsew signal input
rlabel metal3 s 69200 32104 70000 32224 6 sram_dout0[6]
port 155 nsew signal input
rlabel metal3 s 69200 67736 70000 67856 6 sram_dout0[70]
port 156 nsew signal input
rlabel metal3 s 69200 68280 70000 68400 6 sram_dout0[71]
port 157 nsew signal input
rlabel metal3 s 69200 68960 70000 69080 6 sram_dout0[72]
port 158 nsew signal input
rlabel metal3 s 69200 69504 70000 69624 6 sram_dout0[73]
port 159 nsew signal input
rlabel metal3 s 69200 70048 70000 70168 6 sram_dout0[74]
port 160 nsew signal input
rlabel metal3 s 69200 70592 70000 70712 6 sram_dout0[75]
port 161 nsew signal input
rlabel metal3 s 69200 71136 70000 71256 6 sram_dout0[76]
port 162 nsew signal input
rlabel metal3 s 69200 71680 70000 71800 6 sram_dout0[77]
port 163 nsew signal input
rlabel metal3 s 69200 72224 70000 72344 6 sram_dout0[78]
port 164 nsew signal input
rlabel metal3 s 69200 72768 70000 72888 6 sram_dout0[79]
port 165 nsew signal input
rlabel metal3 s 69200 32648 70000 32768 6 sram_dout0[7]
port 166 nsew signal input
rlabel metal3 s 69200 73312 70000 73432 6 sram_dout0[80]
port 167 nsew signal input
rlabel metal3 s 69200 73992 70000 74112 6 sram_dout0[81]
port 168 nsew signal input
rlabel metal3 s 69200 74536 70000 74656 6 sram_dout0[82]
port 169 nsew signal input
rlabel metal3 s 69200 75080 70000 75200 6 sram_dout0[83]
port 170 nsew signal input
rlabel metal3 s 69200 75624 70000 75744 6 sram_dout0[84]
port 171 nsew signal input
rlabel metal3 s 69200 76168 70000 76288 6 sram_dout0[85]
port 172 nsew signal input
rlabel metal3 s 69200 76712 70000 76832 6 sram_dout0[86]
port 173 nsew signal input
rlabel metal3 s 69200 77256 70000 77376 6 sram_dout0[87]
port 174 nsew signal input
rlabel metal3 s 69200 77800 70000 77920 6 sram_dout0[88]
port 175 nsew signal input
rlabel metal3 s 69200 78344 70000 78464 6 sram_dout0[89]
port 176 nsew signal input
rlabel metal3 s 69200 33192 70000 33312 6 sram_dout0[8]
port 177 nsew signal input
rlabel metal3 s 69200 78888 70000 79008 6 sram_dout0[90]
port 178 nsew signal input
rlabel metal3 s 69200 79568 70000 79688 6 sram_dout0[91]
port 179 nsew signal input
rlabel metal3 s 69200 80112 70000 80232 6 sram_dout0[92]
port 180 nsew signal input
rlabel metal3 s 69200 80656 70000 80776 6 sram_dout0[93]
port 181 nsew signal input
rlabel metal3 s 69200 81200 70000 81320 6 sram_dout0[94]
port 182 nsew signal input
rlabel metal3 s 69200 81744 70000 81864 6 sram_dout0[95]
port 183 nsew signal input
rlabel metal3 s 69200 82288 70000 82408 6 sram_dout0[96]
port 184 nsew signal input
rlabel metal3 s 69200 82832 70000 82952 6 sram_dout0[97]
port 185 nsew signal input
rlabel metal3 s 69200 83376 70000 83496 6 sram_dout0[98]
port 186 nsew signal input
rlabel metal3 s 69200 83920 70000 84040 6 sram_dout0[99]
port 187 nsew signal input
rlabel metal3 s 69200 33736 70000 33856 6 sram_dout0[9]
port 188 nsew signal input
rlabel metal2 s 7102 99200 7158 100000 6 sram_dout1[0]
port 189 nsew signal input
rlabel metal2 s 56322 99200 56378 100000 6 sram_dout1[100]
port 190 nsew signal input
rlabel metal2 s 56874 99200 56930 100000 6 sram_dout1[101]
port 191 nsew signal input
rlabel metal2 s 57334 99200 57390 100000 6 sram_dout1[102]
port 192 nsew signal input
rlabel metal2 s 57886 99200 57942 100000 6 sram_dout1[103]
port 193 nsew signal input
rlabel metal2 s 58346 99200 58402 100000 6 sram_dout1[104]
port 194 nsew signal input
rlabel metal2 s 58806 99200 58862 100000 6 sram_dout1[105]
port 195 nsew signal input
rlabel metal2 s 59358 99200 59414 100000 6 sram_dout1[106]
port 196 nsew signal input
rlabel metal2 s 59818 99200 59874 100000 6 sram_dout1[107]
port 197 nsew signal input
rlabel metal2 s 60278 99200 60334 100000 6 sram_dout1[108]
port 198 nsew signal input
rlabel metal2 s 60830 99200 60886 100000 6 sram_dout1[109]
port 199 nsew signal input
rlabel metal2 s 11978 99200 12034 100000 6 sram_dout1[10]
port 200 nsew signal input
rlabel metal2 s 61290 99200 61346 100000 6 sram_dout1[110]
port 201 nsew signal input
rlabel metal2 s 61750 99200 61806 100000 6 sram_dout1[111]
port 202 nsew signal input
rlabel metal2 s 62302 99200 62358 100000 6 sram_dout1[112]
port 203 nsew signal input
rlabel metal2 s 62762 99200 62818 100000 6 sram_dout1[113]
port 204 nsew signal input
rlabel metal2 s 63222 99200 63278 100000 6 sram_dout1[114]
port 205 nsew signal input
rlabel metal2 s 63774 99200 63830 100000 6 sram_dout1[115]
port 206 nsew signal input
rlabel metal2 s 64234 99200 64290 100000 6 sram_dout1[116]
port 207 nsew signal input
rlabel metal2 s 64786 99200 64842 100000 6 sram_dout1[117]
port 208 nsew signal input
rlabel metal2 s 65246 99200 65302 100000 6 sram_dout1[118]
port 209 nsew signal input
rlabel metal2 s 65706 99200 65762 100000 6 sram_dout1[119]
port 210 nsew signal input
rlabel metal2 s 12438 99200 12494 100000 6 sram_dout1[11]
port 211 nsew signal input
rlabel metal2 s 66258 99200 66314 100000 6 sram_dout1[120]
port 212 nsew signal input
rlabel metal2 s 66718 99200 66774 100000 6 sram_dout1[121]
port 213 nsew signal input
rlabel metal2 s 67178 99200 67234 100000 6 sram_dout1[122]
port 214 nsew signal input
rlabel metal2 s 67730 99200 67786 100000 6 sram_dout1[123]
port 215 nsew signal input
rlabel metal2 s 68190 99200 68246 100000 6 sram_dout1[124]
port 216 nsew signal input
rlabel metal2 s 68650 99200 68706 100000 6 sram_dout1[125]
port 217 nsew signal input
rlabel metal2 s 69202 99200 69258 100000 6 sram_dout1[126]
port 218 nsew signal input
rlabel metal2 s 69662 99200 69718 100000 6 sram_dout1[127]
port 219 nsew signal input
rlabel metal2 s 12990 99200 13046 100000 6 sram_dout1[12]
port 220 nsew signal input
rlabel metal2 s 13450 99200 13506 100000 6 sram_dout1[13]
port 221 nsew signal input
rlabel metal2 s 14002 99200 14058 100000 6 sram_dout1[14]
port 222 nsew signal input
rlabel metal2 s 14462 99200 14518 100000 6 sram_dout1[15]
port 223 nsew signal input
rlabel metal2 s 14922 99200 14978 100000 6 sram_dout1[16]
port 224 nsew signal input
rlabel metal2 s 15474 99200 15530 100000 6 sram_dout1[17]
port 225 nsew signal input
rlabel metal2 s 15934 99200 15990 100000 6 sram_dout1[18]
port 226 nsew signal input
rlabel metal2 s 16394 99200 16450 100000 6 sram_dout1[19]
port 227 nsew signal input
rlabel metal2 s 7562 99200 7618 100000 6 sram_dout1[1]
port 228 nsew signal input
rlabel metal2 s 16946 99200 17002 100000 6 sram_dout1[20]
port 229 nsew signal input
rlabel metal2 s 17406 99200 17462 100000 6 sram_dout1[21]
port 230 nsew signal input
rlabel metal2 s 17866 99200 17922 100000 6 sram_dout1[22]
port 231 nsew signal input
rlabel metal2 s 18418 99200 18474 100000 6 sram_dout1[23]
port 232 nsew signal input
rlabel metal2 s 18878 99200 18934 100000 6 sram_dout1[24]
port 233 nsew signal input
rlabel metal2 s 19430 99200 19486 100000 6 sram_dout1[25]
port 234 nsew signal input
rlabel metal2 s 19890 99200 19946 100000 6 sram_dout1[26]
port 235 nsew signal input
rlabel metal2 s 20350 99200 20406 100000 6 sram_dout1[27]
port 236 nsew signal input
rlabel metal2 s 20902 99200 20958 100000 6 sram_dout1[28]
port 237 nsew signal input
rlabel metal2 s 21362 99200 21418 100000 6 sram_dout1[29]
port 238 nsew signal input
rlabel metal2 s 8022 99200 8078 100000 6 sram_dout1[2]
port 239 nsew signal input
rlabel metal2 s 21822 99200 21878 100000 6 sram_dout1[30]
port 240 nsew signal input
rlabel metal2 s 22374 99200 22430 100000 6 sram_dout1[31]
port 241 nsew signal input
rlabel metal2 s 22834 99200 22890 100000 6 sram_dout1[32]
port 242 nsew signal input
rlabel metal2 s 23294 99200 23350 100000 6 sram_dout1[33]
port 243 nsew signal input
rlabel metal2 s 23846 99200 23902 100000 6 sram_dout1[34]
port 244 nsew signal input
rlabel metal2 s 24306 99200 24362 100000 6 sram_dout1[35]
port 245 nsew signal input
rlabel metal2 s 24766 99200 24822 100000 6 sram_dout1[36]
port 246 nsew signal input
rlabel metal2 s 25318 99200 25374 100000 6 sram_dout1[37]
port 247 nsew signal input
rlabel metal2 s 25778 99200 25834 100000 6 sram_dout1[38]
port 248 nsew signal input
rlabel metal2 s 26330 99200 26386 100000 6 sram_dout1[39]
port 249 nsew signal input
rlabel metal2 s 8574 99200 8630 100000 6 sram_dout1[3]
port 250 nsew signal input
rlabel metal2 s 26790 99200 26846 100000 6 sram_dout1[40]
port 251 nsew signal input
rlabel metal2 s 27250 99200 27306 100000 6 sram_dout1[41]
port 252 nsew signal input
rlabel metal2 s 27802 99200 27858 100000 6 sram_dout1[42]
port 253 nsew signal input
rlabel metal2 s 28262 99200 28318 100000 6 sram_dout1[43]
port 254 nsew signal input
rlabel metal2 s 28722 99200 28778 100000 6 sram_dout1[44]
port 255 nsew signal input
rlabel metal2 s 29274 99200 29330 100000 6 sram_dout1[45]
port 256 nsew signal input
rlabel metal2 s 29734 99200 29790 100000 6 sram_dout1[46]
port 257 nsew signal input
rlabel metal2 s 30194 99200 30250 100000 6 sram_dout1[47]
port 258 nsew signal input
rlabel metal2 s 30746 99200 30802 100000 6 sram_dout1[48]
port 259 nsew signal input
rlabel metal2 s 31206 99200 31262 100000 6 sram_dout1[49]
port 260 nsew signal input
rlabel metal2 s 9034 99200 9090 100000 6 sram_dout1[4]
port 261 nsew signal input
rlabel metal2 s 31666 99200 31722 100000 6 sram_dout1[50]
port 262 nsew signal input
rlabel metal2 s 32218 99200 32274 100000 6 sram_dout1[51]
port 263 nsew signal input
rlabel metal2 s 32678 99200 32734 100000 6 sram_dout1[52]
port 264 nsew signal input
rlabel metal2 s 33230 99200 33286 100000 6 sram_dout1[53]
port 265 nsew signal input
rlabel metal2 s 33690 99200 33746 100000 6 sram_dout1[54]
port 266 nsew signal input
rlabel metal2 s 34150 99200 34206 100000 6 sram_dout1[55]
port 267 nsew signal input
rlabel metal2 s 34702 99200 34758 100000 6 sram_dout1[56]
port 268 nsew signal input
rlabel metal2 s 35162 99200 35218 100000 6 sram_dout1[57]
port 269 nsew signal input
rlabel metal2 s 35622 99200 35678 100000 6 sram_dout1[58]
port 270 nsew signal input
rlabel metal2 s 36174 99200 36230 100000 6 sram_dout1[59]
port 271 nsew signal input
rlabel metal2 s 9494 99200 9550 100000 6 sram_dout1[5]
port 272 nsew signal input
rlabel metal2 s 36634 99200 36690 100000 6 sram_dout1[60]
port 273 nsew signal input
rlabel metal2 s 37094 99200 37150 100000 6 sram_dout1[61]
port 274 nsew signal input
rlabel metal2 s 37646 99200 37702 100000 6 sram_dout1[62]
port 275 nsew signal input
rlabel metal2 s 38106 99200 38162 100000 6 sram_dout1[63]
port 276 nsew signal input
rlabel metal2 s 38658 99200 38714 100000 6 sram_dout1[64]
port 277 nsew signal input
rlabel metal2 s 39118 99200 39174 100000 6 sram_dout1[65]
port 278 nsew signal input
rlabel metal2 s 39578 99200 39634 100000 6 sram_dout1[66]
port 279 nsew signal input
rlabel metal2 s 40130 99200 40186 100000 6 sram_dout1[67]
port 280 nsew signal input
rlabel metal2 s 40590 99200 40646 100000 6 sram_dout1[68]
port 281 nsew signal input
rlabel metal2 s 41050 99200 41106 100000 6 sram_dout1[69]
port 282 nsew signal input
rlabel metal2 s 10046 99200 10102 100000 6 sram_dout1[6]
port 283 nsew signal input
rlabel metal2 s 41602 99200 41658 100000 6 sram_dout1[70]
port 284 nsew signal input
rlabel metal2 s 42062 99200 42118 100000 6 sram_dout1[71]
port 285 nsew signal input
rlabel metal2 s 42522 99200 42578 100000 6 sram_dout1[72]
port 286 nsew signal input
rlabel metal2 s 43074 99200 43130 100000 6 sram_dout1[73]
port 287 nsew signal input
rlabel metal2 s 43534 99200 43590 100000 6 sram_dout1[74]
port 288 nsew signal input
rlabel metal2 s 43994 99200 44050 100000 6 sram_dout1[75]
port 289 nsew signal input
rlabel metal2 s 44546 99200 44602 100000 6 sram_dout1[76]
port 290 nsew signal input
rlabel metal2 s 45006 99200 45062 100000 6 sram_dout1[77]
port 291 nsew signal input
rlabel metal2 s 45558 99200 45614 100000 6 sram_dout1[78]
port 292 nsew signal input
rlabel metal2 s 46018 99200 46074 100000 6 sram_dout1[79]
port 293 nsew signal input
rlabel metal2 s 10506 99200 10562 100000 6 sram_dout1[7]
port 294 nsew signal input
rlabel metal2 s 46478 99200 46534 100000 6 sram_dout1[80]
port 295 nsew signal input
rlabel metal2 s 47030 99200 47086 100000 6 sram_dout1[81]
port 296 nsew signal input
rlabel metal2 s 47490 99200 47546 100000 6 sram_dout1[82]
port 297 nsew signal input
rlabel metal2 s 47950 99200 48006 100000 6 sram_dout1[83]
port 298 nsew signal input
rlabel metal2 s 48502 99200 48558 100000 6 sram_dout1[84]
port 299 nsew signal input
rlabel metal2 s 48962 99200 49018 100000 6 sram_dout1[85]
port 300 nsew signal input
rlabel metal2 s 49422 99200 49478 100000 6 sram_dout1[86]
port 301 nsew signal input
rlabel metal2 s 49974 99200 50030 100000 6 sram_dout1[87]
port 302 nsew signal input
rlabel metal2 s 50434 99200 50490 100000 6 sram_dout1[88]
port 303 nsew signal input
rlabel metal2 s 50894 99200 50950 100000 6 sram_dout1[89]
port 304 nsew signal input
rlabel metal2 s 10966 99200 11022 100000 6 sram_dout1[8]
port 305 nsew signal input
rlabel metal2 s 51446 99200 51502 100000 6 sram_dout1[90]
port 306 nsew signal input
rlabel metal2 s 51906 99200 51962 100000 6 sram_dout1[91]
port 307 nsew signal input
rlabel metal2 s 52458 99200 52514 100000 6 sram_dout1[92]
port 308 nsew signal input
rlabel metal2 s 52918 99200 52974 100000 6 sram_dout1[93]
port 309 nsew signal input
rlabel metal2 s 53378 99200 53434 100000 6 sram_dout1[94]
port 310 nsew signal input
rlabel metal2 s 53930 99200 53986 100000 6 sram_dout1[95]
port 311 nsew signal input
rlabel metal2 s 54390 99200 54446 100000 6 sram_dout1[96]
port 312 nsew signal input
rlabel metal2 s 54850 99200 54906 100000 6 sram_dout1[97]
port 313 nsew signal input
rlabel metal2 s 55402 99200 55458 100000 6 sram_dout1[98]
port 314 nsew signal input
rlabel metal2 s 55862 99200 55918 100000 6 sram_dout1[99]
port 315 nsew signal input
rlabel metal2 s 11518 99200 11574 100000 6 sram_dout1[9]
port 316 nsew signal input
rlabel metal3 s 69200 3000 70000 3120 6 sram_web0
port 317 nsew signal output
rlabel metal3 s 69200 3544 70000 3664 6 sram_wmask0[0]
port 318 nsew signal output
rlabel metal3 s 69200 4088 70000 4208 6 sram_wmask0[1]
port 319 nsew signal output
rlabel metal3 s 69200 4632 70000 4752 6 sram_wmask0[2]
port 320 nsew signal output
rlabel metal3 s 69200 5176 70000 5296 6 sram_wmask0[3]
port 321 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal2 s 66350 0 66406 800 6 vga_b[0]
port 323 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 vga_b[1]
port 324 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 vga_g[0]
port 325 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 vga_g[1]
port 326 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 vga_hsync
port 327 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 vga_r[0]
port 328 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 vga_r[1]
port 329 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 vga_vsync
port 330 nsew signal output
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 331 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 331 nsew ground bidirectional
rlabel metal2 s 294 0 350 800 6 wb_ack_o
port 332 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 wb_adr_i[0]
port 333 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wb_adr_i[10]
port 334 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wb_adr_i[11]
port 335 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wb_adr_i[12]
port 336 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wb_adr_i[13]
port 337 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wb_adr_i[14]
port 338 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wb_adr_i[15]
port 339 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wb_adr_i[16]
port 340 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wb_adr_i[17]
port 341 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wb_adr_i[18]
port 342 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wb_adr_i[19]
port 343 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wb_adr_i[1]
port 344 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wb_adr_i[20]
port 345 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wb_adr_i[21]
port 346 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wb_adr_i[22]
port 347 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wb_adr_i[23]
port 348 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_adr_i[2]
port 349 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wb_adr_i[3]
port 350 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wb_adr_i[4]
port 351 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wb_adr_i[5]
port 352 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wb_adr_i[6]
port 353 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wb_adr_i[7]
port 354 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wb_adr_i[8]
port 355 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wb_adr_i[9]
port 356 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_clk_i
port 357 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wb_cyc_i
port 358 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wb_data_i[0]
port 359 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wb_data_i[10]
port 360 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wb_data_i[11]
port 361 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wb_data_i[12]
port 362 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wb_data_i[13]
port 363 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wb_data_i[14]
port 364 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wb_data_i[15]
port 365 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wb_data_i[16]
port 366 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wb_data_i[17]
port 367 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wb_data_i[18]
port 368 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wb_data_i[19]
port 369 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wb_data_i[1]
port 370 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wb_data_i[20]
port 371 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wb_data_i[21]
port 372 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 wb_data_i[22]
port 373 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wb_data_i[23]
port 374 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 wb_data_i[24]
port 375 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 wb_data_i[25]
port 376 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wb_data_i[26]
port 377 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 wb_data_i[27]
port 378 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wb_data_i[28]
port 379 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wb_data_i[29]
port 380 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wb_data_i[2]
port 381 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 wb_data_i[30]
port 382 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 wb_data_i[31]
port 383 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wb_data_i[3]
port 384 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wb_data_i[4]
port 385 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wb_data_i[5]
port 386 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wb_data_i[6]
port 387 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wb_data_i[7]
port 388 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wb_data_i[8]
port 389 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wb_data_i[9]
port 390 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wb_data_o[0]
port 391 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wb_data_o[10]
port 392 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wb_data_o[11]
port 393 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 wb_data_o[12]
port 394 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wb_data_o[13]
port 395 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wb_data_o[14]
port 396 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wb_data_o[15]
port 397 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 wb_data_o[16]
port 398 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 wb_data_o[17]
port 399 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wb_data_o[18]
port 400 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wb_data_o[19]
port 401 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wb_data_o[1]
port 402 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wb_data_o[20]
port 403 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wb_data_o[21]
port 404 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wb_data_o[22]
port 405 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wb_data_o[23]
port 406 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wb_data_o[24]
port 407 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wb_data_o[25]
port 408 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 wb_data_o[26]
port 409 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 wb_data_o[27]
port 410 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 wb_data_o[28]
port 411 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 wb_data_o[29]
port 412 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wb_data_o[2]
port 413 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 wb_data_o[30]
port 414 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 wb_data_o[31]
port 415 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wb_data_o[3]
port 416 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wb_data_o[4]
port 417 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 wb_data_o[5]
port 418 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wb_data_o[6]
port 419 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wb_data_o[7]
port 420 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wb_data_o[8]
port 421 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 wb_data_o[9]
port 422 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wb_error_o
port 423 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 wb_rst_i
port 424 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wb_sel_i[0]
port 425 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wb_sel_i[1]
port 426 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wb_sel_i[2]
port 427 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wb_sel_i[3]
port 428 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wb_stall_o
port 429 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wb_stb_i
port 430 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wb_we_i
port 431 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6569284
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Video/runs/Video/results/signoff/Video.magic.gds
string GDS_START 696274
<< end >>

