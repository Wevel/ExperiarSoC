magic
tech sky130A
magscale 1 2
timestamp 1653219018
<< obsli1 >>
rect 1104 2159 78844 157777
<< obsm1 >>
rect 658 1300 79290 158432
<< metal2 >>
rect 1030 159200 1086 160000
rect 3054 159200 3110 160000
rect 5078 159200 5134 160000
rect 7102 159200 7158 160000
rect 9218 159200 9274 160000
rect 11242 159200 11298 160000
rect 13266 159200 13322 160000
rect 15382 159200 15438 160000
rect 17406 159200 17462 160000
rect 19430 159200 19486 160000
rect 21546 159200 21602 160000
rect 23570 159200 23626 160000
rect 25594 159200 25650 160000
rect 27710 159200 27766 160000
rect 29734 159200 29790 160000
rect 31758 159200 31814 160000
rect 33782 159200 33838 160000
rect 35898 159200 35954 160000
rect 37922 159200 37978 160000
rect 39946 159200 40002 160000
rect 42062 159200 42118 160000
rect 44086 159200 44142 160000
rect 46110 159200 46166 160000
rect 48226 159200 48282 160000
rect 50250 159200 50306 160000
rect 52274 159200 52330 160000
rect 54390 159200 54446 160000
rect 56414 159200 56470 160000
rect 58438 159200 58494 160000
rect 60462 159200 60518 160000
rect 62578 159200 62634 160000
rect 64602 159200 64658 160000
rect 66626 159200 66682 160000
rect 68742 159200 68798 160000
rect 70766 159200 70822 160000
rect 72790 159200 72846 160000
rect 74906 159200 74962 160000
rect 76930 159200 76986 160000
rect 78954 159200 79010 160000
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4986 0 5042 800
rect 6458 0 6514 800
rect 7930 0 7986 800
rect 9310 0 9366 800
rect 10782 0 10838 800
rect 12254 0 12310 800
rect 13726 0 13782 800
rect 15198 0 15254 800
rect 16670 0 16726 800
rect 18050 0 18106 800
rect 19522 0 19578 800
rect 20994 0 21050 800
rect 22466 0 22522 800
rect 23938 0 23994 800
rect 25318 0 25374 800
rect 26790 0 26846 800
rect 28262 0 28318 800
rect 29734 0 29790 800
rect 31206 0 31262 800
rect 32678 0 32734 800
rect 34058 0 34114 800
rect 35530 0 35586 800
rect 37002 0 37058 800
rect 38474 0 38530 800
rect 39946 0 40002 800
rect 41326 0 41382 800
rect 42798 0 42854 800
rect 44270 0 44326 800
rect 45742 0 45798 800
rect 47214 0 47270 800
rect 48686 0 48742 800
rect 50066 0 50122 800
rect 51538 0 51594 800
rect 53010 0 53066 800
rect 54482 0 54538 800
rect 55954 0 56010 800
rect 57334 0 57390 800
rect 58806 0 58862 800
rect 60278 0 60334 800
rect 61750 0 61806 800
rect 63222 0 63278 800
rect 64694 0 64750 800
rect 66074 0 66130 800
rect 67546 0 67602 800
rect 69018 0 69074 800
rect 70490 0 70546 800
rect 71962 0 72018 800
rect 73342 0 73398 800
rect 74814 0 74870 800
rect 76286 0 76342 800
rect 77758 0 77814 800
rect 79230 0 79286 800
<< obsm2 >>
rect 664 159144 974 159497
rect 1142 159144 2998 159497
rect 3166 159144 5022 159497
rect 5190 159144 7046 159497
rect 7214 159144 9162 159497
rect 9330 159144 11186 159497
rect 11354 159144 13210 159497
rect 13378 159144 15326 159497
rect 15494 159144 17350 159497
rect 17518 159144 19374 159497
rect 19542 159144 21490 159497
rect 21658 159144 23514 159497
rect 23682 159144 25538 159497
rect 25706 159144 27654 159497
rect 27822 159144 29678 159497
rect 29846 159144 31702 159497
rect 31870 159144 33726 159497
rect 33894 159144 35842 159497
rect 36010 159144 37866 159497
rect 38034 159144 39890 159497
rect 40058 159144 42006 159497
rect 42174 159144 44030 159497
rect 44198 159144 46054 159497
rect 46222 159144 48170 159497
rect 48338 159144 50194 159497
rect 50362 159144 52218 159497
rect 52386 159144 54334 159497
rect 54502 159144 56358 159497
rect 56526 159144 58382 159497
rect 58550 159144 60406 159497
rect 60574 159144 62522 159497
rect 62690 159144 64546 159497
rect 64714 159144 66570 159497
rect 66738 159144 68686 159497
rect 68854 159144 70710 159497
rect 70878 159144 72734 159497
rect 72902 159144 74850 159497
rect 75018 159144 76874 159497
rect 77042 159144 78898 159497
rect 79066 159144 79284 159497
rect 664 856 79284 159144
rect 774 303 1986 856
rect 2154 303 3458 856
rect 3626 303 4930 856
rect 5098 303 6402 856
rect 6570 303 7874 856
rect 8042 303 9254 856
rect 9422 303 10726 856
rect 10894 303 12198 856
rect 12366 303 13670 856
rect 13838 303 15142 856
rect 15310 303 16614 856
rect 16782 303 17994 856
rect 18162 303 19466 856
rect 19634 303 20938 856
rect 21106 303 22410 856
rect 22578 303 23882 856
rect 24050 303 25262 856
rect 25430 303 26734 856
rect 26902 303 28206 856
rect 28374 303 29678 856
rect 29846 303 31150 856
rect 31318 303 32622 856
rect 32790 303 34002 856
rect 34170 303 35474 856
rect 35642 303 36946 856
rect 37114 303 38418 856
rect 38586 303 39890 856
rect 40058 303 41270 856
rect 41438 303 42742 856
rect 42910 303 44214 856
rect 44382 303 45686 856
rect 45854 303 47158 856
rect 47326 303 48630 856
rect 48798 303 50010 856
rect 50178 303 51482 856
rect 51650 303 52954 856
rect 53122 303 54426 856
rect 54594 303 55898 856
rect 56066 303 57278 856
rect 57446 303 58750 856
rect 58918 303 60222 856
rect 60390 303 61694 856
rect 61862 303 63166 856
rect 63334 303 64638 856
rect 64806 303 66018 856
rect 66186 303 67490 856
rect 67658 303 68962 856
rect 69130 303 70434 856
rect 70602 303 71906 856
rect 72074 303 73286 856
rect 73454 303 74758 856
rect 74926 303 76230 856
rect 76398 303 77702 856
rect 77870 303 79174 856
<< metal3 >>
rect 0 159400 800 159520
rect 79200 159400 80000 159520
rect 0 158584 800 158704
rect 79200 158584 80000 158704
rect 0 157768 800 157888
rect 79200 157768 80000 157888
rect 0 156952 800 157072
rect 79200 156952 80000 157072
rect 0 156136 800 156256
rect 79200 156136 80000 156256
rect 0 155320 800 155440
rect 79200 155456 80000 155576
rect 0 154504 800 154624
rect 79200 154640 80000 154760
rect 0 153688 800 153808
rect 79200 153824 80000 153944
rect 0 152872 800 152992
rect 79200 153008 80000 153128
rect 0 152056 800 152176
rect 79200 152192 80000 152312
rect 79200 151376 80000 151496
rect 0 151104 800 151224
rect 79200 150696 80000 150816
rect 0 150288 800 150408
rect 79200 149880 80000 150000
rect 0 149472 800 149592
rect 79200 149064 80000 149184
rect 0 148656 800 148776
rect 79200 148248 80000 148368
rect 0 147840 800 147960
rect 79200 147432 80000 147552
rect 0 147024 800 147144
rect 79200 146752 80000 146872
rect 0 146208 800 146328
rect 79200 145936 80000 146056
rect 0 145392 800 145512
rect 79200 145120 80000 145240
rect 0 144576 800 144696
rect 79200 144304 80000 144424
rect 0 143760 800 143880
rect 79200 143488 80000 143608
rect 0 142944 800 143064
rect 79200 142672 80000 142792
rect 0 141992 800 142112
rect 79200 141992 80000 142112
rect 0 141176 800 141296
rect 79200 141176 80000 141296
rect 0 140360 800 140480
rect 79200 140360 80000 140480
rect 0 139544 800 139664
rect 79200 139544 80000 139664
rect 0 138728 800 138848
rect 79200 138728 80000 138848
rect 0 137912 800 138032
rect 79200 137912 80000 138032
rect 0 137096 800 137216
rect 79200 137232 80000 137352
rect 0 136280 800 136400
rect 79200 136416 80000 136536
rect 0 135464 800 135584
rect 79200 135600 80000 135720
rect 0 134648 800 134768
rect 79200 134784 80000 134904
rect 0 133832 800 133952
rect 79200 133968 80000 134088
rect 79200 133288 80000 133408
rect 0 132880 800 133000
rect 79200 132472 80000 132592
rect 0 132064 800 132184
rect 79200 131656 80000 131776
rect 0 131248 800 131368
rect 79200 130840 80000 130960
rect 0 130432 800 130552
rect 79200 130024 80000 130144
rect 0 129616 800 129736
rect 79200 129208 80000 129328
rect 0 128800 800 128920
rect 79200 128528 80000 128648
rect 0 127984 800 128104
rect 79200 127712 80000 127832
rect 0 127168 800 127288
rect 79200 126896 80000 127016
rect 0 126352 800 126472
rect 79200 126080 80000 126200
rect 0 125536 800 125656
rect 79200 125264 80000 125384
rect 0 124584 800 124704
rect 79200 124584 80000 124704
rect 0 123768 800 123888
rect 79200 123768 80000 123888
rect 0 122952 800 123072
rect 79200 122952 80000 123072
rect 0 122136 800 122256
rect 79200 122136 80000 122256
rect 0 121320 800 121440
rect 79200 121320 80000 121440
rect 0 120504 800 120624
rect 79200 120504 80000 120624
rect 0 119688 800 119808
rect 79200 119824 80000 119944
rect 0 118872 800 118992
rect 79200 119008 80000 119128
rect 0 118056 800 118176
rect 79200 118192 80000 118312
rect 0 117240 800 117360
rect 79200 117376 80000 117496
rect 0 116424 800 116544
rect 79200 116560 80000 116680
rect 79200 115744 80000 115864
rect 0 115472 800 115592
rect 79200 115064 80000 115184
rect 0 114656 800 114776
rect 79200 114248 80000 114368
rect 0 113840 800 113960
rect 79200 113432 80000 113552
rect 0 113024 800 113144
rect 79200 112616 80000 112736
rect 0 112208 800 112328
rect 79200 111800 80000 111920
rect 0 111392 800 111512
rect 79200 111120 80000 111240
rect 0 110576 800 110696
rect 79200 110304 80000 110424
rect 0 109760 800 109880
rect 79200 109488 80000 109608
rect 0 108944 800 109064
rect 79200 108672 80000 108792
rect 0 108128 800 108248
rect 79200 107856 80000 107976
rect 0 107312 800 107432
rect 79200 107040 80000 107160
rect 0 106360 800 106480
rect 79200 106360 80000 106480
rect 0 105544 800 105664
rect 79200 105544 80000 105664
rect 0 104728 800 104848
rect 79200 104728 80000 104848
rect 0 103912 800 104032
rect 79200 103912 80000 104032
rect 0 103096 800 103216
rect 79200 103096 80000 103216
rect 0 102280 800 102400
rect 79200 102416 80000 102536
rect 0 101464 800 101584
rect 79200 101600 80000 101720
rect 0 100648 800 100768
rect 79200 100784 80000 100904
rect 0 99832 800 99952
rect 79200 99968 80000 100088
rect 0 99016 800 99136
rect 79200 99152 80000 99272
rect 0 98200 800 98320
rect 79200 98336 80000 98456
rect 79200 97656 80000 97776
rect 0 97248 800 97368
rect 79200 96840 80000 96960
rect 0 96432 800 96552
rect 79200 96024 80000 96144
rect 0 95616 800 95736
rect 79200 95208 80000 95328
rect 0 94800 800 94920
rect 79200 94392 80000 94512
rect 0 93984 800 94104
rect 79200 93576 80000 93696
rect 0 93168 800 93288
rect 79200 92896 80000 93016
rect 0 92352 800 92472
rect 79200 92080 80000 92200
rect 0 91536 800 91656
rect 79200 91264 80000 91384
rect 0 90720 800 90840
rect 79200 90448 80000 90568
rect 0 89904 800 90024
rect 79200 89632 80000 89752
rect 0 88952 800 89072
rect 79200 88952 80000 89072
rect 0 88136 800 88256
rect 79200 88136 80000 88256
rect 0 87320 800 87440
rect 79200 87320 80000 87440
rect 0 86504 800 86624
rect 79200 86504 80000 86624
rect 0 85688 800 85808
rect 79200 85688 80000 85808
rect 0 84872 800 84992
rect 79200 84872 80000 84992
rect 0 84056 800 84176
rect 79200 84192 80000 84312
rect 0 83240 800 83360
rect 79200 83376 80000 83496
rect 0 82424 800 82544
rect 79200 82560 80000 82680
rect 0 81608 800 81728
rect 79200 81744 80000 81864
rect 0 80792 800 80912
rect 79200 80928 80000 81048
rect 79200 80248 80000 80368
rect 0 79840 800 79960
rect 79200 79432 80000 79552
rect 0 79024 800 79144
rect 79200 78616 80000 78736
rect 0 78208 800 78328
rect 79200 77800 80000 77920
rect 0 77392 800 77512
rect 79200 76984 80000 77104
rect 0 76576 800 76696
rect 79200 76168 80000 76288
rect 0 75760 800 75880
rect 79200 75488 80000 75608
rect 0 74944 800 75064
rect 79200 74672 80000 74792
rect 0 74128 800 74248
rect 79200 73856 80000 73976
rect 0 73312 800 73432
rect 79200 73040 80000 73160
rect 0 72496 800 72616
rect 79200 72224 80000 72344
rect 0 71680 800 71800
rect 79200 71408 80000 71528
rect 0 70728 800 70848
rect 79200 70728 80000 70848
rect 0 69912 800 70032
rect 79200 69912 80000 70032
rect 0 69096 800 69216
rect 79200 69096 80000 69216
rect 0 68280 800 68400
rect 79200 68280 80000 68400
rect 0 67464 800 67584
rect 79200 67464 80000 67584
rect 0 66648 800 66768
rect 79200 66784 80000 66904
rect 0 65832 800 65952
rect 79200 65968 80000 66088
rect 0 65016 800 65136
rect 79200 65152 80000 65272
rect 0 64200 800 64320
rect 79200 64336 80000 64456
rect 0 63384 800 63504
rect 79200 63520 80000 63640
rect 79200 62704 80000 62824
rect 0 62432 800 62552
rect 79200 62024 80000 62144
rect 0 61616 800 61736
rect 79200 61208 80000 61328
rect 0 60800 800 60920
rect 79200 60392 80000 60512
rect 0 59984 800 60104
rect 79200 59576 80000 59696
rect 0 59168 800 59288
rect 79200 58760 80000 58880
rect 0 58352 800 58472
rect 79200 57944 80000 58064
rect 0 57536 800 57656
rect 79200 57264 80000 57384
rect 0 56720 800 56840
rect 79200 56448 80000 56568
rect 0 55904 800 56024
rect 79200 55632 80000 55752
rect 0 55088 800 55208
rect 79200 54816 80000 54936
rect 0 54272 800 54392
rect 79200 54000 80000 54120
rect 0 53320 800 53440
rect 79200 53320 80000 53440
rect 0 52504 800 52624
rect 79200 52504 80000 52624
rect 0 51688 800 51808
rect 79200 51688 80000 51808
rect 0 50872 800 50992
rect 79200 50872 80000 50992
rect 0 50056 800 50176
rect 79200 50056 80000 50176
rect 0 49240 800 49360
rect 79200 49240 80000 49360
rect 0 48424 800 48544
rect 79200 48560 80000 48680
rect 0 47608 800 47728
rect 79200 47744 80000 47864
rect 0 46792 800 46912
rect 79200 46928 80000 47048
rect 0 45976 800 46096
rect 79200 46112 80000 46232
rect 0 45160 800 45280
rect 79200 45296 80000 45416
rect 79200 44616 80000 44736
rect 0 44208 800 44328
rect 79200 43800 80000 43920
rect 0 43392 800 43512
rect 79200 42984 80000 43104
rect 0 42576 800 42696
rect 79200 42168 80000 42288
rect 0 41760 800 41880
rect 79200 41352 80000 41472
rect 0 40944 800 41064
rect 79200 40536 80000 40656
rect 0 40128 800 40248
rect 79200 39856 80000 39976
rect 0 39312 800 39432
rect 79200 39040 80000 39160
rect 0 38496 800 38616
rect 79200 38224 80000 38344
rect 0 37680 800 37800
rect 79200 37408 80000 37528
rect 0 36864 800 36984
rect 79200 36592 80000 36712
rect 0 36048 800 36168
rect 79200 35776 80000 35896
rect 0 35096 800 35216
rect 79200 35096 80000 35216
rect 0 34280 800 34400
rect 79200 34280 80000 34400
rect 0 33464 800 33584
rect 79200 33464 80000 33584
rect 0 32648 800 32768
rect 79200 32648 80000 32768
rect 0 31832 800 31952
rect 79200 31832 80000 31952
rect 0 31016 800 31136
rect 79200 31152 80000 31272
rect 0 30200 800 30320
rect 79200 30336 80000 30456
rect 0 29384 800 29504
rect 79200 29520 80000 29640
rect 0 28568 800 28688
rect 79200 28704 80000 28824
rect 0 27752 800 27872
rect 79200 27888 80000 28008
rect 79200 27072 80000 27192
rect 0 26800 800 26920
rect 79200 26392 80000 26512
rect 0 25984 800 26104
rect 79200 25576 80000 25696
rect 0 25168 800 25288
rect 79200 24760 80000 24880
rect 0 24352 800 24472
rect 79200 23944 80000 24064
rect 0 23536 800 23656
rect 79200 23128 80000 23248
rect 0 22720 800 22840
rect 79200 22448 80000 22568
rect 0 21904 800 22024
rect 79200 21632 80000 21752
rect 0 21088 800 21208
rect 79200 20816 80000 20936
rect 0 20272 800 20392
rect 79200 20000 80000 20120
rect 0 19456 800 19576
rect 79200 19184 80000 19304
rect 0 18640 800 18760
rect 79200 18368 80000 18488
rect 0 17688 800 17808
rect 79200 17688 80000 17808
rect 0 16872 800 16992
rect 79200 16872 80000 16992
rect 0 16056 800 16176
rect 79200 16056 80000 16176
rect 0 15240 800 15360
rect 79200 15240 80000 15360
rect 0 14424 800 14544
rect 79200 14424 80000 14544
rect 0 13608 800 13728
rect 79200 13608 80000 13728
rect 0 12792 800 12912
rect 79200 12928 80000 13048
rect 0 11976 800 12096
rect 79200 12112 80000 12232
rect 0 11160 800 11280
rect 79200 11296 80000 11416
rect 0 10344 800 10464
rect 79200 10480 80000 10600
rect 0 9528 800 9648
rect 79200 9664 80000 9784
rect 79200 8984 80000 9104
rect 0 8576 800 8696
rect 79200 8168 80000 8288
rect 0 7760 800 7880
rect 79200 7352 80000 7472
rect 0 6944 800 7064
rect 79200 6536 80000 6656
rect 0 6128 800 6248
rect 79200 5720 80000 5840
rect 0 5312 800 5432
rect 79200 4904 80000 5024
rect 0 4496 800 4616
rect 79200 4224 80000 4344
rect 0 3680 800 3800
rect 79200 3408 80000 3528
rect 0 2864 800 2984
rect 79200 2592 80000 2712
rect 0 2048 800 2168
rect 79200 1776 80000 1896
rect 0 1232 800 1352
rect 79200 960 80000 1080
rect 0 416 800 536
rect 79200 280 80000 400
<< obsm3 >>
rect 880 159320 79120 159493
rect 800 158784 79200 159320
rect 880 158504 79120 158784
rect 800 157968 79200 158504
rect 880 157688 79120 157968
rect 800 157152 79200 157688
rect 880 156872 79120 157152
rect 800 156336 79200 156872
rect 880 156056 79120 156336
rect 800 155656 79200 156056
rect 800 155520 79120 155656
rect 880 155376 79120 155520
rect 880 155240 79200 155376
rect 800 154840 79200 155240
rect 800 154704 79120 154840
rect 880 154560 79120 154704
rect 880 154424 79200 154560
rect 800 154024 79200 154424
rect 800 153888 79120 154024
rect 880 153744 79120 153888
rect 880 153608 79200 153744
rect 800 153208 79200 153608
rect 800 153072 79120 153208
rect 880 152928 79120 153072
rect 880 152792 79200 152928
rect 800 152392 79200 152792
rect 800 152256 79120 152392
rect 880 152112 79120 152256
rect 880 151976 79200 152112
rect 800 151576 79200 151976
rect 800 151304 79120 151576
rect 880 151296 79120 151304
rect 880 151024 79200 151296
rect 800 150896 79200 151024
rect 800 150616 79120 150896
rect 800 150488 79200 150616
rect 880 150208 79200 150488
rect 800 150080 79200 150208
rect 800 149800 79120 150080
rect 800 149672 79200 149800
rect 880 149392 79200 149672
rect 800 149264 79200 149392
rect 800 148984 79120 149264
rect 800 148856 79200 148984
rect 880 148576 79200 148856
rect 800 148448 79200 148576
rect 800 148168 79120 148448
rect 800 148040 79200 148168
rect 880 147760 79200 148040
rect 800 147632 79200 147760
rect 800 147352 79120 147632
rect 800 147224 79200 147352
rect 880 146952 79200 147224
rect 880 146944 79120 146952
rect 800 146672 79120 146944
rect 800 146408 79200 146672
rect 880 146136 79200 146408
rect 880 146128 79120 146136
rect 800 145856 79120 146128
rect 800 145592 79200 145856
rect 880 145320 79200 145592
rect 880 145312 79120 145320
rect 800 145040 79120 145312
rect 800 144776 79200 145040
rect 880 144504 79200 144776
rect 880 144496 79120 144504
rect 800 144224 79120 144496
rect 800 143960 79200 144224
rect 880 143688 79200 143960
rect 880 143680 79120 143688
rect 800 143408 79120 143680
rect 800 143144 79200 143408
rect 880 142872 79200 143144
rect 880 142864 79120 142872
rect 800 142592 79120 142864
rect 800 142192 79200 142592
rect 880 141912 79120 142192
rect 800 141376 79200 141912
rect 880 141096 79120 141376
rect 800 140560 79200 141096
rect 880 140280 79120 140560
rect 800 139744 79200 140280
rect 880 139464 79120 139744
rect 800 138928 79200 139464
rect 880 138648 79120 138928
rect 800 138112 79200 138648
rect 880 137832 79120 138112
rect 800 137432 79200 137832
rect 800 137296 79120 137432
rect 880 137152 79120 137296
rect 880 137016 79200 137152
rect 800 136616 79200 137016
rect 800 136480 79120 136616
rect 880 136336 79120 136480
rect 880 136200 79200 136336
rect 800 135800 79200 136200
rect 800 135664 79120 135800
rect 880 135520 79120 135664
rect 880 135384 79200 135520
rect 800 134984 79200 135384
rect 800 134848 79120 134984
rect 880 134704 79120 134848
rect 880 134568 79200 134704
rect 800 134168 79200 134568
rect 800 134032 79120 134168
rect 880 133888 79120 134032
rect 880 133752 79200 133888
rect 800 133488 79200 133752
rect 800 133208 79120 133488
rect 800 133080 79200 133208
rect 880 132800 79200 133080
rect 800 132672 79200 132800
rect 800 132392 79120 132672
rect 800 132264 79200 132392
rect 880 131984 79200 132264
rect 800 131856 79200 131984
rect 800 131576 79120 131856
rect 800 131448 79200 131576
rect 880 131168 79200 131448
rect 800 131040 79200 131168
rect 800 130760 79120 131040
rect 800 130632 79200 130760
rect 880 130352 79200 130632
rect 800 130224 79200 130352
rect 800 129944 79120 130224
rect 800 129816 79200 129944
rect 880 129536 79200 129816
rect 800 129408 79200 129536
rect 800 129128 79120 129408
rect 800 129000 79200 129128
rect 880 128728 79200 129000
rect 880 128720 79120 128728
rect 800 128448 79120 128720
rect 800 128184 79200 128448
rect 880 127912 79200 128184
rect 880 127904 79120 127912
rect 800 127632 79120 127904
rect 800 127368 79200 127632
rect 880 127096 79200 127368
rect 880 127088 79120 127096
rect 800 126816 79120 127088
rect 800 126552 79200 126816
rect 880 126280 79200 126552
rect 880 126272 79120 126280
rect 800 126000 79120 126272
rect 800 125736 79200 126000
rect 880 125464 79200 125736
rect 880 125456 79120 125464
rect 800 125184 79120 125456
rect 800 124784 79200 125184
rect 880 124504 79120 124784
rect 800 123968 79200 124504
rect 880 123688 79120 123968
rect 800 123152 79200 123688
rect 880 122872 79120 123152
rect 800 122336 79200 122872
rect 880 122056 79120 122336
rect 800 121520 79200 122056
rect 880 121240 79120 121520
rect 800 120704 79200 121240
rect 880 120424 79120 120704
rect 800 120024 79200 120424
rect 800 119888 79120 120024
rect 880 119744 79120 119888
rect 880 119608 79200 119744
rect 800 119208 79200 119608
rect 800 119072 79120 119208
rect 880 118928 79120 119072
rect 880 118792 79200 118928
rect 800 118392 79200 118792
rect 800 118256 79120 118392
rect 880 118112 79120 118256
rect 880 117976 79200 118112
rect 800 117576 79200 117976
rect 800 117440 79120 117576
rect 880 117296 79120 117440
rect 880 117160 79200 117296
rect 800 116760 79200 117160
rect 800 116624 79120 116760
rect 880 116480 79120 116624
rect 880 116344 79200 116480
rect 800 115944 79200 116344
rect 800 115672 79120 115944
rect 880 115664 79120 115672
rect 880 115392 79200 115664
rect 800 115264 79200 115392
rect 800 114984 79120 115264
rect 800 114856 79200 114984
rect 880 114576 79200 114856
rect 800 114448 79200 114576
rect 800 114168 79120 114448
rect 800 114040 79200 114168
rect 880 113760 79200 114040
rect 800 113632 79200 113760
rect 800 113352 79120 113632
rect 800 113224 79200 113352
rect 880 112944 79200 113224
rect 800 112816 79200 112944
rect 800 112536 79120 112816
rect 800 112408 79200 112536
rect 880 112128 79200 112408
rect 800 112000 79200 112128
rect 800 111720 79120 112000
rect 800 111592 79200 111720
rect 880 111320 79200 111592
rect 880 111312 79120 111320
rect 800 111040 79120 111312
rect 800 110776 79200 111040
rect 880 110504 79200 110776
rect 880 110496 79120 110504
rect 800 110224 79120 110496
rect 800 109960 79200 110224
rect 880 109688 79200 109960
rect 880 109680 79120 109688
rect 800 109408 79120 109680
rect 800 109144 79200 109408
rect 880 108872 79200 109144
rect 880 108864 79120 108872
rect 800 108592 79120 108864
rect 800 108328 79200 108592
rect 880 108056 79200 108328
rect 880 108048 79120 108056
rect 800 107776 79120 108048
rect 800 107512 79200 107776
rect 880 107240 79200 107512
rect 880 107232 79120 107240
rect 800 106960 79120 107232
rect 800 106560 79200 106960
rect 880 106280 79120 106560
rect 800 105744 79200 106280
rect 880 105464 79120 105744
rect 800 104928 79200 105464
rect 880 104648 79120 104928
rect 800 104112 79200 104648
rect 880 103832 79120 104112
rect 800 103296 79200 103832
rect 880 103016 79120 103296
rect 800 102616 79200 103016
rect 800 102480 79120 102616
rect 880 102336 79120 102480
rect 880 102200 79200 102336
rect 800 101800 79200 102200
rect 800 101664 79120 101800
rect 880 101520 79120 101664
rect 880 101384 79200 101520
rect 800 100984 79200 101384
rect 800 100848 79120 100984
rect 880 100704 79120 100848
rect 880 100568 79200 100704
rect 800 100168 79200 100568
rect 800 100032 79120 100168
rect 880 99888 79120 100032
rect 880 99752 79200 99888
rect 800 99352 79200 99752
rect 800 99216 79120 99352
rect 880 99072 79120 99216
rect 880 98936 79200 99072
rect 800 98536 79200 98936
rect 800 98400 79120 98536
rect 880 98256 79120 98400
rect 880 98120 79200 98256
rect 800 97856 79200 98120
rect 800 97576 79120 97856
rect 800 97448 79200 97576
rect 880 97168 79200 97448
rect 800 97040 79200 97168
rect 800 96760 79120 97040
rect 800 96632 79200 96760
rect 880 96352 79200 96632
rect 800 96224 79200 96352
rect 800 95944 79120 96224
rect 800 95816 79200 95944
rect 880 95536 79200 95816
rect 800 95408 79200 95536
rect 800 95128 79120 95408
rect 800 95000 79200 95128
rect 880 94720 79200 95000
rect 800 94592 79200 94720
rect 800 94312 79120 94592
rect 800 94184 79200 94312
rect 880 93904 79200 94184
rect 800 93776 79200 93904
rect 800 93496 79120 93776
rect 800 93368 79200 93496
rect 880 93096 79200 93368
rect 880 93088 79120 93096
rect 800 92816 79120 93088
rect 800 92552 79200 92816
rect 880 92280 79200 92552
rect 880 92272 79120 92280
rect 800 92000 79120 92272
rect 800 91736 79200 92000
rect 880 91464 79200 91736
rect 880 91456 79120 91464
rect 800 91184 79120 91456
rect 800 90920 79200 91184
rect 880 90648 79200 90920
rect 880 90640 79120 90648
rect 800 90368 79120 90640
rect 800 90104 79200 90368
rect 880 89832 79200 90104
rect 880 89824 79120 89832
rect 800 89552 79120 89824
rect 800 89152 79200 89552
rect 880 88872 79120 89152
rect 800 88336 79200 88872
rect 880 88056 79120 88336
rect 800 87520 79200 88056
rect 880 87240 79120 87520
rect 800 86704 79200 87240
rect 880 86424 79120 86704
rect 800 85888 79200 86424
rect 880 85608 79120 85888
rect 800 85072 79200 85608
rect 880 84792 79120 85072
rect 800 84392 79200 84792
rect 800 84256 79120 84392
rect 880 84112 79120 84256
rect 880 83976 79200 84112
rect 800 83576 79200 83976
rect 800 83440 79120 83576
rect 880 83296 79120 83440
rect 880 83160 79200 83296
rect 800 82760 79200 83160
rect 800 82624 79120 82760
rect 880 82480 79120 82624
rect 880 82344 79200 82480
rect 800 81944 79200 82344
rect 800 81808 79120 81944
rect 880 81664 79120 81808
rect 880 81528 79200 81664
rect 800 81128 79200 81528
rect 800 80992 79120 81128
rect 880 80848 79120 80992
rect 880 80712 79200 80848
rect 800 80448 79200 80712
rect 800 80168 79120 80448
rect 800 80040 79200 80168
rect 880 79760 79200 80040
rect 800 79632 79200 79760
rect 800 79352 79120 79632
rect 800 79224 79200 79352
rect 880 78944 79200 79224
rect 800 78816 79200 78944
rect 800 78536 79120 78816
rect 800 78408 79200 78536
rect 880 78128 79200 78408
rect 800 78000 79200 78128
rect 800 77720 79120 78000
rect 800 77592 79200 77720
rect 880 77312 79200 77592
rect 800 77184 79200 77312
rect 800 76904 79120 77184
rect 800 76776 79200 76904
rect 880 76496 79200 76776
rect 800 76368 79200 76496
rect 800 76088 79120 76368
rect 800 75960 79200 76088
rect 880 75688 79200 75960
rect 880 75680 79120 75688
rect 800 75408 79120 75680
rect 800 75144 79200 75408
rect 880 74872 79200 75144
rect 880 74864 79120 74872
rect 800 74592 79120 74864
rect 800 74328 79200 74592
rect 880 74056 79200 74328
rect 880 74048 79120 74056
rect 800 73776 79120 74048
rect 800 73512 79200 73776
rect 880 73240 79200 73512
rect 880 73232 79120 73240
rect 800 72960 79120 73232
rect 800 72696 79200 72960
rect 880 72424 79200 72696
rect 880 72416 79120 72424
rect 800 72144 79120 72416
rect 800 71880 79200 72144
rect 880 71608 79200 71880
rect 880 71600 79120 71608
rect 800 71328 79120 71600
rect 800 70928 79200 71328
rect 880 70648 79120 70928
rect 800 70112 79200 70648
rect 880 69832 79120 70112
rect 800 69296 79200 69832
rect 880 69016 79120 69296
rect 800 68480 79200 69016
rect 880 68200 79120 68480
rect 800 67664 79200 68200
rect 880 67384 79120 67664
rect 800 66984 79200 67384
rect 800 66848 79120 66984
rect 880 66704 79120 66848
rect 880 66568 79200 66704
rect 800 66168 79200 66568
rect 800 66032 79120 66168
rect 880 65888 79120 66032
rect 880 65752 79200 65888
rect 800 65352 79200 65752
rect 800 65216 79120 65352
rect 880 65072 79120 65216
rect 880 64936 79200 65072
rect 800 64536 79200 64936
rect 800 64400 79120 64536
rect 880 64256 79120 64400
rect 880 64120 79200 64256
rect 800 63720 79200 64120
rect 800 63584 79120 63720
rect 880 63440 79120 63584
rect 880 63304 79200 63440
rect 800 62904 79200 63304
rect 800 62632 79120 62904
rect 880 62624 79120 62632
rect 880 62352 79200 62624
rect 800 62224 79200 62352
rect 800 61944 79120 62224
rect 800 61816 79200 61944
rect 880 61536 79200 61816
rect 800 61408 79200 61536
rect 800 61128 79120 61408
rect 800 61000 79200 61128
rect 880 60720 79200 61000
rect 800 60592 79200 60720
rect 800 60312 79120 60592
rect 800 60184 79200 60312
rect 880 59904 79200 60184
rect 800 59776 79200 59904
rect 800 59496 79120 59776
rect 800 59368 79200 59496
rect 880 59088 79200 59368
rect 800 58960 79200 59088
rect 800 58680 79120 58960
rect 800 58552 79200 58680
rect 880 58272 79200 58552
rect 800 58144 79200 58272
rect 800 57864 79120 58144
rect 800 57736 79200 57864
rect 880 57464 79200 57736
rect 880 57456 79120 57464
rect 800 57184 79120 57456
rect 800 56920 79200 57184
rect 880 56648 79200 56920
rect 880 56640 79120 56648
rect 800 56368 79120 56640
rect 800 56104 79200 56368
rect 880 55832 79200 56104
rect 880 55824 79120 55832
rect 800 55552 79120 55824
rect 800 55288 79200 55552
rect 880 55016 79200 55288
rect 880 55008 79120 55016
rect 800 54736 79120 55008
rect 800 54472 79200 54736
rect 880 54200 79200 54472
rect 880 54192 79120 54200
rect 800 53920 79120 54192
rect 800 53520 79200 53920
rect 880 53240 79120 53520
rect 800 52704 79200 53240
rect 880 52424 79120 52704
rect 800 51888 79200 52424
rect 880 51608 79120 51888
rect 800 51072 79200 51608
rect 880 50792 79120 51072
rect 800 50256 79200 50792
rect 880 49976 79120 50256
rect 800 49440 79200 49976
rect 880 49160 79120 49440
rect 800 48760 79200 49160
rect 800 48624 79120 48760
rect 880 48480 79120 48624
rect 880 48344 79200 48480
rect 800 47944 79200 48344
rect 800 47808 79120 47944
rect 880 47664 79120 47808
rect 880 47528 79200 47664
rect 800 47128 79200 47528
rect 800 46992 79120 47128
rect 880 46848 79120 46992
rect 880 46712 79200 46848
rect 800 46312 79200 46712
rect 800 46176 79120 46312
rect 880 46032 79120 46176
rect 880 45896 79200 46032
rect 800 45496 79200 45896
rect 800 45360 79120 45496
rect 880 45216 79120 45360
rect 880 45080 79200 45216
rect 800 44816 79200 45080
rect 800 44536 79120 44816
rect 800 44408 79200 44536
rect 880 44128 79200 44408
rect 800 44000 79200 44128
rect 800 43720 79120 44000
rect 800 43592 79200 43720
rect 880 43312 79200 43592
rect 800 43184 79200 43312
rect 800 42904 79120 43184
rect 800 42776 79200 42904
rect 880 42496 79200 42776
rect 800 42368 79200 42496
rect 800 42088 79120 42368
rect 800 41960 79200 42088
rect 880 41680 79200 41960
rect 800 41552 79200 41680
rect 800 41272 79120 41552
rect 800 41144 79200 41272
rect 880 40864 79200 41144
rect 800 40736 79200 40864
rect 800 40456 79120 40736
rect 800 40328 79200 40456
rect 880 40056 79200 40328
rect 880 40048 79120 40056
rect 800 39776 79120 40048
rect 800 39512 79200 39776
rect 880 39240 79200 39512
rect 880 39232 79120 39240
rect 800 38960 79120 39232
rect 800 38696 79200 38960
rect 880 38424 79200 38696
rect 880 38416 79120 38424
rect 800 38144 79120 38416
rect 800 37880 79200 38144
rect 880 37608 79200 37880
rect 880 37600 79120 37608
rect 800 37328 79120 37600
rect 800 37064 79200 37328
rect 880 36792 79200 37064
rect 880 36784 79120 36792
rect 800 36512 79120 36784
rect 800 36248 79200 36512
rect 880 35976 79200 36248
rect 880 35968 79120 35976
rect 800 35696 79120 35968
rect 800 35296 79200 35696
rect 880 35016 79120 35296
rect 800 34480 79200 35016
rect 880 34200 79120 34480
rect 800 33664 79200 34200
rect 880 33384 79120 33664
rect 800 32848 79200 33384
rect 880 32568 79120 32848
rect 800 32032 79200 32568
rect 880 31752 79120 32032
rect 800 31352 79200 31752
rect 800 31216 79120 31352
rect 880 31072 79120 31216
rect 880 30936 79200 31072
rect 800 30536 79200 30936
rect 800 30400 79120 30536
rect 880 30256 79120 30400
rect 880 30120 79200 30256
rect 800 29720 79200 30120
rect 800 29584 79120 29720
rect 880 29440 79120 29584
rect 880 29304 79200 29440
rect 800 28904 79200 29304
rect 800 28768 79120 28904
rect 880 28624 79120 28768
rect 880 28488 79200 28624
rect 800 28088 79200 28488
rect 800 27952 79120 28088
rect 880 27808 79120 27952
rect 880 27672 79200 27808
rect 800 27272 79200 27672
rect 800 27000 79120 27272
rect 880 26992 79120 27000
rect 880 26720 79200 26992
rect 800 26592 79200 26720
rect 800 26312 79120 26592
rect 800 26184 79200 26312
rect 880 25904 79200 26184
rect 800 25776 79200 25904
rect 800 25496 79120 25776
rect 800 25368 79200 25496
rect 880 25088 79200 25368
rect 800 24960 79200 25088
rect 800 24680 79120 24960
rect 800 24552 79200 24680
rect 880 24272 79200 24552
rect 800 24144 79200 24272
rect 800 23864 79120 24144
rect 800 23736 79200 23864
rect 880 23456 79200 23736
rect 800 23328 79200 23456
rect 800 23048 79120 23328
rect 800 22920 79200 23048
rect 880 22648 79200 22920
rect 880 22640 79120 22648
rect 800 22368 79120 22640
rect 800 22104 79200 22368
rect 880 21832 79200 22104
rect 880 21824 79120 21832
rect 800 21552 79120 21824
rect 800 21288 79200 21552
rect 880 21016 79200 21288
rect 880 21008 79120 21016
rect 800 20736 79120 21008
rect 800 20472 79200 20736
rect 880 20200 79200 20472
rect 880 20192 79120 20200
rect 800 19920 79120 20192
rect 800 19656 79200 19920
rect 880 19384 79200 19656
rect 880 19376 79120 19384
rect 800 19104 79120 19376
rect 800 18840 79200 19104
rect 880 18568 79200 18840
rect 880 18560 79120 18568
rect 800 18288 79120 18560
rect 800 17888 79200 18288
rect 880 17608 79120 17888
rect 800 17072 79200 17608
rect 880 16792 79120 17072
rect 800 16256 79200 16792
rect 880 15976 79120 16256
rect 800 15440 79200 15976
rect 880 15160 79120 15440
rect 800 14624 79200 15160
rect 880 14344 79120 14624
rect 800 13808 79200 14344
rect 880 13528 79120 13808
rect 800 13128 79200 13528
rect 800 12992 79120 13128
rect 880 12848 79120 12992
rect 880 12712 79200 12848
rect 800 12312 79200 12712
rect 800 12176 79120 12312
rect 880 12032 79120 12176
rect 880 11896 79200 12032
rect 800 11496 79200 11896
rect 800 11360 79120 11496
rect 880 11216 79120 11360
rect 880 11080 79200 11216
rect 800 10680 79200 11080
rect 800 10544 79120 10680
rect 880 10400 79120 10544
rect 880 10264 79200 10400
rect 800 9864 79200 10264
rect 800 9728 79120 9864
rect 880 9584 79120 9728
rect 880 9448 79200 9584
rect 800 9184 79200 9448
rect 800 8904 79120 9184
rect 800 8776 79200 8904
rect 880 8496 79200 8776
rect 800 8368 79200 8496
rect 800 8088 79120 8368
rect 800 7960 79200 8088
rect 880 7680 79200 7960
rect 800 7552 79200 7680
rect 800 7272 79120 7552
rect 800 7144 79200 7272
rect 880 6864 79200 7144
rect 800 6736 79200 6864
rect 800 6456 79120 6736
rect 800 6328 79200 6456
rect 880 6048 79200 6328
rect 800 5920 79200 6048
rect 800 5640 79120 5920
rect 800 5512 79200 5640
rect 880 5232 79200 5512
rect 800 5104 79200 5232
rect 800 4824 79120 5104
rect 800 4696 79200 4824
rect 880 4424 79200 4696
rect 880 4416 79120 4424
rect 800 4144 79120 4416
rect 800 3880 79200 4144
rect 880 3608 79200 3880
rect 880 3600 79120 3608
rect 800 3328 79120 3600
rect 800 3064 79200 3328
rect 880 2792 79200 3064
rect 880 2784 79120 2792
rect 800 2512 79120 2784
rect 800 2248 79200 2512
rect 880 1976 79200 2248
rect 880 1968 79120 1976
rect 800 1696 79120 1968
rect 800 1432 79200 1696
rect 880 1160 79200 1432
rect 880 1152 79120 1160
rect 800 880 79120 1152
rect 800 616 79200 880
rect 880 480 79200 616
rect 880 336 79120 480
rect 800 307 79120 336
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
<< obsm4 >>
rect 35387 110739 35453 124677
<< labels >>
rlabel metal3 s 0 10344 800 10464 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 103912 800 104032 6 addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 clk0
port 19 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 clk1
port 20 nsew signal output
rlabel metal2 s 1030 159200 1086 160000 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 3054 159200 3110 160000 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 5078 159200 5134 160000 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 7102 159200 7158 160000 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 9218 159200 9274 160000 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 11242 159200 11298 160000 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 13266 159200 13322 160000 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 15382 159200 15438 160000 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 79200 1776 80000 1896 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 79200 6536 80000 6656 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 79200 33464 80000 33584 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 79200 35776 80000 35896 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 79200 38224 80000 38344 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 79200 40536 80000 40656 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 79200 42984 80000 43104 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 79200 45296 80000 45416 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 79200 47744 80000 47864 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 79200 50056 80000 50176 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 79200 52504 80000 52624 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 79200 54816 80000 54936 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 79200 9664 80000 9784 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 79200 57264 80000 57384 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 79200 59576 80000 59696 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 79200 62024 80000 62144 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 79200 64336 80000 64456 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 79200 66784 80000 66904 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 79200 69096 80000 69216 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 79200 71408 80000 71528 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 79200 73856 80000 73976 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 79200 12928 80000 13048 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 79200 16056 80000 16176 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 79200 19184 80000 19304 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 79200 21632 80000 21752 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 79200 23944 80000 24064 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 79200 26392 80000 26512 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 79200 28704 80000 28824 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 79200 31152 80000 31272 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 79200 2592 80000 2712 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 79200 7352 80000 7472 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 79200 34280 80000 34400 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 79200 36592 80000 36712 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 79200 39040 80000 39160 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 79200 41352 80000 41472 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 79200 43800 80000 43920 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 79200 46112 80000 46232 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 79200 48560 80000 48680 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 79200 50872 80000 50992 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 79200 53320 80000 53440 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 79200 55632 80000 55752 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 79200 10480 80000 10600 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 79200 57944 80000 58064 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 79200 60392 80000 60512 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 79200 62704 80000 62824 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 79200 65152 80000 65272 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 79200 67464 80000 67584 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 79200 69912 80000 70032 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 79200 72224 80000 72344 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 79200 74672 80000 74792 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 79200 76168 80000 76288 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 79200 77800 80000 77920 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 79200 13608 80000 13728 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 79200 79432 80000 79552 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 79200 80928 80000 81048 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 79200 16872 80000 16992 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 79200 20000 80000 20120 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 79200 22448 80000 22568 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 79200 24760 80000 24880 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 79200 27072 80000 27192 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 79200 29520 80000 29640 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 79200 31832 80000 31952 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 79200 8168 80000 8288 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 79200 35096 80000 35216 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 79200 37408 80000 37528 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 79200 39856 80000 39976 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 79200 42168 80000 42288 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 79200 44616 80000 44736 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 79200 46928 80000 47048 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 79200 49240 80000 49360 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 79200 51688 80000 51808 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 79200 54000 80000 54120 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 79200 56448 80000 56568 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 79200 11296 80000 11416 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 79200 58760 80000 58880 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 79200 61208 80000 61328 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 79200 63520 80000 63640 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 79200 65968 80000 66088 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 79200 68280 80000 68400 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 79200 70728 80000 70848 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 79200 73040 80000 73160 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 79200 75488 80000 75608 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 79200 76984 80000 77104 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 79200 78616 80000 78736 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 79200 14424 80000 14544 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 79200 80248 80000 80368 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 79200 81744 80000 81864 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 79200 17688 80000 17808 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 79200 20816 80000 20936 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 79200 23128 80000 23248 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 79200 25576 80000 25696 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 79200 27888 80000 28008 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 79200 30336 80000 30456 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 79200 32648 80000 32768 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 79200 3408 80000 3528 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 79200 8984 80000 9104 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 79200 12112 80000 12232 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 79200 15240 80000 15360 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 79200 18368 80000 18488 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 79200 4224 80000 4344 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 79200 4904 80000 5024 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 79200 5720 80000 5840 6 core_wb_we_o
port 130 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 csb0[0]
port 131 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 csb0[1]
port 132 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 csb1[1]
port 134 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 din0[0]
port 135 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 din0[10]
port 136 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 din0[11]
port 137 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 din0[12]
port 138 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 din0[13]
port 139 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 din0[14]
port 140 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 din0[15]
port 141 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 din0[16]
port 142 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 din0[17]
port 143 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 din0[18]
port 144 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 din0[19]
port 145 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 din0[1]
port 146 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 din0[20]
port 147 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 din0[21]
port 148 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 din0[22]
port 149 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 din0[23]
port 150 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 din0[24]
port 151 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 din0[25]
port 152 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 din0[26]
port 153 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 din0[27]
port 154 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 din0[28]
port 155 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 din0[29]
port 156 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 din0[2]
port 157 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 din0[30]
port 158 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 din0[31]
port 159 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 din0[3]
port 160 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 din0[4]
port 161 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 din0[5]
port 162 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 din0[6]
port 163 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 din0[7]
port 164 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 din0[8]
port 165 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 din0[9]
port 166 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 dout0[0]
port 167 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 dout0[10]
port 168 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 dout0[11]
port 169 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 dout0[12]
port 170 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 dout0[13]
port 171 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 dout0[14]
port 172 nsew signal input
rlabel metal3 s 0 56720 800 56840 6 dout0[15]
port 173 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 dout0[16]
port 174 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 dout0[17]
port 175 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 dout0[18]
port 176 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 dout0[19]
port 177 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 dout0[1]
port 178 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 dout0[20]
port 179 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 dout0[21]
port 180 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 dout0[22]
port 181 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 dout0[23]
port 182 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 dout0[24]
port 183 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 dout0[25]
port 184 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 dout0[26]
port 185 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 dout0[27]
port 186 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 dout0[28]
port 187 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 dout0[29]
port 188 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 dout0[2]
port 189 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 dout0[30]
port 190 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 dout0[31]
port 191 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 dout0[32]
port 192 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 dout0[33]
port 193 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 dout0[34]
port 194 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 dout0[35]
port 195 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 dout0[36]
port 196 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 dout0[37]
port 197 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 dout0[38]
port 198 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 dout0[39]
port 199 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 dout0[3]
port 200 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 dout0[40]
port 201 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 dout0[41]
port 202 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 dout0[42]
port 203 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 dout0[43]
port 204 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 dout0[44]
port 205 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 dout0[45]
port 206 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 dout0[46]
port 207 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 dout0[47]
port 208 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 dout0[48]
port 209 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 dout0[49]
port 210 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 dout0[4]
port 211 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 dout0[50]
port 212 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 dout0[51]
port 213 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 dout0[52]
port 214 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 dout0[53]
port 215 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 dout0[54]
port 216 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 dout0[55]
port 217 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 dout0[56]
port 218 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 dout0[57]
port 219 nsew signal input
rlabel metal3 s 0 92352 800 92472 6 dout0[58]
port 220 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 dout0[59]
port 221 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 dout0[5]
port 222 nsew signal input
rlabel metal3 s 0 93984 800 94104 6 dout0[60]
port 223 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 dout0[61]
port 224 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 dout0[62]
port 225 nsew signal input
rlabel metal3 s 0 96432 800 96552 6 dout0[63]
port 226 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 dout0[6]
port 227 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 dout0[7]
port 228 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 dout0[8]
port 229 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 dout0[9]
port 230 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 dout1[0]
port 231 nsew signal input
rlabel metal3 s 0 115472 800 115592 6 dout1[10]
port 232 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 dout1[11]
port 233 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 dout1[12]
port 234 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 dout1[13]
port 235 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 dout1[14]
port 236 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 dout1[15]
port 237 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 dout1[16]
port 238 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 dout1[17]
port 239 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 dout1[18]
port 240 nsew signal input
rlabel metal3 s 0 122952 800 123072 6 dout1[19]
port 241 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 dout1[1]
port 242 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 dout1[20]
port 243 nsew signal input
rlabel metal3 s 0 124584 800 124704 6 dout1[21]
port 244 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 dout1[22]
port 245 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 dout1[23]
port 246 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 dout1[24]
port 247 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 dout1[25]
port 248 nsew signal input
rlabel metal3 s 0 128800 800 128920 6 dout1[26]
port 249 nsew signal input
rlabel metal3 s 0 129616 800 129736 6 dout1[27]
port 250 nsew signal input
rlabel metal3 s 0 130432 800 130552 6 dout1[28]
port 251 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 dout1[29]
port 252 nsew signal input
rlabel metal3 s 0 108944 800 109064 6 dout1[2]
port 253 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 dout1[30]
port 254 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 dout1[31]
port 255 nsew signal input
rlabel metal3 s 0 133832 800 133952 6 dout1[32]
port 256 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 dout1[33]
port 257 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 dout1[34]
port 258 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 dout1[35]
port 259 nsew signal input
rlabel metal3 s 0 137096 800 137216 6 dout1[36]
port 260 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 dout1[37]
port 261 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 dout1[38]
port 262 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 dout1[39]
port 263 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 dout1[3]
port 264 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 dout1[40]
port 265 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 dout1[41]
port 266 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 dout1[42]
port 267 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 dout1[43]
port 268 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 dout1[44]
port 269 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 dout1[45]
port 270 nsew signal input
rlabel metal3 s 0 145392 800 145512 6 dout1[46]
port 271 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 dout1[47]
port 272 nsew signal input
rlabel metal3 s 0 147024 800 147144 6 dout1[48]
port 273 nsew signal input
rlabel metal3 s 0 147840 800 147960 6 dout1[49]
port 274 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 dout1[4]
port 275 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 dout1[50]
port 276 nsew signal input
rlabel metal3 s 0 149472 800 149592 6 dout1[51]
port 277 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 dout1[52]
port 278 nsew signal input
rlabel metal3 s 0 151104 800 151224 6 dout1[53]
port 279 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 dout1[54]
port 280 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 dout1[55]
port 281 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 dout1[56]
port 282 nsew signal input
rlabel metal3 s 0 154504 800 154624 6 dout1[57]
port 283 nsew signal input
rlabel metal3 s 0 155320 800 155440 6 dout1[58]
port 284 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 dout1[59]
port 285 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 dout1[5]
port 286 nsew signal input
rlabel metal3 s 0 156952 800 157072 6 dout1[60]
port 287 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 dout1[61]
port 288 nsew signal input
rlabel metal3 s 0 158584 800 158704 6 dout1[62]
port 289 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 dout1[63]
port 290 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 dout1[6]
port 291 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 dout1[7]
port 292 nsew signal input
rlabel metal3 s 0 113840 800 113960 6 dout1[8]
port 293 nsew signal input
rlabel metal3 s 0 114656 800 114776 6 dout1[9]
port 294 nsew signal input
rlabel metal3 s 0 416 800 536 6 jtag_tck
port 295 nsew signal input
rlabel metal3 s 0 1232 800 1352 6 jtag_tdi
port 296 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 jtag_tdo
port 297 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 jtag_tms
port 298 nsew signal input
rlabel metal3 s 79200 82560 80000 82680 6 localMemory_wb_ack_o
port 299 nsew signal output
rlabel metal3 s 79200 87320 80000 87440 6 localMemory_wb_adr_i[0]
port 300 nsew signal input
rlabel metal3 s 79200 114248 80000 114368 6 localMemory_wb_adr_i[10]
port 301 nsew signal input
rlabel metal3 s 79200 116560 80000 116680 6 localMemory_wb_adr_i[11]
port 302 nsew signal input
rlabel metal3 s 79200 119008 80000 119128 6 localMemory_wb_adr_i[12]
port 303 nsew signal input
rlabel metal3 s 79200 121320 80000 121440 6 localMemory_wb_adr_i[13]
port 304 nsew signal input
rlabel metal3 s 79200 123768 80000 123888 6 localMemory_wb_adr_i[14]
port 305 nsew signal input
rlabel metal3 s 79200 126080 80000 126200 6 localMemory_wb_adr_i[15]
port 306 nsew signal input
rlabel metal3 s 79200 128528 80000 128648 6 localMemory_wb_adr_i[16]
port 307 nsew signal input
rlabel metal3 s 79200 130840 80000 130960 6 localMemory_wb_adr_i[17]
port 308 nsew signal input
rlabel metal3 s 79200 133288 80000 133408 6 localMemory_wb_adr_i[18]
port 309 nsew signal input
rlabel metal3 s 79200 135600 80000 135720 6 localMemory_wb_adr_i[19]
port 310 nsew signal input
rlabel metal3 s 79200 90448 80000 90568 6 localMemory_wb_adr_i[1]
port 311 nsew signal input
rlabel metal3 s 79200 137912 80000 138032 6 localMemory_wb_adr_i[20]
port 312 nsew signal input
rlabel metal3 s 79200 140360 80000 140480 6 localMemory_wb_adr_i[21]
port 313 nsew signal input
rlabel metal3 s 79200 142672 80000 142792 6 localMemory_wb_adr_i[22]
port 314 nsew signal input
rlabel metal3 s 79200 145120 80000 145240 6 localMemory_wb_adr_i[23]
port 315 nsew signal input
rlabel metal3 s 79200 93576 80000 93696 6 localMemory_wb_adr_i[2]
port 316 nsew signal input
rlabel metal3 s 79200 96840 80000 96960 6 localMemory_wb_adr_i[3]
port 317 nsew signal input
rlabel metal3 s 79200 99968 80000 100088 6 localMemory_wb_adr_i[4]
port 318 nsew signal input
rlabel metal3 s 79200 102416 80000 102536 6 localMemory_wb_adr_i[5]
port 319 nsew signal input
rlabel metal3 s 79200 104728 80000 104848 6 localMemory_wb_adr_i[6]
port 320 nsew signal input
rlabel metal3 s 79200 107040 80000 107160 6 localMemory_wb_adr_i[7]
port 321 nsew signal input
rlabel metal3 s 79200 109488 80000 109608 6 localMemory_wb_adr_i[8]
port 322 nsew signal input
rlabel metal3 s 79200 111800 80000 111920 6 localMemory_wb_adr_i[9]
port 323 nsew signal input
rlabel metal3 s 79200 83376 80000 83496 6 localMemory_wb_cyc_i
port 324 nsew signal input
rlabel metal3 s 79200 88136 80000 88256 6 localMemory_wb_data_i[0]
port 325 nsew signal input
rlabel metal3 s 79200 115064 80000 115184 6 localMemory_wb_data_i[10]
port 326 nsew signal input
rlabel metal3 s 79200 117376 80000 117496 6 localMemory_wb_data_i[11]
port 327 nsew signal input
rlabel metal3 s 79200 119824 80000 119944 6 localMemory_wb_data_i[12]
port 328 nsew signal input
rlabel metal3 s 79200 122136 80000 122256 6 localMemory_wb_data_i[13]
port 329 nsew signal input
rlabel metal3 s 79200 124584 80000 124704 6 localMemory_wb_data_i[14]
port 330 nsew signal input
rlabel metal3 s 79200 126896 80000 127016 6 localMemory_wb_data_i[15]
port 331 nsew signal input
rlabel metal3 s 79200 129208 80000 129328 6 localMemory_wb_data_i[16]
port 332 nsew signal input
rlabel metal3 s 79200 131656 80000 131776 6 localMemory_wb_data_i[17]
port 333 nsew signal input
rlabel metal3 s 79200 133968 80000 134088 6 localMemory_wb_data_i[18]
port 334 nsew signal input
rlabel metal3 s 79200 136416 80000 136536 6 localMemory_wb_data_i[19]
port 335 nsew signal input
rlabel metal3 s 79200 91264 80000 91384 6 localMemory_wb_data_i[1]
port 336 nsew signal input
rlabel metal3 s 79200 138728 80000 138848 6 localMemory_wb_data_i[20]
port 337 nsew signal input
rlabel metal3 s 79200 141176 80000 141296 6 localMemory_wb_data_i[21]
port 338 nsew signal input
rlabel metal3 s 79200 143488 80000 143608 6 localMemory_wb_data_i[22]
port 339 nsew signal input
rlabel metal3 s 79200 145936 80000 146056 6 localMemory_wb_data_i[23]
port 340 nsew signal input
rlabel metal3 s 79200 147432 80000 147552 6 localMemory_wb_data_i[24]
port 341 nsew signal input
rlabel metal3 s 79200 149064 80000 149184 6 localMemory_wb_data_i[25]
port 342 nsew signal input
rlabel metal3 s 79200 150696 80000 150816 6 localMemory_wb_data_i[26]
port 343 nsew signal input
rlabel metal3 s 79200 152192 80000 152312 6 localMemory_wb_data_i[27]
port 344 nsew signal input
rlabel metal3 s 79200 153824 80000 153944 6 localMemory_wb_data_i[28]
port 345 nsew signal input
rlabel metal3 s 79200 155456 80000 155576 6 localMemory_wb_data_i[29]
port 346 nsew signal input
rlabel metal3 s 79200 94392 80000 94512 6 localMemory_wb_data_i[2]
port 347 nsew signal input
rlabel metal3 s 79200 156952 80000 157072 6 localMemory_wb_data_i[30]
port 348 nsew signal input
rlabel metal3 s 79200 158584 80000 158704 6 localMemory_wb_data_i[31]
port 349 nsew signal input
rlabel metal3 s 79200 97656 80000 97776 6 localMemory_wb_data_i[3]
port 350 nsew signal input
rlabel metal3 s 79200 100784 80000 100904 6 localMemory_wb_data_i[4]
port 351 nsew signal input
rlabel metal3 s 79200 103096 80000 103216 6 localMemory_wb_data_i[5]
port 352 nsew signal input
rlabel metal3 s 79200 105544 80000 105664 6 localMemory_wb_data_i[6]
port 353 nsew signal input
rlabel metal3 s 79200 107856 80000 107976 6 localMemory_wb_data_i[7]
port 354 nsew signal input
rlabel metal3 s 79200 110304 80000 110424 6 localMemory_wb_data_i[8]
port 355 nsew signal input
rlabel metal3 s 79200 112616 80000 112736 6 localMemory_wb_data_i[9]
port 356 nsew signal input
rlabel metal3 s 79200 88952 80000 89072 6 localMemory_wb_data_o[0]
port 357 nsew signal output
rlabel metal3 s 79200 115744 80000 115864 6 localMemory_wb_data_o[10]
port 358 nsew signal output
rlabel metal3 s 79200 118192 80000 118312 6 localMemory_wb_data_o[11]
port 359 nsew signal output
rlabel metal3 s 79200 120504 80000 120624 6 localMemory_wb_data_o[12]
port 360 nsew signal output
rlabel metal3 s 79200 122952 80000 123072 6 localMemory_wb_data_o[13]
port 361 nsew signal output
rlabel metal3 s 79200 125264 80000 125384 6 localMemory_wb_data_o[14]
port 362 nsew signal output
rlabel metal3 s 79200 127712 80000 127832 6 localMemory_wb_data_o[15]
port 363 nsew signal output
rlabel metal3 s 79200 130024 80000 130144 6 localMemory_wb_data_o[16]
port 364 nsew signal output
rlabel metal3 s 79200 132472 80000 132592 6 localMemory_wb_data_o[17]
port 365 nsew signal output
rlabel metal3 s 79200 134784 80000 134904 6 localMemory_wb_data_o[18]
port 366 nsew signal output
rlabel metal3 s 79200 137232 80000 137352 6 localMemory_wb_data_o[19]
port 367 nsew signal output
rlabel metal3 s 79200 92080 80000 92200 6 localMemory_wb_data_o[1]
port 368 nsew signal output
rlabel metal3 s 79200 139544 80000 139664 6 localMemory_wb_data_o[20]
port 369 nsew signal output
rlabel metal3 s 79200 141992 80000 142112 6 localMemory_wb_data_o[21]
port 370 nsew signal output
rlabel metal3 s 79200 144304 80000 144424 6 localMemory_wb_data_o[22]
port 371 nsew signal output
rlabel metal3 s 79200 146752 80000 146872 6 localMemory_wb_data_o[23]
port 372 nsew signal output
rlabel metal3 s 79200 148248 80000 148368 6 localMemory_wb_data_o[24]
port 373 nsew signal output
rlabel metal3 s 79200 149880 80000 150000 6 localMemory_wb_data_o[25]
port 374 nsew signal output
rlabel metal3 s 79200 151376 80000 151496 6 localMemory_wb_data_o[26]
port 375 nsew signal output
rlabel metal3 s 79200 153008 80000 153128 6 localMemory_wb_data_o[27]
port 376 nsew signal output
rlabel metal3 s 79200 154640 80000 154760 6 localMemory_wb_data_o[28]
port 377 nsew signal output
rlabel metal3 s 79200 156136 80000 156256 6 localMemory_wb_data_o[29]
port 378 nsew signal output
rlabel metal3 s 79200 95208 80000 95328 6 localMemory_wb_data_o[2]
port 379 nsew signal output
rlabel metal3 s 79200 157768 80000 157888 6 localMemory_wb_data_o[30]
port 380 nsew signal output
rlabel metal3 s 79200 159400 80000 159520 6 localMemory_wb_data_o[31]
port 381 nsew signal output
rlabel metal3 s 79200 98336 80000 98456 6 localMemory_wb_data_o[3]
port 382 nsew signal output
rlabel metal3 s 79200 101600 80000 101720 6 localMemory_wb_data_o[4]
port 383 nsew signal output
rlabel metal3 s 79200 103912 80000 104032 6 localMemory_wb_data_o[5]
port 384 nsew signal output
rlabel metal3 s 79200 106360 80000 106480 6 localMemory_wb_data_o[6]
port 385 nsew signal output
rlabel metal3 s 79200 108672 80000 108792 6 localMemory_wb_data_o[7]
port 386 nsew signal output
rlabel metal3 s 79200 111120 80000 111240 6 localMemory_wb_data_o[8]
port 387 nsew signal output
rlabel metal3 s 79200 113432 80000 113552 6 localMemory_wb_data_o[9]
port 388 nsew signal output
rlabel metal3 s 79200 84192 80000 84312 6 localMemory_wb_error_o
port 389 nsew signal output
rlabel metal3 s 79200 89632 80000 89752 6 localMemory_wb_sel_i[0]
port 390 nsew signal input
rlabel metal3 s 79200 92896 80000 93016 6 localMemory_wb_sel_i[1]
port 391 nsew signal input
rlabel metal3 s 79200 96024 80000 96144 6 localMemory_wb_sel_i[2]
port 392 nsew signal input
rlabel metal3 s 79200 99152 80000 99272 6 localMemory_wb_sel_i[3]
port 393 nsew signal input
rlabel metal3 s 79200 84872 80000 84992 6 localMemory_wb_stall_o
port 394 nsew signal output
rlabel metal3 s 79200 85688 80000 85808 6 localMemory_wb_stb_i
port 395 nsew signal input
rlabel metal3 s 79200 86504 80000 86624 6 localMemory_wb_we_i
port 396 nsew signal input
rlabel metal2 s 17406 159200 17462 160000 6 manufacturerID[0]
port 397 nsew signal input
rlabel metal2 s 37922 159200 37978 160000 6 manufacturerID[10]
port 398 nsew signal input
rlabel metal2 s 19430 159200 19486 160000 6 manufacturerID[1]
port 399 nsew signal input
rlabel metal2 s 21546 159200 21602 160000 6 manufacturerID[2]
port 400 nsew signal input
rlabel metal2 s 23570 159200 23626 160000 6 manufacturerID[3]
port 401 nsew signal input
rlabel metal2 s 25594 159200 25650 160000 6 manufacturerID[4]
port 402 nsew signal input
rlabel metal2 s 27710 159200 27766 160000 6 manufacturerID[5]
port 403 nsew signal input
rlabel metal2 s 29734 159200 29790 160000 6 manufacturerID[6]
port 404 nsew signal input
rlabel metal2 s 31758 159200 31814 160000 6 manufacturerID[7]
port 405 nsew signal input
rlabel metal2 s 33782 159200 33838 160000 6 manufacturerID[8]
port 406 nsew signal input
rlabel metal2 s 35898 159200 35954 160000 6 manufacturerID[9]
port 407 nsew signal input
rlabel metal2 s 39946 159200 40002 160000 6 partID[0]
port 408 nsew signal input
rlabel metal2 s 60462 159200 60518 160000 6 partID[10]
port 409 nsew signal input
rlabel metal2 s 62578 159200 62634 160000 6 partID[11]
port 410 nsew signal input
rlabel metal2 s 64602 159200 64658 160000 6 partID[12]
port 411 nsew signal input
rlabel metal2 s 66626 159200 66682 160000 6 partID[13]
port 412 nsew signal input
rlabel metal2 s 68742 159200 68798 160000 6 partID[14]
port 413 nsew signal input
rlabel metal2 s 70766 159200 70822 160000 6 partID[15]
port 414 nsew signal input
rlabel metal2 s 42062 159200 42118 160000 6 partID[1]
port 415 nsew signal input
rlabel metal2 s 44086 159200 44142 160000 6 partID[2]
port 416 nsew signal input
rlabel metal2 s 46110 159200 46166 160000 6 partID[3]
port 417 nsew signal input
rlabel metal2 s 48226 159200 48282 160000 6 partID[4]
port 418 nsew signal input
rlabel metal2 s 50250 159200 50306 160000 6 partID[5]
port 419 nsew signal input
rlabel metal2 s 52274 159200 52330 160000 6 partID[6]
port 420 nsew signal input
rlabel metal2 s 54390 159200 54446 160000 6 partID[7]
port 421 nsew signal input
rlabel metal2 s 56414 159200 56470 160000 6 partID[8]
port 422 nsew signal input
rlabel metal2 s 58438 159200 58494 160000 6 partID[9]
port 423 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 probe_errorCode[0]
port 424 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 probe_errorCode[1]
port 425 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 probe_errorCode[2]
port 426 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 probe_errorCode[3]
port 427 nsew signal output
rlabel metal2 s 662 0 718 800 6 probe_isBranch
port 428 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 probe_isCompressed
port 429 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 probe_isLoad
port 430 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 probe_isStore
port 431 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 probe_jtagInstruction[0]
port 432 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 probe_jtagInstruction[1]
port 433 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 probe_jtagInstruction[2]
port 434 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 probe_jtagInstruction[3]
port 435 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 probe_jtagInstruction[4]
port 436 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 probe_opcode[0]
port 437 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 probe_opcode[1]
port 438 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 probe_opcode[2]
port 439 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 probe_opcode[3]
port 440 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 probe_opcode[4]
port 441 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 probe_opcode[5]
port 442 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 probe_opcode[6]
port 443 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 probe_programCounter[0]
port 444 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 probe_programCounter[10]
port 445 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 probe_programCounter[11]
port 446 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 probe_programCounter[12]
port 447 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 probe_programCounter[13]
port 448 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 probe_programCounter[14]
port 449 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 probe_programCounter[15]
port 450 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 probe_programCounter[16]
port 451 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 probe_programCounter[17]
port 452 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 probe_programCounter[18]
port 453 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 probe_programCounter[19]
port 454 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 probe_programCounter[1]
port 455 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 probe_programCounter[20]
port 456 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 probe_programCounter[21]
port 457 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 probe_programCounter[22]
port 458 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 probe_programCounter[23]
port 459 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 probe_programCounter[24]
port 460 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 probe_programCounter[25]
port 461 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 probe_programCounter[26]
port 462 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 probe_programCounter[27]
port 463 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 probe_programCounter[28]
port 464 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 probe_programCounter[29]
port 465 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 probe_programCounter[2]
port 466 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 probe_programCounter[30]
port 467 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 probe_programCounter[31]
port 468 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 probe_programCounter[3]
port 469 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 probe_programCounter[4]
port 470 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 probe_programCounter[5]
port 471 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 probe_programCounter[6]
port 472 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 probe_programCounter[7]
port 473 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 probe_programCounter[8]
port 474 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 probe_programCounter[9]
port 475 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 probe_state[0]
port 476 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 probe_state[1]
port 477 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 probe_takeBranch
port 478 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 479 nsew power bidirectional
rlabel metal2 s 72790 159200 72846 160000 6 versionID[0]
port 480 nsew signal input
rlabel metal2 s 74906 159200 74962 160000 6 versionID[1]
port 481 nsew signal input
rlabel metal2 s 76930 159200 76986 160000 6 versionID[2]
port 482 nsew signal input
rlabel metal2 s 78954 159200 79010 160000 6 versionID[3]
port 483 nsew signal input
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 484 nsew ground bidirectional
rlabel metal3 s 79200 280 80000 400 6 wb_clk_i
port 485 nsew signal input
rlabel metal3 s 79200 960 80000 1080 6 wb_rst_i
port 486 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 web0
port 487 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 wmask0[0]
port 488 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 wmask0[1]
port 489 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 wmask0[2]
port 490 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 wmask0[3]
port 491 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6182128
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/signoff/ExperiarCore.magic.gds
string GDS_START 518744
<< end >>

