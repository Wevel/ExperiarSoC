// This is the unpowered netlist.
module Flash (flash_csb,
    flash_io0_read,
    flash_io0_we,
    flash_io0_write,
    flash_io1_read,
    flash_io1_we,
    flash_io1_write,
    flash_sck,
    sram_clk0,
    sram_clk1,
    sram_csb0,
    sram_csb1,
    sram_web0,
    wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_error_o,
    wb_rst_i,
    wb_stall_o,
    wb_stb_i,
    wb_we_i,
    sram_addr0,
    sram_addr1,
    sram_din0,
    sram_dout0,
    sram_dout1,
    sram_wmask0,
    wb_adr_i,
    wb_data_i,
    wb_data_o,
    wb_sel_i);
 output flash_csb;
 input flash_io0_read;
 output flash_io0_we;
 output flash_io0_write;
 input flash_io1_read;
 output flash_io1_we;
 output flash_io1_write;
 output flash_sck;
 output sram_clk0;
 output sram_clk1;
 output sram_csb0;
 output sram_csb1;
 output sram_web0;
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 output wb_error_o;
 input wb_rst_i;
 output wb_stall_o;
 input wb_stb_i;
 input wb_we_i;
 output [8:0] sram_addr0;
 output [8:0] sram_addr1;
 output [31:0] sram_din0;
 input [31:0] sram_dout0;
 input [31:0] sram_dout1;
 output [3:0] sram_wmask0;
 input [23:0] wb_adr_i;
 input [31:0] wb_data_i;
 output [31:0] wb_data_o;
 input [3:0] wb_sel_i;

 wire net242;
 wire net238;
 wire net239;
 wire net240;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net241;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire \flashBuffer.baseAddress[0] ;
 wire \flashBuffer.baseAddress[10] ;
 wire \flashBuffer.baseAddress[11] ;
 wire \flashBuffer.baseAddress[12] ;
 wire \flashBuffer.baseAddress[13] ;
 wire \flashBuffer.baseAddress[14] ;
 wire \flashBuffer.baseAddress[15] ;
 wire \flashBuffer.baseAddress[16] ;
 wire \flashBuffer.baseAddress[17] ;
 wire \flashBuffer.baseAddress[18] ;
 wire \flashBuffer.baseAddress[19] ;
 wire \flashBuffer.baseAddress[1] ;
 wire \flashBuffer.baseAddress[20] ;
 wire \flashBuffer.baseAddress[21] ;
 wire \flashBuffer.baseAddress[22] ;
 wire \flashBuffer.baseAddress[23] ;
 wire \flashBuffer.baseAddress[2] ;
 wire \flashBuffer.baseAddress[3] ;
 wire \flashBuffer.baseAddress[4] ;
 wire \flashBuffer.baseAddress[5] ;
 wire \flashBuffer.baseAddress[6] ;
 wire \flashBuffer.baseAddress[7] ;
 wire \flashBuffer.baseAddress[8] ;
 wire \flashBuffer.baseAddress[9] ;
 wire \flashBuffer.cachedAddress[11] ;
 wire \flashBuffer.cachedAddress[12] ;
 wire \flashBuffer.cachedAddress[13] ;
 wire \flashBuffer.cachedAddress[14] ;
 wire \flashBuffer.cachedAddress[15] ;
 wire \flashBuffer.cachedAddress[16] ;
 wire \flashBuffer.cachedAddress[17] ;
 wire \flashBuffer.cachedAddress[18] ;
 wire \flashBuffer.cachedAddress[19] ;
 wire \flashBuffer.cachedAddress[20] ;
 wire \flashBuffer.cachedAddress[21] ;
 wire \flashBuffer.cachedAddress[22] ;
 wire \flashBuffer.cachedAddress[23] ;
 wire \flashBuffer.cachedCount[0] ;
 wire \flashBuffer.cachedCount[1] ;
 wire \flashBuffer.cachedCount[2] ;
 wire \flashBuffer.cachedCount[3] ;
 wire \flashBuffer.cachedCount[4] ;
 wire \flashBuffer.cachedCount[5] ;
 wire \flashBuffer.cachedCount[6] ;
 wire \flashBuffer.cachedCount[7] ;
 wire \flashBuffer.cachedCount[8] ;
 wire \flashBuffer.cachedCount[9] ;
 wire \flashBuffer.configuration ;
 wire \flashBuffer.flashCacheReadReady ;
 wire \flashBuffer.qspi_readDataValid ;
 wire \flashBuffer.qspi_requestData ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \qspiDevice.bitCounter[0] ;
 wire \qspiDevice.bitCounter[1] ;
 wire \qspiDevice.bitCounter[2] ;
 wire \qspiDevice.bitCounter[3] ;
 wire \qspiDevice.bitCounter[4] ;
 wire \qspiDevice.outputClock ;
 wire \qspiDevice.register.outputBit ;
 wire \qspiDevice.resetState[0] ;
 wire \qspiDevice.resetState[1] ;
 wire \qspiDevice.settingAddress ;
 wire \qspiDevice.state[0] ;
 wire \qspiDevice.state[1] ;
 wire \wbPeripheralBusInterface.currentAddress[10] ;
 wire \wbPeripheralBusInterface.currentAddress[11] ;
 wire \wbPeripheralBusInterface.currentAddress[12] ;
 wire \wbPeripheralBusInterface.currentAddress[13] ;
 wire \wbPeripheralBusInterface.currentAddress[14] ;
 wire \wbPeripheralBusInterface.currentAddress[15] ;
 wire \wbPeripheralBusInterface.currentAddress[16] ;
 wire \wbPeripheralBusInterface.currentAddress[17] ;
 wire \wbPeripheralBusInterface.currentAddress[18] ;
 wire \wbPeripheralBusInterface.currentAddress[19] ;
 wire \wbPeripheralBusInterface.currentAddress[20] ;
 wire \wbPeripheralBusInterface.currentAddress[21] ;
 wire \wbPeripheralBusInterface.currentAddress[22] ;
 wire \wbPeripheralBusInterface.currentAddress[23] ;
 wire \wbPeripheralBusInterface.currentAddress[2] ;
 wire \wbPeripheralBusInterface.currentAddress[3] ;
 wire \wbPeripheralBusInterface.currentAddress[4] ;
 wire \wbPeripheralBusInterface.currentAddress[5] ;
 wire \wbPeripheralBusInterface.currentAddress[6] ;
 wire \wbPeripheralBusInterface.currentAddress[7] ;
 wire \wbPeripheralBusInterface.currentAddress[8] ;
 wire \wbPeripheralBusInterface.currentAddress[9] ;
 wire \wbPeripheralBusInterface.currentByteSelect[0] ;
 wire \wbPeripheralBusInterface.currentByteSelect[1] ;
 wire \wbPeripheralBusInterface.currentByteSelect[2] ;
 wire \wbPeripheralBusInterface.state[0] ;
 wire \wbPeripheralBusInterface.state[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net58));
 sky130_fd_sc_hd__decap_4 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_94 ();
 sky130_fd_sc_hd__conb_1 Flash_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 Flash_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 Flash_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 Flash_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 Flash_242 (.HI(net242));
 sky130_fd_sc_hd__conb_1 Flash_243 (.HI(net243));
 sky130_fd_sc_hd__conb_1 Flash_244 (.HI(net244));
 sky130_fd_sc_hd__conb_1 Flash_245 (.HI(net245));
 sky130_fd_sc_hd__conb_1 Flash_246 (.HI(net246));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__clkinv_2 _0475_ (.A(\wbPeripheralBusInterface.state[0] ),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _0476_ (.A(\flashBuffer.cachedAddress[11] ),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _0477_ (.A(\qspiDevice.bitCounter[4] ),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(\qspiDevice.bitCounter[0] ),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\flashBuffer.qspi_readDataValid ),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _0480_ (.A(net226),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _0481_ (.A(\qspiDevice.resetState[1] ),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _0482_ (.A(\flashBuffer.cachedCount[8] ),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _0483_ (.A(\flashBuffer.cachedCount[7] ),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _0484_ (.A(\wbPeripheralBusInterface.currentAddress[3] ),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(net237),
    .Y(_0176_));
 sky130_fd_sc_hd__nor2_4 _0486_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .Y(_0177_));
 sky130_fd_sc_hd__or2_2 _0487_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .X(_0178_));
 sky130_fd_sc_hd__nor2_1 _0488_ (.A(_0175_),
    .B(_0177_),
    .Y(net100));
 sky130_fd_sc_hd__and2_2 _0489_ (.A(\wbPeripheralBusInterface.currentAddress[2] ),
    .B(net220),
    .X(net99));
 sky130_fd_sc_hd__nand2_4 _0490_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(_0166_),
    .Y(_0179_));
 sky130_fd_sc_hd__or4_1 _0491_ (.A(\wbPeripheralBusInterface.currentAddress[11] ),
    .B(\wbPeripheralBusInterface.currentAddress[19] ),
    .C(\wbPeripheralBusInterface.currentAddress[21] ),
    .D(\wbPeripheralBusInterface.currentAddress[22] ),
    .X(_0180_));
 sky130_fd_sc_hd__o31a_1 _0492_ (.A1(\wbPeripheralBusInterface.currentAddress[20] ),
    .A2(\wbPeripheralBusInterface.currentAddress[23] ),
    .A3(_0180_),
    .B1(net221),
    .X(_0181_));
 sky130_fd_sc_hd__or4_1 _0493_ (.A(\wbPeripheralBusInterface.currentAddress[15] ),
    .B(\wbPeripheralBusInterface.currentAddress[16] ),
    .C(\wbPeripheralBusInterface.currentAddress[17] ),
    .D(\wbPeripheralBusInterface.currentAddress[18] ),
    .X(_0182_));
 sky130_fd_sc_hd__or3_1 _0494_ (.A(\wbPeripheralBusInterface.currentAddress[13] ),
    .B(\wbPeripheralBusInterface.currentAddress[14] ),
    .C(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__or4_4 _0495_ (.A(\wbPeripheralBusInterface.currentAddress[12] ),
    .B(_0179_),
    .C(_0181_),
    .D(_0183_),
    .X(net111));
 sky130_fd_sc_hd__nor2_8 _0496_ (.A(net226),
    .B(\qspiDevice.state[0] ),
    .Y(net87));
 sky130_fd_sc_hd__and2_1 _0497_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(net220),
    .X(net101));
 sky130_fd_sc_hd__and2_1 _0498_ (.A(\wbPeripheralBusInterface.currentAddress[5] ),
    .B(net220),
    .X(net102));
 sky130_fd_sc_hd__and2_1 _0499_ (.A(\wbPeripheralBusInterface.currentAddress[6] ),
    .B(net220),
    .X(net103));
 sky130_fd_sc_hd__and2_1 _0500_ (.A(\wbPeripheralBusInterface.currentAddress[7] ),
    .B(net220),
    .X(net104));
 sky130_fd_sc_hd__and2_1 _0501_ (.A(\wbPeripheralBusInterface.currentAddress[8] ),
    .B(net221),
    .X(net105));
 sky130_fd_sc_hd__and2_1 _0502_ (.A(\wbPeripheralBusInterface.currentAddress[9] ),
    .B(net221),
    .X(net106));
 sky130_fd_sc_hd__and2_1 _0503_ (.A(\wbPeripheralBusInterface.currentAddress[10] ),
    .B(net220),
    .X(net107));
 sky130_fd_sc_hd__and2_2 _0504_ (.A(\flashBuffer.qspi_readDataValid ),
    .B(\flashBuffer.qspi_requestData ),
    .X(_0184_));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(_0184_),
    .Y(net110));
 sky130_fd_sc_hd__o21a_1 _0506_ (.A1(net226),
    .A2(net227),
    .B1(\qspiDevice.register.outputBit ),
    .X(net88));
 sky130_fd_sc_hd__and4_1 _0507_ (.A(\flashBuffer.cachedCount[5] ),
    .B(\flashBuffer.cachedCount[4] ),
    .C(\flashBuffer.cachedCount[3] ),
    .D(\flashBuffer.cachedCount[0] ),
    .X(_0185_));
 sky130_fd_sc_hd__and4_1 _0508_ (.A(\flashBuffer.cachedCount[7] ),
    .B(\flashBuffer.cachedCount[6] ),
    .C(\flashBuffer.cachedCount[2] ),
    .D(\flashBuffer.cachedCount[1] ),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_1 _0509_ (.A(_0185_),
    .B(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__o41a_1 _0510_ (.A1(_0170_),
    .A2(\flashBuffer.cachedCount[9] ),
    .A3(_0173_),
    .A4(_0187_),
    .B1(\flashBuffer.qspi_requestData ),
    .X(_0188_));
 sky130_fd_sc_hd__or3_1 _0511_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(\wbPeripheralBusInterface.currentAddress[5] ),
    .C(\wbPeripheralBusInterface.currentAddress[10] ),
    .X(_0189_));
 sky130_fd_sc_hd__o41a_1 _0512_ (.A1(\wbPeripheralBusInterface.currentAddress[6] ),
    .A2(\wbPeripheralBusInterface.currentAddress[7] ),
    .A3(\wbPeripheralBusInterface.currentAddress[8] ),
    .A4(\wbPeripheralBusInterface.currentAddress[9] ),
    .B1(net221),
    .X(_0190_));
 sky130_fd_sc_hd__or3b_4 _0513_ (.A(_0190_),
    .B(\wbPeripheralBusInterface.currentAddress[3] ),
    .C_N(net99),
    .X(_0191_));
 sky130_fd_sc_hd__or4_1 _0514_ (.A(\wbPeripheralBusInterface.currentAddress[14] ),
    .B(\wbPeripheralBusInterface.currentAddress[15] ),
    .C(\wbPeripheralBusInterface.currentAddress[17] ),
    .D(\wbPeripheralBusInterface.currentAddress[18] ),
    .X(_0192_));
 sky130_fd_sc_hd__or4b_1 _0515_ (.A(\wbPeripheralBusInterface.currentAddress[13] ),
    .B(\wbPeripheralBusInterface.currentAddress[16] ),
    .C(\wbPeripheralBusInterface.currentAddress[19] ),
    .D_N(\wbPeripheralBusInterface.currentAddress[12] ),
    .X(_0193_));
 sky130_fd_sc_hd__or3_1 _0516_ (.A(_0177_),
    .B(_0189_),
    .C(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__or3_4 _0517_ (.A(_0181_),
    .B(_0192_),
    .C(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__nor4_1 _0518_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(_0166_),
    .C(_0191_),
    .D(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__o21a_1 _0519_ (.A1(_0188_),
    .A2(net205),
    .B1(net229),
    .X(_0000_));
 sky130_fd_sc_hd__nor2_4 _0520_ (.A(net237),
    .B(net205),
    .Y(_0197_));
 sky130_fd_sc_hd__or2_4 _0521_ (.A(net237),
    .B(net208),
    .X(_0198_));
 sky130_fd_sc_hd__a21oi_1 _0522_ (.A1(\flashBuffer.cachedCount[0] ),
    .A2(_0184_),
    .B1(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__o21a_1 _0523_ (.A1(\flashBuffer.cachedCount[0] ),
    .A2(_0184_),
    .B1(_0199_),
    .X(_0001_));
 sky130_fd_sc_hd__a31o_1 _0524_ (.A1(\flashBuffer.qspi_readDataValid ),
    .A2(\flashBuffer.cachedCount[0] ),
    .A3(\flashBuffer.qspi_requestData ),
    .B1(\flashBuffer.cachedCount[1] ),
    .X(_0200_));
 sky130_fd_sc_hd__and3_1 _0525_ (.A(\flashBuffer.cachedCount[1] ),
    .B(\flashBuffer.cachedCount[0] ),
    .C(_0184_),
    .X(_0201_));
 sky130_fd_sc_hd__and3b_1 _0526_ (.A_N(_0201_),
    .B(net196),
    .C(_0200_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _0527_ (.A(\flashBuffer.cachedCount[2] ),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__o21ai_1 _0528_ (.A1(\flashBuffer.cachedCount[2] ),
    .A2(_0201_),
    .B1(net196),
    .Y(_0203_));
 sky130_fd_sc_hd__nor2_1 _0529_ (.A(_0202_),
    .B(_0203_),
    .Y(_0003_));
 sky130_fd_sc_hd__and3_2 _0530_ (.A(\flashBuffer.cachedCount[3] ),
    .B(\flashBuffer.cachedCount[2] ),
    .C(_0201_),
    .X(_0204_));
 sky130_fd_sc_hd__o21ai_1 _0531_ (.A1(\flashBuffer.cachedCount[3] ),
    .A2(_0202_),
    .B1(net196),
    .Y(_0205_));
 sky130_fd_sc_hd__nor2_1 _0532_ (.A(_0204_),
    .B(_0205_),
    .Y(_0004_));
 sky130_fd_sc_hd__and2_2 _0533_ (.A(\flashBuffer.cachedCount[4] ),
    .B(_0204_),
    .X(_0206_));
 sky130_fd_sc_hd__o21ai_1 _0534_ (.A1(\flashBuffer.cachedCount[4] ),
    .A2(_0204_),
    .B1(net196),
    .Y(_0207_));
 sky130_fd_sc_hd__nor2_1 _0535_ (.A(_0206_),
    .B(_0207_),
    .Y(_0005_));
 sky130_fd_sc_hd__o21ai_1 _0536_ (.A1(\flashBuffer.cachedCount[5] ),
    .A2(_0206_),
    .B1(net196),
    .Y(_0208_));
 sky130_fd_sc_hd__a21oi_1 _0537_ (.A1(\flashBuffer.cachedCount[5] ),
    .A2(_0206_),
    .B1(_0208_),
    .Y(_0006_));
 sky130_fd_sc_hd__nand3_1 _0538_ (.A(\flashBuffer.cachedCount[6] ),
    .B(\flashBuffer.cachedCount[5] ),
    .C(_0206_),
    .Y(_0209_));
 sky130_fd_sc_hd__a31o_1 _0539_ (.A1(\flashBuffer.cachedCount[5] ),
    .A2(\flashBuffer.cachedCount[4] ),
    .A3(_0204_),
    .B1(\flashBuffer.cachedCount[6] ),
    .X(_0210_));
 sky130_fd_sc_hd__and3_1 _0540_ (.A(net196),
    .B(_0209_),
    .C(_0210_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_1 _0541_ (.A(net110),
    .B(_0187_),
    .Y(_0211_));
 sky130_fd_sc_hd__a211oi_1 _0542_ (.A1(_0174_),
    .A2(_0209_),
    .B1(_0211_),
    .C1(_0198_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_1 _0543_ (.A(\flashBuffer.cachedCount[8] ),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__or2_1 _0544_ (.A(\flashBuffer.cachedCount[8] ),
    .B(_0211_),
    .X(_0213_));
 sky130_fd_sc_hd__and3_1 _0545_ (.A(net196),
    .B(_0212_),
    .C(_0213_),
    .X(_0009_));
 sky130_fd_sc_hd__xor2_1 _0546_ (.A(\flashBuffer.cachedCount[9] ),
    .B(_0212_),
    .X(_0214_));
 sky130_fd_sc_hd__nor2_1 _0547_ (.A(_0198_),
    .B(_0214_),
    .Y(_0010_));
 sky130_fd_sc_hd__and3_1 _0548_ (.A(net228),
    .B(net57),
    .C(net204),
    .X(_0215_));
 sky130_fd_sc_hd__a21o_1 _0549_ (.A1(\flashBuffer.baseAddress[0] ),
    .A2(net195),
    .B1(_0215_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _0550_ (.A(net228),
    .B(net68),
    .C(net204),
    .X(_0216_));
 sky130_fd_sc_hd__a21o_1 _0551_ (.A1(\flashBuffer.baseAddress[1] ),
    .A2(net195),
    .B1(_0216_),
    .X(_0012_));
 sky130_fd_sc_hd__and3_4 _0552_ (.A(net228),
    .B(net73),
    .C(net204),
    .X(_0217_));
 sky130_fd_sc_hd__a21o_1 _0553_ (.A1(\flashBuffer.baseAddress[2] ),
    .A2(net195),
    .B1(_0217_),
    .X(_0013_));
 sky130_fd_sc_hd__and3_4 _0554_ (.A(net228),
    .B(net74),
    .C(net204),
    .X(_0218_));
 sky130_fd_sc_hd__a21o_1 _0555_ (.A1(\flashBuffer.baseAddress[3] ),
    .A2(net195),
    .B1(_0218_),
    .X(_0014_));
 sky130_fd_sc_hd__and3_4 _0556_ (.A(net228),
    .B(net75),
    .C(net204),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_1 _0557_ (.A1(\flashBuffer.baseAddress[4] ),
    .A2(net194),
    .B1(_0219_),
    .X(_0015_));
 sky130_fd_sc_hd__nand2_1 _0558_ (.A(net76),
    .B(net204),
    .Y(_0220_));
 sky130_fd_sc_hd__a2bb2o_1 _0559_ (.A1_N(net237),
    .A2_N(_0220_),
    .B1(net195),
    .B2(\flashBuffer.baseAddress[5] ),
    .X(_0016_));
 sky130_fd_sc_hd__and3_4 _0560_ (.A(net228),
    .B(net77),
    .C(net204),
    .X(_0221_));
 sky130_fd_sc_hd__a21o_1 _0561_ (.A1(\flashBuffer.baseAddress[6] ),
    .A2(net194),
    .B1(_0221_),
    .X(_0017_));
 sky130_fd_sc_hd__and3_4 _0562_ (.A(net228),
    .B(net78),
    .C(net205),
    .X(_0222_));
 sky130_fd_sc_hd__a21o_1 _0563_ (.A1(\flashBuffer.baseAddress[7] ),
    .A2(net194),
    .B1(_0222_),
    .X(_0018_));
 sky130_fd_sc_hd__and3_4 _0564_ (.A(net228),
    .B(net79),
    .C(net204),
    .X(_0223_));
 sky130_fd_sc_hd__a21o_1 _0565_ (.A1(\flashBuffer.baseAddress[8] ),
    .A2(net194),
    .B1(_0223_),
    .X(_0019_));
 sky130_fd_sc_hd__and3_4 _0566_ (.A(net229),
    .B(net80),
    .C(net205),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _0567_ (.A1(\flashBuffer.baseAddress[9] ),
    .A2(net196),
    .B1(_0224_),
    .X(_0020_));
 sky130_fd_sc_hd__and3_1 _0568_ (.A(net231),
    .B(net58),
    .C(net207),
    .X(_0225_));
 sky130_fd_sc_hd__a21o_1 _0569_ (.A1(\flashBuffer.baseAddress[10] ),
    .A2(net194),
    .B1(_0225_),
    .X(_0021_));
 sky130_fd_sc_hd__nand2_1 _0570_ (.A(net59),
    .B(net204),
    .Y(_0226_));
 sky130_fd_sc_hd__a2bb2o_1 _0571_ (.A1_N(net237),
    .A2_N(_0226_),
    .B1(net197),
    .B2(\flashBuffer.baseAddress[11] ),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _0572_ (.A(net60),
    .B(net205),
    .Y(_0227_));
 sky130_fd_sc_hd__a2bb2o_1 _0573_ (.A1_N(net237),
    .A2_N(_0227_),
    .B1(net197),
    .B2(\flashBuffer.baseAddress[12] ),
    .X(_0023_));
 sky130_fd_sc_hd__and3_4 _0574_ (.A(net229),
    .B(net61),
    .C(net208),
    .X(_0228_));
 sky130_fd_sc_hd__a21o_1 _0575_ (.A1(\flashBuffer.baseAddress[13] ),
    .A2(net195),
    .B1(_0228_),
    .X(_0024_));
 sky130_fd_sc_hd__nand2_1 _0576_ (.A(net62),
    .B(net206),
    .Y(_0229_));
 sky130_fd_sc_hd__a2bb2o_1 _0577_ (.A1_N(net234),
    .A2_N(_0229_),
    .B1(net196),
    .B2(\flashBuffer.baseAddress[14] ),
    .X(_0025_));
 sky130_fd_sc_hd__nand2_1 _0578_ (.A(net63),
    .B(net206),
    .Y(_0230_));
 sky130_fd_sc_hd__a2bb2o_1 _0579_ (.A1_N(net234),
    .A2_N(_0230_),
    .B1(net198),
    .B2(\flashBuffer.baseAddress[15] ),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _0580_ (.A(net64),
    .B(net206),
    .Y(_0231_));
 sky130_fd_sc_hd__a2bb2o_1 _0581_ (.A1_N(net234),
    .A2_N(_0231_),
    .B1(net198),
    .B2(\flashBuffer.baseAddress[16] ),
    .X(_0027_));
 sky130_fd_sc_hd__and3_1 _0582_ (.A(net232),
    .B(net65),
    .C(net206),
    .X(_0232_));
 sky130_fd_sc_hd__a21o_1 _0583_ (.A1(\flashBuffer.baseAddress[17] ),
    .A2(net198),
    .B1(_0232_),
    .X(_0028_));
 sky130_fd_sc_hd__nand2_1 _0584_ (.A(net66),
    .B(net206),
    .Y(_0233_));
 sky130_fd_sc_hd__a2bb2o_1 _0585_ (.A1_N(net234),
    .A2_N(_0233_),
    .B1(net198),
    .B2(\flashBuffer.baseAddress[18] ),
    .X(_0029_));
 sky130_fd_sc_hd__nand2_1 _0586_ (.A(net67),
    .B(net206),
    .Y(_0234_));
 sky130_fd_sc_hd__a2bb2o_1 _0587_ (.A1_N(net234),
    .A2_N(_0234_),
    .B1(net198),
    .B2(\flashBuffer.baseAddress[19] ),
    .X(_0030_));
 sky130_fd_sc_hd__and3_1 _0588_ (.A(net233),
    .B(net69),
    .C(net207),
    .X(_0235_));
 sky130_fd_sc_hd__a21o_1 _0589_ (.A1(\flashBuffer.baseAddress[20] ),
    .A2(net198),
    .B1(_0235_),
    .X(_0031_));
 sky130_fd_sc_hd__and3_4 _0590_ (.A(net229),
    .B(net70),
    .C(net205),
    .X(_0236_));
 sky130_fd_sc_hd__a21o_1 _0591_ (.A1(\flashBuffer.baseAddress[21] ),
    .A2(net198),
    .B1(_0236_),
    .X(_0032_));
 sky130_fd_sc_hd__and3_4 _0592_ (.A(net229),
    .B(net71),
    .C(net205),
    .X(_0237_));
 sky130_fd_sc_hd__a21o_1 _0593_ (.A1(\flashBuffer.baseAddress[22] ),
    .A2(net197),
    .B1(_0237_),
    .X(_0033_));
 sky130_fd_sc_hd__and3_4 _0594_ (.A(net229),
    .B(net72),
    .C(net205),
    .X(_0238_));
 sky130_fd_sc_hd__a21o_1 _0595_ (.A1(\flashBuffer.baseAddress[23] ),
    .A2(net196),
    .B1(_0238_),
    .X(_0034_));
 sky130_fd_sc_hd__or2_2 _0596_ (.A(\qspiDevice.resetState[1] ),
    .B(\qspiDevice.resetState[0] ),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _0597_ (.A(_0171_),
    .B(\qspiDevice.state[0] ),
    .Y(_0240_));
 sky130_fd_sc_hd__and3_2 _0598_ (.A(_0171_),
    .B(net227),
    .C(_0239_),
    .X(_0241_));
 sky130_fd_sc_hd__a21oi_4 _0599_ (.A1(net87),
    .A2(net206),
    .B1(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _0600_ (.A(net192),
    .Y(_0243_));
 sky130_fd_sc_hd__o21a_2 _0601_ (.A1(net226),
    .A2(net227),
    .B1(\qspiDevice.outputClock ),
    .X(_0244_));
 sky130_fd_sc_hd__o21ai_4 _0602_ (.A1(\qspiDevice.state[1] ),
    .A2(net227),
    .B1(\qspiDevice.outputClock ),
    .Y(_0245_));
 sky130_fd_sc_hd__and2_4 _0603_ (.A(net191),
    .B(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_2 _0604_ (.A(net191),
    .B(_0245_),
    .Y(_0247_));
 sky130_fd_sc_hd__nor2_1 _0605_ (.A(_0241_),
    .B(_0245_),
    .Y(_0248_));
 sky130_fd_sc_hd__or2_2 _0606_ (.A(_0241_),
    .B(_0245_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_2 _0607_ (.A(_0172_),
    .B(\qspiDevice.resetState[0] ),
    .Y(_0250_));
 sky130_fd_sc_hd__or2_1 _0608_ (.A(_0172_),
    .B(\qspiDevice.resetState[0] ),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_2 _0609_ (.A(_0250_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__nor2_1 _0610_ (.A(net191),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__or2_1 _0611_ (.A(net128),
    .B(net218),
    .X(_0254_));
 sky130_fd_sc_hd__o211a_1 _0612_ (.A1(net1),
    .A2(_0245_),
    .B1(_0254_),
    .C1(net191),
    .X(_0255_));
 sky130_fd_sc_hd__a31o_1 _0613_ (.A1(net57),
    .A2(net207),
    .A3(net182),
    .B1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__and2_1 _0614_ (.A(net230),
    .B(_0256_),
    .X(_0035_));
 sky130_fd_sc_hd__or2_1 _0615_ (.A(net129),
    .B(net219),
    .X(_0257_));
 sky130_fd_sc_hd__o211a_1 _0616_ (.A1(net128),
    .A2(_0245_),
    .B1(_0257_),
    .C1(net193),
    .X(_0258_));
 sky130_fd_sc_hd__a31o_1 _0617_ (.A1(net68),
    .A2(net207),
    .A3(net183),
    .B1(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__and2_1 _0618_ (.A(net230),
    .B(_0259_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(net130),
    .A1(net129),
    .S(net219),
    .X(_0260_));
 sky130_fd_sc_hd__and2_1 _0620_ (.A(net207),
    .B(net182),
    .X(_0261_));
 sky130_fd_sc_hd__a32o_1 _0621_ (.A1(net230),
    .A2(net193),
    .A3(_0260_),
    .B1(net182),
    .B2(_0217_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0622_ (.A0(net131),
    .A1(net130),
    .S(net219),
    .X(_0262_));
 sky130_fd_sc_hd__a32o_1 _0623_ (.A1(net230),
    .A2(net193),
    .A3(_0262_),
    .B1(net182),
    .B2(_0218_),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_1 _0624_ (.A1(net132),
    .A2(_0246_),
    .B1(net209),
    .B2(net131),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _0625_ (.A1(_0219_),
    .A2(net182),
    .B1(_0263_),
    .B2(net230),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_1 _0626_ (.A1(net133),
    .A2(_0246_),
    .B1(net209),
    .B2(net132),
    .X(_0264_));
 sky130_fd_sc_hd__a21oi_1 _0627_ (.A1(net76),
    .A2(net178),
    .B1(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor2_1 _0628_ (.A(net236),
    .B(_0265_),
    .Y(_0040_));
 sky130_fd_sc_hd__mux2_1 _0629_ (.A0(net135),
    .A1(net133),
    .S(net219),
    .X(_0266_));
 sky130_fd_sc_hd__a32o_1 _0630_ (.A1(net230),
    .A2(net193),
    .A3(_0266_),
    .B1(net183),
    .B2(_0221_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0631_ (.A0(net136),
    .A1(net135),
    .S(net219),
    .X(_0267_));
 sky130_fd_sc_hd__a32o_1 _0632_ (.A1(net230),
    .A2(net193),
    .A3(_0267_),
    .B1(net183),
    .B2(_0222_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0633_ (.A0(net119),
    .A1(net136),
    .S(net218),
    .X(_0268_));
 sky130_fd_sc_hd__a32o_1 _0634_ (.A1(net230),
    .A2(_0242_),
    .A3(_0268_),
    .B1(net183),
    .B2(_0223_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0635_ (.A0(net120),
    .A1(net119),
    .S(net218),
    .X(_0269_));
 sky130_fd_sc_hd__a32o_1 _0636_ (.A1(net231),
    .A2(net191),
    .A3(_0269_),
    .B1(net182),
    .B2(_0224_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0637_ (.A0(net121),
    .A1(net120),
    .S(net218),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _0638_ (.A1(net58),
    .A2(net178),
    .B1(_0270_),
    .B2(net191),
    .X(_0271_));
 sky130_fd_sc_hd__and2_1 _0639_ (.A(net230),
    .B(_0271_),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _0640_ (.A1(net122),
    .A2(_0246_),
    .B1(net209),
    .B2(net121),
    .X(_0272_));
 sky130_fd_sc_hd__a21oi_1 _0641_ (.A1(net59),
    .A2(net178),
    .B1(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__nor2_1 _0642_ (.A(net236),
    .B(_0273_),
    .Y(_0046_));
 sky130_fd_sc_hd__mux2_1 _0643_ (.A0(net124),
    .A1(net122),
    .S(net218),
    .X(_0274_));
 sky130_fd_sc_hd__a22o_1 _0644_ (.A1(net60),
    .A2(net178),
    .B1(_0274_),
    .B2(net193),
    .X(_0275_));
 sky130_fd_sc_hd__and2_1 _0645_ (.A(net232),
    .B(_0275_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(net125),
    .A1(net124),
    .S(net219),
    .X(_0276_));
 sky130_fd_sc_hd__a32o_1 _0647_ (.A1(net232),
    .A2(net193),
    .A3(_0276_),
    .B1(net182),
    .B2(_0228_),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _0648_ (.A1(net126),
    .A2(_0246_),
    .B1(net209),
    .B2(net125),
    .X(_0277_));
 sky130_fd_sc_hd__a21oi_1 _0649_ (.A1(net62),
    .A2(net178),
    .B1(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__nor2_1 _0650_ (.A(net236),
    .B(_0278_),
    .Y(_0049_));
 sky130_fd_sc_hd__a22o_1 _0651_ (.A1(net127),
    .A2(_0246_),
    .B1(net209),
    .B2(net126),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_1 _0652_ (.A1(net63),
    .A2(net178),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nor2_1 _0653_ (.A(net236),
    .B(_0280_),
    .Y(_0050_));
 sky130_fd_sc_hd__mux2_1 _0654_ (.A0(net142),
    .A1(net127),
    .S(net218),
    .X(_0281_));
 sky130_fd_sc_hd__a22o_1 _0655_ (.A1(net64),
    .A2(net178),
    .B1(_0281_),
    .B2(net192),
    .X(_0282_));
 sky130_fd_sc_hd__and2_1 _0656_ (.A(net232),
    .B(_0282_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0657_ (.A0(net143),
    .A1(net142),
    .S(net218),
    .X(_0283_));
 sky130_fd_sc_hd__a22o_1 _0658_ (.A1(net65),
    .A2(_0261_),
    .B1(_0283_),
    .B2(net192),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _0659_ (.A(net232),
    .B(_0284_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0660_ (.A0(net113),
    .A1(net143),
    .S(net218),
    .X(_0285_));
 sky130_fd_sc_hd__a22o_1 _0661_ (.A1(net66),
    .A2(net178),
    .B1(_0285_),
    .B2(net192),
    .X(_0286_));
 sky130_fd_sc_hd__and2_1 _0662_ (.A(net231),
    .B(_0286_),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_1 _0663_ (.A1(net114),
    .A2(_0246_),
    .B1(net209),
    .B2(net113),
    .X(_0287_));
 sky130_fd_sc_hd__a21oi_1 _0664_ (.A1(net67),
    .A2(net178),
    .B1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nor2_1 _0665_ (.A(net236),
    .B(_0288_),
    .Y(_0054_));
 sky130_fd_sc_hd__a22o_1 _0666_ (.A1(net115),
    .A2(_0246_),
    .B1(net209),
    .B2(net114),
    .X(_0289_));
 sky130_fd_sc_hd__a21oi_1 _0667_ (.A1(net69),
    .A2(net178),
    .B1(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__nor2_1 _0668_ (.A(net236),
    .B(_0290_),
    .Y(_0055_));
 sky130_fd_sc_hd__mux2_1 _0669_ (.A0(net116),
    .A1(net115),
    .S(net218),
    .X(_0291_));
 sky130_fd_sc_hd__a32o_1 _0670_ (.A1(net232),
    .A2(net193),
    .A3(_0291_),
    .B1(net183),
    .B2(_0236_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0671_ (.A0(net117),
    .A1(net116),
    .S(net218),
    .X(_0292_));
 sky130_fd_sc_hd__a32o_1 _0672_ (.A1(net231),
    .A2(net191),
    .A3(_0292_),
    .B1(net182),
    .B2(_0237_),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _0673_ (.A(net118),
    .B(net191),
    .X(_0293_));
 sky130_fd_sc_hd__o22a_1 _0674_ (.A1(net117),
    .A2(_0245_),
    .B1(net209),
    .B2(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_1 _0675_ (.A1(_0238_),
    .A2(net182),
    .B1(_0294_),
    .B2(net231),
    .X(_0058_));
 sky130_fd_sc_hd__o31a_1 _0676_ (.A1(net207),
    .A2(net191),
    .A3(_0252_),
    .B1(_0249_),
    .X(_0295_));
 sky130_fd_sc_hd__o221a_1 _0677_ (.A1(net112),
    .A2(_0247_),
    .B1(_0293_),
    .B2(_0295_),
    .C1(net231),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _0678_ (.A(net112),
    .B(net191),
    .X(_0296_));
 sky130_fd_sc_hd__o221a_1 _0679_ (.A1(net123),
    .A2(_0247_),
    .B1(_0295_),
    .B2(_0296_),
    .C1(net231),
    .X(_0060_));
 sky130_fd_sc_hd__nor2_2 _0680_ (.A(net192),
    .B(_0250_),
    .Y(_0297_));
 sky130_fd_sc_hd__a221o_1 _0681_ (.A1(net134),
    .A2(_0246_),
    .B1(net209),
    .B2(net123),
    .C1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__and2_1 _0682_ (.A(net231),
    .B(_0298_),
    .X(_0061_));
 sky130_fd_sc_hd__nor2_2 _0683_ (.A(net236),
    .B(net182),
    .Y(_0299_));
 sky130_fd_sc_hd__o221a_1 _0684_ (.A1(net137),
    .A2(_0247_),
    .B1(_0249_),
    .B2(net134),
    .C1(_0299_),
    .X(_0062_));
 sky130_fd_sc_hd__a221o_1 _0685_ (.A1(net138),
    .A2(_0246_),
    .B1(_0248_),
    .B2(net137),
    .C1(_0297_),
    .X(_0300_));
 sky130_fd_sc_hd__and2_1 _0686_ (.A(net230),
    .B(_0300_),
    .X(_0063_));
 sky130_fd_sc_hd__o221a_1 _0687_ (.A1(net139),
    .A2(_0247_),
    .B1(_0249_),
    .B2(net138),
    .C1(_0299_),
    .X(_0064_));
 sky130_fd_sc_hd__a221o_1 _0688_ (.A1(net140),
    .A2(_0246_),
    .B1(net209),
    .B2(net139),
    .C1(_0297_),
    .X(_0301_));
 sky130_fd_sc_hd__and2_1 _0689_ (.A(net231),
    .B(_0301_),
    .X(_0065_));
 sky130_fd_sc_hd__o221a_1 _0690_ (.A1(net141),
    .A2(_0247_),
    .B1(_0249_),
    .B2(net140),
    .C1(_0299_),
    .X(_0066_));
 sky130_fd_sc_hd__nor2_1 _0691_ (.A(\qspiDevice.outputClock ),
    .B(net87),
    .Y(_0302_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(\qspiDevice.register.outputBit ),
    .A1(net141),
    .S(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__o21a_1 _0693_ (.A1(_0243_),
    .A2(_0303_),
    .B1(_0299_),
    .X(_0067_));
 sky130_fd_sc_hd__nand2_2 _0694_ (.A(net226),
    .B(net227),
    .Y(_0304_));
 sky130_fd_sc_hd__a21o_1 _0695_ (.A1(\qspiDevice.resetState[0] ),
    .A2(_0304_),
    .B1(net234),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(_0250_),
    .A1(_0172_),
    .S(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__nor2_1 _0697_ (.A(net235),
    .B(_0305_),
    .Y(_0069_));
 sky130_fd_sc_hd__o211a_1 _0698_ (.A1(net206),
    .A2(_0239_),
    .B1(\flashBuffer.configuration ),
    .C1(net87),
    .X(_0306_));
 sky130_fd_sc_hd__and3_1 _0699_ (.A(net226),
    .B(net227),
    .C(\flashBuffer.qspi_requestData ),
    .X(_0307_));
 sky130_fd_sc_hd__or3_1 _0700_ (.A(_0171_),
    .B(\qspiDevice.state[0] ),
    .C(net206),
    .X(_0308_));
 sky130_fd_sc_hd__nand3_2 _0701_ (.A(\qspiDevice.bitCounter[2] ),
    .B(\qspiDevice.bitCounter[1] ),
    .C(\qspiDevice.bitCounter[0] ),
    .Y(_0309_));
 sky130_fd_sc_hd__a21oi_1 _0702_ (.A1(_0168_),
    .A2(_0239_),
    .B1(\qspiDevice.bitCounter[3] ),
    .Y(_0310_));
 sky130_fd_sc_hd__a211oi_2 _0703_ (.A1(_0168_),
    .A2(\qspiDevice.bitCounter[3] ),
    .B1(_0309_),
    .C1(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__and2b_1 _0704_ (.A_N(\qspiDevice.outputClock ),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__and2b_1 _0705_ (.A_N(_0308_),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__o31a_1 _0706_ (.A1(_0306_),
    .A2(_0307_),
    .A3(_0313_),
    .B1(net233),
    .X(_0070_));
 sky130_fd_sc_hd__a21oi_1 _0707_ (.A1(_0240_),
    .A2(_0308_),
    .B1(net234),
    .Y(_0071_));
 sky130_fd_sc_hd__and2_1 _0708_ (.A(net226),
    .B(_0312_),
    .X(_0314_));
 sky130_fd_sc_hd__a211o_1 _0709_ (.A1(\qspiDevice.settingAddress ),
    .A2(_0314_),
    .B1(net234),
    .C1(net227),
    .X(_0315_));
 sky130_fd_sc_hd__o21ba_1 _0710_ (.A1(\flashBuffer.qspi_readDataValid ),
    .A2(_0314_),
    .B1_N(_0315_),
    .X(_0072_));
 sky130_fd_sc_hd__nor2_1 _0711_ (.A(net237),
    .B(net111),
    .Y(_0073_));
 sky130_fd_sc_hd__and3b_1 _0712_ (.A_N(_0306_),
    .B(\qspiDevice.settingAddress ),
    .C(_0304_),
    .X(_0316_));
 sky130_fd_sc_hd__and3_1 _0713_ (.A(\flashBuffer.configuration ),
    .B(net87),
    .C(net205),
    .X(_0317_));
 sky130_fd_sc_hd__o21a_1 _0714_ (.A1(_0316_),
    .A2(_0317_),
    .B1(net233),
    .X(_0074_));
 sky130_fd_sc_hd__nor2_1 _0715_ (.A(\qspiDevice.outputClock ),
    .B(net227),
    .Y(_0318_));
 sky130_fd_sc_hd__or3_2 _0716_ (.A(\qspiDevice.outputClock ),
    .B(net227),
    .C(_0311_),
    .X(_0319_));
 sky130_fd_sc_hd__nand2_1 _0717_ (.A(net226),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__o211a_1 _0718_ (.A1(net226),
    .A2(net227),
    .B1(net232),
    .C1(_0320_),
    .X(_0075_));
 sky130_fd_sc_hd__nor2_2 _0719_ (.A(_0171_),
    .B(net235),
    .Y(_0321_));
 sky130_fd_sc_hd__o21a_1 _0720_ (.A1(\qspiDevice.bitCounter[0] ),
    .A2(_0318_),
    .B1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__o21a_1 _0721_ (.A1(_0169_),
    .A2(_0319_),
    .B1(_0322_),
    .X(_0076_));
 sky130_fd_sc_hd__a21o_1 _0722_ (.A1(\qspiDevice.bitCounter[0] ),
    .A2(_0320_),
    .B1(\qspiDevice.bitCounter[1] ),
    .X(_0323_));
 sky130_fd_sc_hd__and4b_1 _0723_ (.A_N(_0311_),
    .B(_0318_),
    .C(\qspiDevice.bitCounter[1] ),
    .D(\qspiDevice.bitCounter[0] ),
    .X(_0324_));
 sky130_fd_sc_hd__and3b_1 _0724_ (.A_N(_0324_),
    .B(_0321_),
    .C(_0323_),
    .X(_0077_));
 sky130_fd_sc_hd__o221a_1 _0725_ (.A1(_0309_),
    .A2(_0319_),
    .B1(_0324_),
    .B2(\qspiDevice.bitCounter[2] ),
    .C1(_0321_),
    .X(_0078_));
 sky130_fd_sc_hd__a41o_1 _0726_ (.A1(\qspiDevice.bitCounter[2] ),
    .A2(\qspiDevice.bitCounter[1] ),
    .A3(\qspiDevice.bitCounter[0] ),
    .A4(_0320_),
    .B1(\qspiDevice.bitCounter[3] ),
    .X(_0325_));
 sky130_fd_sc_hd__nand3_1 _0727_ (.A(\qspiDevice.bitCounter[3] ),
    .B(\qspiDevice.bitCounter[2] ),
    .C(_0324_),
    .Y(_0326_));
 sky130_fd_sc_hd__and4_1 _0728_ (.A(net226),
    .B(net232),
    .C(_0325_),
    .D(_0326_),
    .X(_0079_));
 sky130_fd_sc_hd__a21boi_1 _0729_ (.A1(_0168_),
    .A2(_0326_),
    .B1_N(_0321_),
    .Y(_0080_));
 sky130_fd_sc_hd__and3_1 _0730_ (.A(net90),
    .B(\flashBuffer.qspi_readDataValid ),
    .C(\flashBuffer.qspi_requestData ),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_1 _0731_ (.A(net90),
    .B(_0184_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_1 _0732_ (.A(_0327_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a21o_1 _0733_ (.A1(net195),
    .A2(_0329_),
    .B1(_0217_),
    .X(_0081_));
 sky130_fd_sc_hd__nor2_1 _0734_ (.A(net91),
    .B(_0327_),
    .Y(_0330_));
 sky130_fd_sc_hd__and4_2 _0735_ (.A(net91),
    .B(net90),
    .C(\flashBuffer.qspi_readDataValid ),
    .D(\flashBuffer.qspi_requestData ),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_1 _0736_ (.A(_0330_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a21o_1 _0737_ (.A1(net195),
    .A2(_0332_),
    .B1(_0218_),
    .X(_0082_));
 sky130_fd_sc_hd__nand2_1 _0738_ (.A(net92),
    .B(_0331_),
    .Y(_0333_));
 sky130_fd_sc_hd__or2_1 _0739_ (.A(net92),
    .B(_0331_),
    .X(_0334_));
 sky130_fd_sc_hd__a31o_1 _0740_ (.A1(net195),
    .A2(_0333_),
    .A3(_0334_),
    .B1(_0219_),
    .X(_0083_));
 sky130_fd_sc_hd__and3_1 _0741_ (.A(net93),
    .B(net92),
    .C(_0331_),
    .X(_0335_));
 sky130_fd_sc_hd__a21oi_1 _0742_ (.A1(net92),
    .A2(_0331_),
    .B1(net93),
    .Y(_0336_));
 sky130_fd_sc_hd__o31a_1 _0743_ (.A1(net204),
    .A2(_0335_),
    .A3(_0336_),
    .B1(_0220_),
    .X(_0337_));
 sky130_fd_sc_hd__nor2_1 _0744_ (.A(net237),
    .B(_0337_),
    .Y(_0084_));
 sky130_fd_sc_hd__and4_4 _0745_ (.A(net94),
    .B(net93),
    .C(net92),
    .D(_0331_),
    .X(_0338_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(net94),
    .B(_0335_),
    .X(_0340_));
 sky130_fd_sc_hd__a31o_1 _0748_ (.A1(net195),
    .A2(_0339_),
    .A3(_0340_),
    .B1(_0221_),
    .X(_0085_));
 sky130_fd_sc_hd__xor2_1 _0749_ (.A(net95),
    .B(_0338_),
    .X(_0341_));
 sky130_fd_sc_hd__a21o_1 _0750_ (.A1(net194),
    .A2(_0341_),
    .B1(_0222_),
    .X(_0086_));
 sky130_fd_sc_hd__and3_1 _0751_ (.A(net96),
    .B(net95),
    .C(_0338_),
    .X(_0342_));
 sky130_fd_sc_hd__a21oi_1 _0752_ (.A1(net95),
    .A2(_0338_),
    .B1(net96),
    .Y(_0343_));
 sky130_fd_sc_hd__nor2_1 _0753_ (.A(_0342_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__a21o_1 _0754_ (.A1(net194),
    .A2(_0344_),
    .B1(_0223_),
    .X(_0087_));
 sky130_fd_sc_hd__or2_1 _0755_ (.A(net97),
    .B(_0342_),
    .X(_0345_));
 sky130_fd_sc_hd__and4_4 _0756_ (.A(net97),
    .B(net96),
    .C(net95),
    .D(_0338_),
    .X(_0346_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__a31o_1 _0758_ (.A1(net194),
    .A2(_0345_),
    .A3(_0347_),
    .B1(_0224_),
    .X(_0088_));
 sky130_fd_sc_hd__nand2_1 _0759_ (.A(net98),
    .B(_0346_),
    .Y(_0348_));
 sky130_fd_sc_hd__o211a_1 _0760_ (.A1(net98),
    .A2(_0346_),
    .B1(_0348_),
    .C1(net194),
    .X(_0349_));
 sky130_fd_sc_hd__or2_1 _0761_ (.A(_0225_),
    .B(_0349_),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _0762_ (.A(\flashBuffer.cachedAddress[11] ),
    .B(net98),
    .X(_0350_));
 sky130_fd_sc_hd__and2_2 _0763_ (.A(_0346_),
    .B(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__a211o_1 _0764_ (.A1(_0167_),
    .A2(_0348_),
    .B1(_0351_),
    .C1(net207),
    .X(_0352_));
 sky130_fd_sc_hd__a21oi_1 _0765_ (.A1(_0226_),
    .A2(_0352_),
    .B1(net236),
    .Y(_0090_));
 sky130_fd_sc_hd__o21ai_1 _0766_ (.A1(\flashBuffer.cachedAddress[12] ),
    .A2(_0351_),
    .B1(net194),
    .Y(_0353_));
 sky130_fd_sc_hd__a21o_1 _0767_ (.A1(\flashBuffer.cachedAddress[12] ),
    .A2(_0351_),
    .B1(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__o21ai_1 _0768_ (.A1(net234),
    .A2(_0227_),
    .B1(_0354_),
    .Y(_0091_));
 sky130_fd_sc_hd__and4_4 _0769_ (.A(\flashBuffer.cachedAddress[13] ),
    .B(\flashBuffer.cachedAddress[12] ),
    .C(_0346_),
    .D(_0350_),
    .X(_0355_));
 sky130_fd_sc_hd__a21oi_1 _0770_ (.A1(\flashBuffer.cachedAddress[12] ),
    .A2(_0351_),
    .B1(\flashBuffer.cachedAddress[13] ),
    .Y(_0356_));
 sky130_fd_sc_hd__nor3_1 _0771_ (.A(_0198_),
    .B(_0355_),
    .C(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__or2_1 _0772_ (.A(_0228_),
    .B(_0357_),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_1 _0773_ (.A(\flashBuffer.cachedAddress[14] ),
    .B(_0355_),
    .Y(_0358_));
 sky130_fd_sc_hd__a211o_1 _0774_ (.A1(\flashBuffer.cachedAddress[14] ),
    .A2(_0355_),
    .B1(_0358_),
    .C1(_0198_),
    .X(_0359_));
 sky130_fd_sc_hd__o21ai_1 _0775_ (.A1(net234),
    .A2(_0229_),
    .B1(_0359_),
    .Y(_0093_));
 sky130_fd_sc_hd__a21oi_1 _0776_ (.A1(\flashBuffer.cachedAddress[14] ),
    .A2(_0355_),
    .B1(\flashBuffer.cachedAddress[15] ),
    .Y(_0360_));
 sky130_fd_sc_hd__and3_1 _0777_ (.A(\flashBuffer.cachedAddress[15] ),
    .B(\flashBuffer.cachedAddress[14] ),
    .C(_0355_),
    .X(_0361_));
 sky130_fd_sc_hd__o31a_1 _0778_ (.A1(net207),
    .A2(_0360_),
    .A3(_0361_),
    .B1(_0230_),
    .X(_0362_));
 sky130_fd_sc_hd__nor2_1 _0779_ (.A(net235),
    .B(_0362_),
    .Y(_0094_));
 sky130_fd_sc_hd__and4_4 _0780_ (.A(\flashBuffer.cachedAddress[16] ),
    .B(\flashBuffer.cachedAddress[15] ),
    .C(\flashBuffer.cachedAddress[14] ),
    .D(_0355_),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_1 _0781_ (.A(\flashBuffer.cachedAddress[16] ),
    .B(_0361_),
    .Y(_0364_));
 sky130_fd_sc_hd__o31a_1 _0782_ (.A1(net207),
    .A2(_0363_),
    .A3(_0364_),
    .B1(_0231_),
    .X(_0365_));
 sky130_fd_sc_hd__nor2_1 _0783_ (.A(net235),
    .B(_0365_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_1 _0784_ (.A(\flashBuffer.cachedAddress[17] ),
    .B(_0363_),
    .Y(_0366_));
 sky130_fd_sc_hd__o211a_1 _0785_ (.A1(\flashBuffer.cachedAddress[17] ),
    .A2(_0363_),
    .B1(_0366_),
    .C1(net198),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _0786_ (.A(_0232_),
    .B(_0367_),
    .X(_0096_));
 sky130_fd_sc_hd__and3_1 _0787_ (.A(\flashBuffer.cachedAddress[18] ),
    .B(\flashBuffer.cachedAddress[17] ),
    .C(_0363_),
    .X(_0368_));
 sky130_fd_sc_hd__a21oi_1 _0788_ (.A1(\flashBuffer.cachedAddress[17] ),
    .A2(_0363_),
    .B1(\flashBuffer.cachedAddress[18] ),
    .Y(_0369_));
 sky130_fd_sc_hd__o31a_1 _0789_ (.A1(net208),
    .A2(_0368_),
    .A3(_0369_),
    .B1(_0233_),
    .X(_0370_));
 sky130_fd_sc_hd__nor2_1 _0790_ (.A(net235),
    .B(_0370_),
    .Y(_0097_));
 sky130_fd_sc_hd__nor2_1 _0791_ (.A(\flashBuffer.cachedAddress[19] ),
    .B(_0368_),
    .Y(_0371_));
 sky130_fd_sc_hd__and4_4 _0792_ (.A(\flashBuffer.cachedAddress[19] ),
    .B(\flashBuffer.cachedAddress[18] ),
    .C(\flashBuffer.cachedAddress[17] ),
    .D(_0363_),
    .X(_0372_));
 sky130_fd_sc_hd__o31a_1 _0793_ (.A1(net206),
    .A2(_0371_),
    .A3(_0372_),
    .B1(_0234_),
    .X(_0373_));
 sky130_fd_sc_hd__nor2_1 _0794_ (.A(net235),
    .B(_0373_),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_1 _0795_ (.A(\flashBuffer.cachedAddress[20] ),
    .B(_0372_),
    .Y(_0374_));
 sky130_fd_sc_hd__o211a_1 _0796_ (.A1(\flashBuffer.cachedAddress[20] ),
    .A2(_0372_),
    .B1(_0374_),
    .C1(net198),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _0797_ (.A(_0235_),
    .B(_0375_),
    .X(_0099_));
 sky130_fd_sc_hd__a21o_1 _0798_ (.A1(\flashBuffer.cachedAddress[20] ),
    .A2(_0372_),
    .B1(\flashBuffer.cachedAddress[21] ),
    .X(_0376_));
 sky130_fd_sc_hd__nand3_2 _0799_ (.A(\flashBuffer.cachedAddress[21] ),
    .B(\flashBuffer.cachedAddress[20] ),
    .C(_0372_),
    .Y(_0377_));
 sky130_fd_sc_hd__a31o_1 _0800_ (.A1(_0197_),
    .A2(_0376_),
    .A3(_0377_),
    .B1(_0236_),
    .X(_0100_));
 sky130_fd_sc_hd__and4_1 _0801_ (.A(\flashBuffer.cachedAddress[22] ),
    .B(\flashBuffer.cachedAddress[21] ),
    .C(\flashBuffer.cachedAddress[20] ),
    .D(_0372_),
    .X(_0378_));
 sky130_fd_sc_hd__xnor2_1 _0802_ (.A(\flashBuffer.cachedAddress[22] ),
    .B(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__a21o_1 _0803_ (.A1(net198),
    .A2(_0379_),
    .B1(_0237_),
    .X(_0101_));
 sky130_fd_sc_hd__xor2_1 _0804_ (.A(\flashBuffer.cachedAddress[23] ),
    .B(_0378_),
    .X(_0380_));
 sky130_fd_sc_hd__a21o_1 _0805_ (.A1(_0197_),
    .A2(_0380_),
    .B1(_0238_),
    .X(_0102_));
 sky130_fd_sc_hd__nor2_1 _0806_ (.A(net99),
    .B(_0190_),
    .Y(_0381_));
 sky130_fd_sc_hd__nor3b_1 _0807_ (.A(net100),
    .B(_0195_),
    .C_N(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__and4b_1 _0808_ (.A_N(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .C(net225),
    .D(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(\flashBuffer.configuration ),
    .A1(net57),
    .S(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__and2_1 _0810_ (.A(net228),
    .B(_0384_),
    .X(_0103_));
 sky130_fd_sc_hd__nor4b_4 _0811_ (.A(_0175_),
    .B(_0179_),
    .C(_0195_),
    .D_N(_0381_),
    .Y(_0385_));
 sky130_fd_sc_hd__and2b_1 _0812_ (.A_N(_0385_),
    .B(\flashBuffer.flashCacheReadReady ),
    .X(_0386_));
 sky130_fd_sc_hd__nor3_4 _0813_ (.A(_0179_),
    .B(_0191_),
    .C(_0195_),
    .Y(_0387_));
 sky130_fd_sc_hd__or3_1 _0814_ (.A(_0179_),
    .B(_0191_),
    .C(_0195_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_2 _0815_ (.A(\flashBuffer.flashCacheReadReady ),
    .B(net111),
    .X(_0389_));
 sky130_fd_sc_hd__nand2_2 _0816_ (.A(_0166_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__and3_1 _0817_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(_0166_),
    .C(_0382_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_1 _0818_ (.A(net185),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__and3_4 _0819_ (.A(net188),
    .B(net201),
    .C(net181),
    .X(_0393_));
 sky130_fd_sc_hd__and3_1 _0820_ (.A(\flashBuffer.configuration ),
    .B(net225),
    .C(net220),
    .X(_0394_));
 sky130_fd_sc_hd__xnor2_1 _0821_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .Y(_0395_));
 sky130_fd_sc_hd__or2_1 _0822_ (.A(net237),
    .B(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__and3_1 _0823_ (.A(net225),
    .B(net220),
    .C(net203),
    .X(_0397_));
 sky130_fd_sc_hd__a32o_1 _0824_ (.A1(net2),
    .A2(net188),
    .A3(net201),
    .B1(_0397_),
    .B2(\flashBuffer.baseAddress[0] ),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(_0398_),
    .A1(_0394_),
    .S(_0391_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _0826_ (.A0(_0399_),
    .A1(net145),
    .S(net185),
    .X(_0400_));
 sky130_fd_sc_hd__or2_1 _0827_ (.A(net213),
    .B(_0400_),
    .X(_0104_));
 sky130_fd_sc_hd__a221o_1 _0828_ (.A1(net156),
    .A2(net185),
    .B1(_0397_),
    .B2(\flashBuffer.baseAddress[1] ),
    .C1(net213),
    .X(_0401_));
 sky130_fd_sc_hd__a21o_1 _0829_ (.A1(net13),
    .A2(_0393_),
    .B1(_0401_),
    .X(_0105_));
 sky130_fd_sc_hd__and3_4 _0830_ (.A(net225),
    .B(net224),
    .C(_0385_),
    .X(_0402_));
 sky130_fd_sc_hd__a221o_1 _0831_ (.A1(net24),
    .A2(net188),
    .B1(_0402_),
    .B2(net90),
    .C1(net203),
    .X(_0403_));
 sky130_fd_sc_hd__a31o_1 _0832_ (.A1(\flashBuffer.baseAddress[2] ),
    .A2(net225),
    .A3(net220),
    .B1(net201),
    .X(_0404_));
 sky130_fd_sc_hd__a31o_1 _0833_ (.A1(net181),
    .A2(_0403_),
    .A3(_0404_),
    .B1(net213),
    .X(_0405_));
 sky130_fd_sc_hd__a21o_1 _0834_ (.A1(net167),
    .A2(net185),
    .B1(_0405_),
    .X(_0106_));
 sky130_fd_sc_hd__a221o_1 _0835_ (.A1(net27),
    .A2(net188),
    .B1(_0402_),
    .B2(net91),
    .C1(net203),
    .X(_0406_));
 sky130_fd_sc_hd__a31o_1 _0836_ (.A1(\flashBuffer.baseAddress[3] ),
    .A2(net225),
    .A3(net224),
    .B1(net200),
    .X(_0407_));
 sky130_fd_sc_hd__a31o_1 _0837_ (.A1(net181),
    .A2(_0406_),
    .A3(_0407_),
    .B1(net213),
    .X(_0408_));
 sky130_fd_sc_hd__a21o_1 _0838_ (.A1(net170),
    .A2(net185),
    .B1(_0408_),
    .X(_0107_));
 sky130_fd_sc_hd__a221o_1 _0839_ (.A1(net28),
    .A2(net188),
    .B1(_0402_),
    .B2(net92),
    .C1(net203),
    .X(_0409_));
 sky130_fd_sc_hd__a31o_1 _0840_ (.A1(\flashBuffer.baseAddress[4] ),
    .A2(net225),
    .A3(net224),
    .B1(net200),
    .X(_0410_));
 sky130_fd_sc_hd__a31o_1 _0841_ (.A1(net181),
    .A2(_0409_),
    .A3(_0410_),
    .B1(net216),
    .X(_0411_));
 sky130_fd_sc_hd__a21o_1 _0842_ (.A1(net171),
    .A2(net185),
    .B1(_0411_),
    .X(_0108_));
 sky130_fd_sc_hd__a221o_1 _0843_ (.A1(net29),
    .A2(net188),
    .B1(_0402_),
    .B2(net93),
    .C1(net203),
    .X(_0412_));
 sky130_fd_sc_hd__a31o_1 _0844_ (.A1(\flashBuffer.baseAddress[5] ),
    .A2(net225),
    .A3(net224),
    .B1(net201),
    .X(_0413_));
 sky130_fd_sc_hd__a31o_1 _0845_ (.A1(net181),
    .A2(_0412_),
    .A3(_0413_),
    .B1(net216),
    .X(_0414_));
 sky130_fd_sc_hd__a21o_1 _0846_ (.A1(net172),
    .A2(net185),
    .B1(_0414_),
    .X(_0109_));
 sky130_fd_sc_hd__a221o_1 _0847_ (.A1(net30),
    .A2(net188),
    .B1(_0402_),
    .B2(net94),
    .C1(net203),
    .X(_0415_));
 sky130_fd_sc_hd__a31o_1 _0848_ (.A1(\flashBuffer.baseAddress[6] ),
    .A2(net225),
    .A3(net224),
    .B1(net200),
    .X(_0416_));
 sky130_fd_sc_hd__a31o_1 _0849_ (.A1(net180),
    .A2(_0415_),
    .A3(_0416_),
    .B1(net216),
    .X(_0417_));
 sky130_fd_sc_hd__a21o_1 _0850_ (.A1(net173),
    .A2(net187),
    .B1(_0417_),
    .X(_0110_));
 sky130_fd_sc_hd__a221o_1 _0851_ (.A1(net31),
    .A2(net188),
    .B1(_0402_),
    .B2(net95),
    .C1(net203),
    .X(_0418_));
 sky130_fd_sc_hd__a31o_1 _0852_ (.A1(\flashBuffer.baseAddress[7] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[0] ),
    .A3(net224),
    .B1(net200),
    .X(_0419_));
 sky130_fd_sc_hd__a31o_1 _0853_ (.A1(net180),
    .A2(_0418_),
    .A3(_0419_),
    .B1(net216),
    .X(_0420_));
 sky130_fd_sc_hd__a21o_1 _0854_ (.A1(net174),
    .A2(net185),
    .B1(_0420_),
    .X(_0111_));
 sky130_fd_sc_hd__and3_4 _0855_ (.A(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .B(net224),
    .C(_0385_),
    .X(_0421_));
 sky130_fd_sc_hd__a221o_1 _0856_ (.A1(net32),
    .A2(net188),
    .B1(_0421_),
    .B2(net96),
    .C1(net203),
    .X(_0422_));
 sky130_fd_sc_hd__a31o_1 _0857_ (.A1(\flashBuffer.baseAddress[8] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net222),
    .B1(net200),
    .X(_0423_));
 sky130_fd_sc_hd__a31o_1 _0858_ (.A1(net180),
    .A2(_0422_),
    .A3(_0423_),
    .B1(net214),
    .X(_0424_));
 sky130_fd_sc_hd__a21o_1 _0859_ (.A1(net175),
    .A2(net187),
    .B1(_0424_),
    .X(_0112_));
 sky130_fd_sc_hd__a221o_2 _0860_ (.A1(net33),
    .A2(net188),
    .B1(_0421_),
    .B2(net97),
    .C1(net203),
    .X(_0425_));
 sky130_fd_sc_hd__a31o_1 _0861_ (.A1(\flashBuffer.baseAddress[9] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net223),
    .B1(net201),
    .X(_0426_));
 sky130_fd_sc_hd__a31o_1 _0862_ (.A1(net181),
    .A2(_0425_),
    .A3(_0426_),
    .B1(net215),
    .X(_0427_));
 sky130_fd_sc_hd__a21o_1 _0863_ (.A1(net176),
    .A2(net186),
    .B1(_0427_),
    .X(_0113_));
 sky130_fd_sc_hd__a221o_1 _0864_ (.A1(net3),
    .A2(net189),
    .B1(_0421_),
    .B2(net98),
    .C1(net202),
    .X(_0428_));
 sky130_fd_sc_hd__a31o_1 _0865_ (.A1(\flashBuffer.baseAddress[10] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net224),
    .B1(net200),
    .X(_0429_));
 sky130_fd_sc_hd__a31o_1 _0866_ (.A1(net180),
    .A2(_0428_),
    .A3(_0429_),
    .B1(net216),
    .X(_0430_));
 sky130_fd_sc_hd__a21o_1 _0867_ (.A1(net146),
    .A2(net187),
    .B1(_0430_),
    .X(_0114_));
 sky130_fd_sc_hd__a221o_1 _0868_ (.A1(net4),
    .A2(net189),
    .B1(_0421_),
    .B2(\flashBuffer.cachedAddress[11] ),
    .C1(net202),
    .X(_0431_));
 sky130_fd_sc_hd__a31o_1 _0869_ (.A1(\flashBuffer.baseAddress[11] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net222),
    .B1(net200),
    .X(_0432_));
 sky130_fd_sc_hd__a31o_1 _0870_ (.A1(net180),
    .A2(_0431_),
    .A3(_0432_),
    .B1(net214),
    .X(_0433_));
 sky130_fd_sc_hd__a21o_1 _0871_ (.A1(net147),
    .A2(net186),
    .B1(_0433_),
    .X(_0115_));
 sky130_fd_sc_hd__a221o_1 _0872_ (.A1(net5),
    .A2(net190),
    .B1(_0421_),
    .B2(\flashBuffer.cachedAddress[12] ),
    .C1(net203),
    .X(_0434_));
 sky130_fd_sc_hd__a31o_1 _0873_ (.A1(\flashBuffer.baseAddress[12] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net223),
    .B1(net199),
    .X(_0435_));
 sky130_fd_sc_hd__a31o_1 _0874_ (.A1(net179),
    .A2(_0434_),
    .A3(_0435_),
    .B1(net215),
    .X(_0436_));
 sky130_fd_sc_hd__a21o_1 _0875_ (.A1(net148),
    .A2(net187),
    .B1(_0436_),
    .X(_0116_));
 sky130_fd_sc_hd__a221o_2 _0876_ (.A1(net6),
    .A2(net189),
    .B1(_0421_),
    .B2(\flashBuffer.cachedAddress[13] ),
    .C1(net202),
    .X(_0437_));
 sky130_fd_sc_hd__a31o_1 _0877_ (.A1(\flashBuffer.baseAddress[13] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net221),
    .B1(net201),
    .X(_0438_));
 sky130_fd_sc_hd__a31o_1 _0878_ (.A1(net181),
    .A2(_0437_),
    .A3(_0438_),
    .B1(net213),
    .X(_0439_));
 sky130_fd_sc_hd__a21o_1 _0879_ (.A1(net149),
    .A2(net184),
    .B1(_0439_),
    .X(_0117_));
 sky130_fd_sc_hd__a221o_1 _0880_ (.A1(net7),
    .A2(net189),
    .B1(_0421_),
    .B2(\flashBuffer.cachedAddress[14] ),
    .C1(net202),
    .X(_0440_));
 sky130_fd_sc_hd__a31o_1 _0881_ (.A1(\flashBuffer.baseAddress[14] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net222),
    .B1(net200),
    .X(_0441_));
 sky130_fd_sc_hd__a31o_1 _0882_ (.A1(net179),
    .A2(_0440_),
    .A3(_0441_),
    .B1(net214),
    .X(_0442_));
 sky130_fd_sc_hd__a21o_1 _0883_ (.A1(net150),
    .A2(net186),
    .B1(_0442_),
    .X(_0118_));
 sky130_fd_sc_hd__a221o_1 _0884_ (.A1(net8),
    .A2(net189),
    .B1(_0421_),
    .B2(\flashBuffer.cachedAddress[15] ),
    .C1(net202),
    .X(_0443_));
 sky130_fd_sc_hd__a31o_1 _0885_ (.A1(\flashBuffer.baseAddress[15] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A3(net222),
    .B1(net199),
    .X(_0444_));
 sky130_fd_sc_hd__a31o_1 _0886_ (.A1(net179),
    .A2(_0443_),
    .A3(_0444_),
    .B1(net214),
    .X(_0445_));
 sky130_fd_sc_hd__a21o_1 _0887_ (.A1(net151),
    .A2(net186),
    .B1(_0445_),
    .X(_0119_));
 sky130_fd_sc_hd__and3_4 _0888_ (.A(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .B(net222),
    .C(_0385_),
    .X(_0446_));
 sky130_fd_sc_hd__a221o_1 _0889_ (.A1(net9),
    .A2(net189),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[16] ),
    .C1(net202),
    .X(_0447_));
 sky130_fd_sc_hd__a31o_1 _0890_ (.A1(\flashBuffer.baseAddress[16] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net222),
    .B1(net199),
    .X(_0448_));
 sky130_fd_sc_hd__a31o_1 _0891_ (.A1(net179),
    .A2(_0447_),
    .A3(_0448_),
    .B1(net214),
    .X(_0449_));
 sky130_fd_sc_hd__a21o_1 _0892_ (.A1(net152),
    .A2(net184),
    .B1(_0449_),
    .X(_0120_));
 sky130_fd_sc_hd__a221o_1 _0893_ (.A1(net10),
    .A2(net189),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[17] ),
    .C1(net202),
    .X(_0450_));
 sky130_fd_sc_hd__a31o_1 _0894_ (.A1(\flashBuffer.baseAddress[17] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net222),
    .B1(net199),
    .X(_0451_));
 sky130_fd_sc_hd__a31o_1 _0895_ (.A1(net179),
    .A2(_0450_),
    .A3(_0451_),
    .B1(net214),
    .X(_0452_));
 sky130_fd_sc_hd__a21o_1 _0896_ (.A1(net153),
    .A2(net184),
    .B1(_0452_),
    .X(_0121_));
 sky130_fd_sc_hd__a221o_2 _0897_ (.A1(net11),
    .A2(net189),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[18] ),
    .C1(net202),
    .X(_0453_));
 sky130_fd_sc_hd__a31o_1 _0898_ (.A1(\flashBuffer.baseAddress[18] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net222),
    .B1(net199),
    .X(_0454_));
 sky130_fd_sc_hd__a31o_1 _0899_ (.A1(net179),
    .A2(_0453_),
    .A3(_0454_),
    .B1(net214),
    .X(_0455_));
 sky130_fd_sc_hd__a21o_1 _0900_ (.A1(net154),
    .A2(net184),
    .B1(_0455_),
    .X(_0122_));
 sky130_fd_sc_hd__a221o_2 _0901_ (.A1(net12),
    .A2(net189),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[19] ),
    .C1(net202),
    .X(_0456_));
 sky130_fd_sc_hd__a31o_1 _0902_ (.A1(\flashBuffer.baseAddress[19] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net223),
    .B1(net199),
    .X(_0457_));
 sky130_fd_sc_hd__a31o_1 _0903_ (.A1(net179),
    .A2(_0456_),
    .A3(_0457_),
    .B1(net214),
    .X(_0458_));
 sky130_fd_sc_hd__a21o_1 _0904_ (.A1(net155),
    .A2(net186),
    .B1(_0458_),
    .X(_0123_));
 sky130_fd_sc_hd__a221o_2 _0905_ (.A1(net14),
    .A2(net189),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[20] ),
    .C1(net202),
    .X(_0459_));
 sky130_fd_sc_hd__a31o_1 _0906_ (.A1(\flashBuffer.baseAddress[20] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net223),
    .B1(net199),
    .X(_0460_));
 sky130_fd_sc_hd__a31o_1 _0907_ (.A1(net179),
    .A2(_0459_),
    .A3(_0460_),
    .B1(net214),
    .X(_0461_));
 sky130_fd_sc_hd__a21o_1 _0908_ (.A1(net157),
    .A2(net186),
    .B1(_0461_),
    .X(_0124_));
 sky130_fd_sc_hd__a221o_2 _0909_ (.A1(net15),
    .A2(net190),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[21] ),
    .C1(_0387_),
    .X(_0462_));
 sky130_fd_sc_hd__a31o_1 _0910_ (.A1(\flashBuffer.baseAddress[21] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net222),
    .B1(net199),
    .X(_0463_));
 sky130_fd_sc_hd__a31o_1 _0911_ (.A1(net179),
    .A2(_0462_),
    .A3(_0463_),
    .B1(net215),
    .X(_0464_));
 sky130_fd_sc_hd__a21o_1 _0912_ (.A1(net158),
    .A2(net186),
    .B1(_0464_),
    .X(_0125_));
 sky130_fd_sc_hd__a221o_2 _0913_ (.A1(net16),
    .A2(net190),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[22] ),
    .C1(_0387_),
    .X(_0465_));
 sky130_fd_sc_hd__a31o_1 _0914_ (.A1(\flashBuffer.baseAddress[22] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net222),
    .B1(net199),
    .X(_0466_));
 sky130_fd_sc_hd__a31o_1 _0915_ (.A1(net180),
    .A2(_0465_),
    .A3(_0466_),
    .B1(net215),
    .X(_0467_));
 sky130_fd_sc_hd__a21o_1 _0916_ (.A1(net159),
    .A2(net186),
    .B1(_0467_),
    .X(_0126_));
 sky130_fd_sc_hd__a221o_2 _0917_ (.A1(net17),
    .A2(net190),
    .B1(_0446_),
    .B2(\flashBuffer.cachedAddress[23] ),
    .C1(_0387_),
    .X(_0468_));
 sky130_fd_sc_hd__a31o_1 _0918_ (.A1(\flashBuffer.baseAddress[23] ),
    .A2(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A3(net223),
    .B1(net199),
    .X(_0469_));
 sky130_fd_sc_hd__a31o_1 _0919_ (.A1(net179),
    .A2(_0468_),
    .A3(_0469_),
    .B1(net214),
    .X(_0470_));
 sky130_fd_sc_hd__a21o_1 _0920_ (.A1(net160),
    .A2(net187),
    .B1(_0470_),
    .X(_0127_));
 sky130_fd_sc_hd__a221o_1 _0921_ (.A1(net161),
    .A2(net184),
    .B1(_0393_),
    .B2(net18),
    .C1(net213),
    .X(_0128_));
 sky130_fd_sc_hd__a221o_1 _0922_ (.A1(net162),
    .A2(net184),
    .B1(_0393_),
    .B2(net19),
    .C1(net213),
    .X(_0129_));
 sky130_fd_sc_hd__a221o_1 _0923_ (.A1(net163),
    .A2(net184),
    .B1(_0393_),
    .B2(net20),
    .C1(net213),
    .X(_0130_));
 sky130_fd_sc_hd__a221o_1 _0924_ (.A1(net164),
    .A2(net185),
    .B1(_0393_),
    .B2(net21),
    .C1(net213),
    .X(_0131_));
 sky130_fd_sc_hd__a221o_1 _0925_ (.A1(net165),
    .A2(net184),
    .B1(_0393_),
    .B2(net22),
    .C1(net217),
    .X(_0132_));
 sky130_fd_sc_hd__a221o_1 _0926_ (.A1(net166),
    .A2(net184),
    .B1(_0393_),
    .B2(net23),
    .C1(net217),
    .X(_0133_));
 sky130_fd_sc_hd__a221o_1 _0927_ (.A1(net168),
    .A2(net184),
    .B1(_0393_),
    .B2(net25),
    .C1(net217),
    .X(_0134_));
 sky130_fd_sc_hd__a221o_1 _0928_ (.A1(net169),
    .A2(net186),
    .B1(_0393_),
    .B2(net26),
    .C1(net217),
    .X(_0135_));
 sky130_fd_sc_hd__o21ba_1 _0929_ (.A1(net144),
    .A2(_0389_),
    .B1_N(net213),
    .X(_0136_));
 sky130_fd_sc_hd__nand2_1 _0930_ (.A(net85),
    .B(net56),
    .Y(_0471_));
 sky130_fd_sc_hd__o21a_1 _0931_ (.A1(\wbPeripheralBusInterface.state[1] ),
    .A2(_0471_),
    .B1(_0395_),
    .X(_0472_));
 sky130_fd_sc_hd__nor2_1 _0932_ (.A(net237),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__o21a_1 _0933_ (.A1(net177),
    .A2(_0177_),
    .B1(_0473_),
    .X(_0137_));
 sky130_fd_sc_hd__and3b_2 _0934_ (.A_N(_0471_),
    .B(net228),
    .C(_0177_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(\wbPeripheralBusInterface.currentAddress[2] ),
    .A1(net48),
    .S(net212),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(\wbPeripheralBusInterface.currentAddress[3] ),
    .A1(net49),
    .S(net212),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(\wbPeripheralBusInterface.currentAddress[4] ),
    .A1(net50),
    .S(net212),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(\wbPeripheralBusInterface.currentAddress[5] ),
    .A1(net51),
    .S(net212),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0939_ (.A0(\wbPeripheralBusInterface.currentAddress[6] ),
    .A1(net52),
    .S(net212),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(\wbPeripheralBusInterface.currentAddress[7] ),
    .A1(net53),
    .S(net212),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0941_ (.A0(\wbPeripheralBusInterface.currentAddress[8] ),
    .A1(net54),
    .S(net212),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(\wbPeripheralBusInterface.currentAddress[9] ),
    .A1(net55),
    .S(net210),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0943_ (.A0(\wbPeripheralBusInterface.currentAddress[10] ),
    .A1(net34),
    .S(net210),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(\wbPeripheralBusInterface.currentAddress[11] ),
    .A1(net35),
    .S(net210),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0945_ (.A0(\wbPeripheralBusInterface.currentAddress[12] ),
    .A1(net36),
    .S(net210),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(\wbPeripheralBusInterface.currentAddress[13] ),
    .A1(net37),
    .S(net210),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0947_ (.A0(\wbPeripheralBusInterface.currentAddress[14] ),
    .A1(net38),
    .S(net210),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(\wbPeripheralBusInterface.currentAddress[15] ),
    .A1(net39),
    .S(net210),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0949_ (.A0(\wbPeripheralBusInterface.currentAddress[16] ),
    .A1(net40),
    .S(net210),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(\wbPeripheralBusInterface.currentAddress[17] ),
    .A1(net41),
    .S(net210),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0951_ (.A0(\wbPeripheralBusInterface.currentAddress[18] ),
    .A1(net42),
    .S(net211),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(\wbPeripheralBusInterface.currentAddress[19] ),
    .A1(net43),
    .S(net211),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(\wbPeripheralBusInterface.currentAddress[20] ),
    .A1(net44),
    .S(net211),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(\wbPeripheralBusInterface.currentAddress[21] ),
    .A1(net45),
    .S(net211),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _0955_ (.A0(\wbPeripheralBusInterface.currentAddress[22] ),
    .A1(net46),
    .S(net211),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(\wbPeripheralBusInterface.currentAddress[23] ),
    .A1(net47),
    .S(net211),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _0957_ (.A(\qspiDevice.outputClock ),
    .B(net232),
    .X(_0160_));
 sky130_fd_sc_hd__o211a_1 _0958_ (.A1(net86),
    .A2(net220),
    .B1(_0389_),
    .C1(_0473_),
    .X(_0161_));
 sky130_fd_sc_hd__a21boi_1 _0959_ (.A1(net86),
    .A2(_0177_),
    .B1_N(_0473_),
    .Y(_0162_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(net225),
    .A1(net82),
    .S(net212),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .A1(net83),
    .S(net212),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A1(net84),
    .S(net210),
    .X(_0165_));
 sky130_fd_sc_hd__dfxtp_2 _0963_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0000_),
    .Q(\flashBuffer.qspi_requestData ));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0001_),
    .Q(\flashBuffer.cachedCount[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0002_),
    .Q(\flashBuffer.cachedCount[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0003_),
    .Q(\flashBuffer.cachedCount[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0004_),
    .Q(\flashBuffer.cachedCount[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0005_),
    .Q(\flashBuffer.cachedCount[4] ));
 sky130_fd_sc_hd__dfxtp_2 _0969_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0006_),
    .Q(\flashBuffer.cachedCount[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0007_),
    .Q(\flashBuffer.cachedCount[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0008_),
    .Q(\flashBuffer.cachedCount[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0009_),
    .Q(\flashBuffer.cachedCount[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0010_),
    .Q(\flashBuffer.cachedCount[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0974_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0011_),
    .Q(\flashBuffer.baseAddress[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0012_),
    .Q(\flashBuffer.baseAddress[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0976_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0013_),
    .Q(\flashBuffer.baseAddress[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0977_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0014_),
    .Q(\flashBuffer.baseAddress[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0015_),
    .Q(\flashBuffer.baseAddress[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0016_),
    .Q(\flashBuffer.baseAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0017_),
    .Q(\flashBuffer.baseAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0018_),
    .Q(\flashBuffer.baseAddress[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0019_),
    .Q(\flashBuffer.baseAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0020_),
    .Q(\flashBuffer.baseAddress[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0021_),
    .Q(\flashBuffer.baseAddress[10] ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0022_),
    .Q(\flashBuffer.baseAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0023_),
    .Q(\flashBuffer.baseAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0024_),
    .Q(\flashBuffer.baseAddress[13] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0025_),
    .Q(\flashBuffer.baseAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0026_),
    .Q(\flashBuffer.baseAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0027_),
    .Q(\flashBuffer.baseAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0028_),
    .Q(\flashBuffer.baseAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0029_),
    .Q(\flashBuffer.baseAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0030_),
    .Q(\flashBuffer.baseAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0031_),
    .Q(\flashBuffer.baseAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0032_),
    .Q(\flashBuffer.baseAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0033_),
    .Q(\flashBuffer.baseAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0034_),
    .Q(\flashBuffer.baseAddress[23] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0035_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0036_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0037_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0038_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_2 _1002_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0039_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_2 _1003_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0040_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0041_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_2 _1005_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0042_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0043_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0044_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0045_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0046_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0047_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0048_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0049_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_2 _1013_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0050_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_2 _1014_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0051_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_2 _1015_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0052_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0053_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0054_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0055_),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0056_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0057_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0058_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_2 _1022_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0059_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_2 _1023_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0060_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_2 _1024_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0061_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_2 _1025_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0062_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_2 _1026_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0063_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0064_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0065_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_2 _1029_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0066_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0067_),
    .Q(\qspiDevice.register.outputBit ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0068_),
    .Q(\qspiDevice.resetState[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0069_),
    .Q(\qspiDevice.resetState[1] ));
 sky130_fd_sc_hd__dfxtp_4 _1033_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0070_),
    .Q(\qspiDevice.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1034_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0071_),
    .Q(\qspiDevice.state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _1035_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0072_),
    .Q(\flashBuffer.qspi_readDataValid ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0073_),
    .Q(\flashBuffer.flashCacheReadReady ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0074_),
    .Q(\qspiDevice.settingAddress ));
 sky130_fd_sc_hd__dfxtp_4 _1038_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0075_),
    .Q(\qspiDevice.outputClock ));
 sky130_fd_sc_hd__dfxtp_2 _1039_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0076_),
    .Q(\qspiDevice.bitCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0077_),
    .Q(\qspiDevice.bitCounter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1041_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0078_),
    .Q(\qspiDevice.bitCounter[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1042_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0079_),
    .Q(\qspiDevice.bitCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0080_),
    .Q(\qspiDevice.bitCounter[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1044_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0081_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _1045_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0082_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _1046_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0083_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_2 _1047_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0084_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0085_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _1049_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0086_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _1050_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0087_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0088_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_2 _1052_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0089_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0090_),
    .Q(\flashBuffer.cachedAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0091_),
    .Q(\flashBuffer.cachedAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0092_),
    .Q(\flashBuffer.cachedAddress[13] ));
 sky130_fd_sc_hd__dfxtp_2 _1056_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0093_),
    .Q(\flashBuffer.cachedAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0094_),
    .Q(\flashBuffer.cachedAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0095_),
    .Q(\flashBuffer.cachedAddress[16] ));
 sky130_fd_sc_hd__dfxtp_2 _1059_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0096_),
    .Q(\flashBuffer.cachedAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0097_),
    .Q(\flashBuffer.cachedAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0098_),
    .Q(\flashBuffer.cachedAddress[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1062_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0099_),
    .Q(\flashBuffer.cachedAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0100_),
    .Q(\flashBuffer.cachedAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0101_),
    .Q(\flashBuffer.cachedAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0102_),
    .Q(\flashBuffer.cachedAddress[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1066_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0103_),
    .Q(\flashBuffer.configuration ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0104_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0105_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0106_),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0107_),
    .Q(net170));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0108_),
    .Q(net171));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0109_),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0110_),
    .Q(net173));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0111_),
    .Q(net174));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0112_),
    .Q(net175));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0113_),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0114_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_2 _1078_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0115_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_2 _1079_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0116_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0117_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0118_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0119_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0120_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0121_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0122_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0123_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_2 _1087_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0124_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_2 _1088_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0125_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_2 _1089_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0126_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_2 _1090_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0127_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_2 _1091_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0128_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_2 _1092_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0129_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_2 _1093_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0130_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_2 _1094_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0131_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_2 _1095_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0132_),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_2 _1096_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0133_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_2 _1097_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0134_),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_2 _1098_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0135_),
    .Q(net169));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0136_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0137_),
    .Q(net177));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0138_),
    .Q(\wbPeripheralBusInterface.currentAddress[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0139_),
    .Q(\wbPeripheralBusInterface.currentAddress[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0140_),
    .Q(\wbPeripheralBusInterface.currentAddress[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0141_),
    .Q(\wbPeripheralBusInterface.currentAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0142_),
    .Q(\wbPeripheralBusInterface.currentAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0143_),
    .Q(\wbPeripheralBusInterface.currentAddress[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0144_),
    .Q(\wbPeripheralBusInterface.currentAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0145_),
    .Q(\wbPeripheralBusInterface.currentAddress[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0146_),
    .Q(\wbPeripheralBusInterface.currentAddress[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0147_),
    .Q(\wbPeripheralBusInterface.currentAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0148_),
    .Q(\wbPeripheralBusInterface.currentAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0149_),
    .Q(\wbPeripheralBusInterface.currentAddress[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0150_),
    .Q(\wbPeripheralBusInterface.currentAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0151_),
    .Q(\wbPeripheralBusInterface.currentAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0152_),
    .Q(\wbPeripheralBusInterface.currentAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0153_),
    .Q(\wbPeripheralBusInterface.currentAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0154_),
    .Q(\wbPeripheralBusInterface.currentAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0155_),
    .Q(\wbPeripheralBusInterface.currentAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0156_),
    .Q(\wbPeripheralBusInterface.currentAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0157_),
    .Q(\wbPeripheralBusInterface.currentAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0158_),
    .Q(\wbPeripheralBusInterface.currentAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0159_),
    .Q(\wbPeripheralBusInterface.currentAddress[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1123_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0160_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _1124_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0161_),
    .Q(\wbPeripheralBusInterface.state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1125_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0162_),
    .Q(\wbPeripheralBusInterface.state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1126_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0163_),
    .Q(\wbPeripheralBusInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1127_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0164_),
    .Q(\wbPeripheralBusInterface.currentByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_4 _1128_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0165_),
    .Q(\wbPeripheralBusInterface.currentByteSelect[2] ));
 sky130_fd_sc_hd__buf_2 _1138_ (.A(clknet_4_0_0_wb_clk_i),
    .X(net108));
 sky130_fd_sc_hd__buf_2 _1139_ (.A(clknet_4_0_0_wb_clk_i),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(_0261_),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(_0392_),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_0253_),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(_0253_),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_6 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_6 fanout186 (.A(_0390_),
    .X(net186));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(_0390_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(net190),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(_0386_),
    .X(net190));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__buf_2 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(_0242_),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net197),
    .X(net194));
 sky130_fd_sc_hd__buf_4 fanout195 (.A(net197),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(_0197_),
    .X(net197));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(_0197_),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(_0388_),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(_0387_),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(_0387_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_6 fanout205 (.A(net208),
    .X(net205));
 sky130_fd_sc_hd__buf_6 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_6 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_6 fanout208 (.A(_0196_),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(_0248_),
    .X(net209));
 sky130_fd_sc_hd__buf_6 fanout210 (.A(_0474_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_6 fanout212 (.A(_0474_),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net217),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_4 fanout217 (.A(_0396_),
    .X(net217));
 sky130_fd_sc_hd__buf_6 fanout218 (.A(_0244_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(_0244_),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_4 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(_0178_),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(_0178_),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(\wbPeripheralBusInterface.currentByteSelect[0] ),
    .X(net225));
 sky130_fd_sc_hd__buf_6 fanout226 (.A(\qspiDevice.state[1] ),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_8 fanout227 (.A(\qspiDevice.state[0] ),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net233),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net233),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 fanout233 (.A(_0176_),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net236),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_6 fanout236 (.A(net81),
    .X(net236));
 sky130_fd_sc_hd__buf_6 fanout237 (.A(net81),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(flash_io1_read),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(sram_dout1[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(sram_dout1[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(sram_dout1[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(sram_dout1[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(sram_dout1[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(sram_dout1[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(sram_dout1[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(sram_dout1[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(sram_dout1[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(sram_dout1[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(sram_dout1[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(sram_dout1[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(sram_dout1[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(sram_dout1[28]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(sram_dout1[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(sram_dout1[2]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(sram_dout1[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(sram_dout1[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(sram_dout1[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(sram_dout1[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(sram_dout1[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(sram_dout1[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(sram_dout1[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(sram_dout1[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(sram_dout1[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(sram_dout1[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(wb_adr_i[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(wb_adr_i[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(wb_adr_i[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(wb_adr_i[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(wb_adr_i[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(wb_adr_i[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(sram_dout1[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(wb_adr_i[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(wb_adr_i[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(wb_adr_i[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(wb_adr_i[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(wb_adr_i[20]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(wb_adr_i[21]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(wb_adr_i[22]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(wb_adr_i[23]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(wb_adr_i[2]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(wb_adr_i[3]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(sram_dout1[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(wb_adr_i[4]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(wb_adr_i[5]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(wb_adr_i[6]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(wb_adr_i[7]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(wb_adr_i[8]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(wb_adr_i[9]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(wb_cyc_i),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(wb_data_i[0]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(wb_data_i[10]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(wb_data_i[11]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(sram_dout1[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(wb_data_i[12]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(wb_data_i[13]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(wb_data_i[14]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(wb_data_i[15]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(wb_data_i[16]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(wb_data_i[17]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input66 (.A(wb_data_i[18]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(wb_data_i[19]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(wb_data_i[1]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(wb_data_i[20]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(sram_dout1[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(wb_data_i[21]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(wb_data_i[22]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(wb_data_i[23]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(wb_data_i[2]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(wb_data_i[3]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(wb_data_i[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(wb_data_i[5]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(wb_data_i[6]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(wb_data_i[7]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(wb_data_i[8]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(sram_dout1[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(wb_data_i[9]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(wb_rst_i),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(wb_sel_i[0]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(wb_sel_i[1]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(wb_sel_i[2]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(wb_stb_i),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(wb_we_i),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(sram_dout1[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 output100 (.A(net100),
    .X(sram_addr1[1]));
 sky130_fd_sc_hd__buf_4 output101 (.A(net101),
    .X(sram_addr1[2]));
 sky130_fd_sc_hd__buf_4 output102 (.A(net102),
    .X(sram_addr1[3]));
 sky130_fd_sc_hd__buf_4 output103 (.A(net103),
    .X(sram_addr1[4]));
 sky130_fd_sc_hd__buf_4 output104 (.A(net104),
    .X(sram_addr1[5]));
 sky130_fd_sc_hd__buf_4 output105 (.A(net105),
    .X(sram_addr1[6]));
 sky130_fd_sc_hd__buf_4 output106 (.A(net106),
    .X(sram_addr1[7]));
 sky130_fd_sc_hd__buf_4 output107 (.A(net107),
    .X(sram_addr1[8]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(sram_clk0));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(sram_clk1));
 sky130_fd_sc_hd__buf_4 output110 (.A(net110),
    .X(sram_csb0));
 sky130_fd_sc_hd__buf_4 output111 (.A(net111),
    .X(sram_csb1));
 sky130_fd_sc_hd__buf_4 output112 (.A(net112),
    .X(sram_din0[0]));
 sky130_fd_sc_hd__buf_4 output113 (.A(net113),
    .X(sram_din0[10]));
 sky130_fd_sc_hd__buf_4 output114 (.A(net114),
    .X(sram_din0[11]));
 sky130_fd_sc_hd__buf_4 output115 (.A(net115),
    .X(sram_din0[12]));
 sky130_fd_sc_hd__buf_4 output116 (.A(net116),
    .X(sram_din0[13]));
 sky130_fd_sc_hd__buf_4 output117 (.A(net117),
    .X(sram_din0[14]));
 sky130_fd_sc_hd__buf_4 output118 (.A(net118),
    .X(sram_din0[15]));
 sky130_fd_sc_hd__buf_4 output119 (.A(net119),
    .X(sram_din0[16]));
 sky130_fd_sc_hd__buf_4 output120 (.A(net120),
    .X(sram_din0[17]));
 sky130_fd_sc_hd__buf_4 output121 (.A(net121),
    .X(sram_din0[18]));
 sky130_fd_sc_hd__buf_4 output122 (.A(net122),
    .X(sram_din0[19]));
 sky130_fd_sc_hd__buf_4 output123 (.A(net123),
    .X(sram_din0[1]));
 sky130_fd_sc_hd__buf_4 output124 (.A(net124),
    .X(sram_din0[20]));
 sky130_fd_sc_hd__buf_4 output125 (.A(net125),
    .X(sram_din0[21]));
 sky130_fd_sc_hd__buf_4 output126 (.A(net126),
    .X(sram_din0[22]));
 sky130_fd_sc_hd__buf_4 output127 (.A(net127),
    .X(sram_din0[23]));
 sky130_fd_sc_hd__buf_4 output128 (.A(net128),
    .X(sram_din0[24]));
 sky130_fd_sc_hd__buf_4 output129 (.A(net129),
    .X(sram_din0[25]));
 sky130_fd_sc_hd__buf_4 output130 (.A(net130),
    .X(sram_din0[26]));
 sky130_fd_sc_hd__buf_4 output131 (.A(net131),
    .X(sram_din0[27]));
 sky130_fd_sc_hd__buf_4 output132 (.A(net132),
    .X(sram_din0[28]));
 sky130_fd_sc_hd__buf_4 output133 (.A(net133),
    .X(sram_din0[29]));
 sky130_fd_sc_hd__buf_4 output134 (.A(net134),
    .X(sram_din0[2]));
 sky130_fd_sc_hd__buf_4 output135 (.A(net135),
    .X(sram_din0[30]));
 sky130_fd_sc_hd__buf_4 output136 (.A(net136),
    .X(sram_din0[31]));
 sky130_fd_sc_hd__buf_4 output137 (.A(net137),
    .X(sram_din0[3]));
 sky130_fd_sc_hd__buf_4 output138 (.A(net138),
    .X(sram_din0[4]));
 sky130_fd_sc_hd__buf_4 output139 (.A(net139),
    .X(sram_din0[5]));
 sky130_fd_sc_hd__buf_4 output140 (.A(net140),
    .X(sram_din0[6]));
 sky130_fd_sc_hd__buf_4 output141 (.A(net141),
    .X(sram_din0[7]));
 sky130_fd_sc_hd__buf_4 output142 (.A(net142),
    .X(sram_din0[8]));
 sky130_fd_sc_hd__buf_4 output143 (.A(net143),
    .X(sram_din0[9]));
 sky130_fd_sc_hd__buf_4 output144 (.A(net144),
    .X(wb_ack_o));
 sky130_fd_sc_hd__buf_4 output145 (.A(net145),
    .X(wb_data_o[0]));
 sky130_fd_sc_hd__buf_4 output146 (.A(net146),
    .X(wb_data_o[10]));
 sky130_fd_sc_hd__buf_4 output147 (.A(net147),
    .X(wb_data_o[11]));
 sky130_fd_sc_hd__buf_4 output148 (.A(net148),
    .X(wb_data_o[12]));
 sky130_fd_sc_hd__buf_4 output149 (.A(net149),
    .X(wb_data_o[13]));
 sky130_fd_sc_hd__buf_4 output150 (.A(net150),
    .X(wb_data_o[14]));
 sky130_fd_sc_hd__buf_4 output151 (.A(net151),
    .X(wb_data_o[15]));
 sky130_fd_sc_hd__buf_4 output152 (.A(net152),
    .X(wb_data_o[16]));
 sky130_fd_sc_hd__buf_4 output153 (.A(net153),
    .X(wb_data_o[17]));
 sky130_fd_sc_hd__buf_4 output154 (.A(net154),
    .X(wb_data_o[18]));
 sky130_fd_sc_hd__buf_4 output155 (.A(net155),
    .X(wb_data_o[19]));
 sky130_fd_sc_hd__buf_4 output156 (.A(net156),
    .X(wb_data_o[1]));
 sky130_fd_sc_hd__buf_4 output157 (.A(net157),
    .X(wb_data_o[20]));
 sky130_fd_sc_hd__buf_4 output158 (.A(net158),
    .X(wb_data_o[21]));
 sky130_fd_sc_hd__buf_4 output159 (.A(net159),
    .X(wb_data_o[22]));
 sky130_fd_sc_hd__buf_4 output160 (.A(net160),
    .X(wb_data_o[23]));
 sky130_fd_sc_hd__buf_4 output161 (.A(net161),
    .X(wb_data_o[24]));
 sky130_fd_sc_hd__buf_4 output162 (.A(net162),
    .X(wb_data_o[25]));
 sky130_fd_sc_hd__buf_4 output163 (.A(net163),
    .X(wb_data_o[26]));
 sky130_fd_sc_hd__buf_4 output164 (.A(net164),
    .X(wb_data_o[27]));
 sky130_fd_sc_hd__buf_4 output165 (.A(net165),
    .X(wb_data_o[28]));
 sky130_fd_sc_hd__buf_4 output166 (.A(net166),
    .X(wb_data_o[29]));
 sky130_fd_sc_hd__buf_4 output167 (.A(net167),
    .X(wb_data_o[2]));
 sky130_fd_sc_hd__buf_4 output168 (.A(net168),
    .X(wb_data_o[30]));
 sky130_fd_sc_hd__buf_4 output169 (.A(net169),
    .X(wb_data_o[31]));
 sky130_fd_sc_hd__buf_4 output170 (.A(net170),
    .X(wb_data_o[3]));
 sky130_fd_sc_hd__buf_4 output171 (.A(net171),
    .X(wb_data_o[4]));
 sky130_fd_sc_hd__buf_4 output172 (.A(net172),
    .X(wb_data_o[5]));
 sky130_fd_sc_hd__buf_4 output173 (.A(net173),
    .X(wb_data_o[6]));
 sky130_fd_sc_hd__buf_4 output174 (.A(net174),
    .X(wb_data_o[7]));
 sky130_fd_sc_hd__buf_4 output175 (.A(net175),
    .X(wb_data_o[8]));
 sky130_fd_sc_hd__buf_4 output176 (.A(net176),
    .X(wb_data_o[9]));
 sky130_fd_sc_hd__buf_4 output177 (.A(net177),
    .X(wb_stall_o));
 sky130_fd_sc_hd__buf_4 output87 (.A(net87),
    .X(flash_csb));
 sky130_fd_sc_hd__buf_4 output88 (.A(net88),
    .X(flash_io0_write));
 sky130_fd_sc_hd__buf_4 output89 (.A(net89),
    .X(flash_sck));
 sky130_fd_sc_hd__buf_4 output90 (.A(net90),
    .X(sram_addr0[0]));
 sky130_fd_sc_hd__buf_4 output91 (.A(net91),
    .X(sram_addr0[1]));
 sky130_fd_sc_hd__buf_4 output92 (.A(net92),
    .X(sram_addr0[2]));
 sky130_fd_sc_hd__buf_4 output93 (.A(net93),
    .X(sram_addr0[3]));
 sky130_fd_sc_hd__buf_4 output94 (.A(net94),
    .X(sram_addr0[4]));
 sky130_fd_sc_hd__buf_4 output95 (.A(net95),
    .X(sram_addr0[5]));
 sky130_fd_sc_hd__buf_4 output96 (.A(net96),
    .X(sram_addr0[6]));
 sky130_fd_sc_hd__buf_4 output97 (.A(net97),
    .X(sram_addr0[7]));
 sky130_fd_sc_hd__buf_4 output98 (.A(net98),
    .X(sram_addr0[8]));
 sky130_fd_sc_hd__buf_4 output99 (.A(net99),
    .X(sram_addr1[0]));
 assign flash_io0_we = net242;
 assign flash_io1_we = net238;
 assign flash_io1_write = net239;
 assign sram_web0 = net240;
 assign sram_wmask0[0] = net243;
 assign sram_wmask0[1] = net244;
 assign sram_wmask0[2] = net245;
 assign sram_wmask0[3] = net246;
 assign wb_error_o = net241;
endmodule

