VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 950.000 ;
  PIN flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END flash_csb
  PIN flash_io0_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END flash_io0_read
  PIN flash_io0_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END flash_io0_we
  PIN flash_io0_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END flash_io0_write
  PIN flash_io1_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END flash_io1_read
  PIN flash_io1_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END flash_io1_we
  PIN flash_io1_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END flash_io1_write
  PIN flash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END flash_sck
  PIN internal_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END internal_uart_rx
  PIN internal_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END internal_uart_tx
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 946.000 4.050 950.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 946.000 81.790 950.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 946.000 89.610 950.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 946.000 97.430 950.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 946.000 105.250 950.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 946.000 113.070 950.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 946.000 120.890 950.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 946.000 128.250 950.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 946.000 136.070 950.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 946.000 143.890 950.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 946.000 151.710 950.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 946.000 11.410 950.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 946.000 159.530 950.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 946.000 167.350 950.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 946.000 175.170 950.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 946.000 182.990 950.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 946.000 190.810 950.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 946.000 198.630 950.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 946.000 206.450 950.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 946.000 214.270 950.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 946.000 222.090 950.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 946.000 229.910 950.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 946.000 19.230 950.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 946.000 237.730 950.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 946.000 245.090 950.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 946.000 252.910 950.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 946.000 260.730 950.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 946.000 268.550 950.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 946.000 276.370 950.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 946.000 284.190 950.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 946.000 292.010 950.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 946.000 27.050 950.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 946.000 34.870 950.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 946.000 42.690 950.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 946.000 50.510 950.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 946.000 58.330 950.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 946.000 66.150 950.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 946.000 73.970 950.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 946.000 299.830 950.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 946.000 377.570 950.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 946.000 385.390 950.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 946.000 393.210 950.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 946.000 401.030 950.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 946.000 408.850 950.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 946.000 416.670 950.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 946.000 424.490 950.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 946.000 432.310 950.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 946.000 440.130 950.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 946.000 447.950 950.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 946.000 307.650 950.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 946.000 455.770 950.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 946.000 463.590 950.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 946.000 471.410 950.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 946.000 479.230 950.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 946.000 486.590 950.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 946.000 494.410 950.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 946.000 502.230 950.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 946.000 510.050 950.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 946.000 517.870 950.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 946.000 525.690 950.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 946.000 315.470 950.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 946.000 533.510 950.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 946.000 541.330 950.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 946.000 549.150 950.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 946.000 556.970 950.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 946.000 564.790 950.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 946.000 572.610 950.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 946.000 580.430 950.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 946.000 588.250 950.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 946.000 323.290 950.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 946.000 331.110 950.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 946.000 338.930 950.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 946.000 346.750 950.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 946.000 354.570 950.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 946.000 362.390 950.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 946.000 369.750 950.000 ;
    END
  END io_out[9]
  PIN jtag_tck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 395.120 600.000 395.720 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 553.560 600.000 554.160 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 712.000 600.000 712.600 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 870.440 600.000 871.040 ;
    END
  END jtag_tms
  PIN peripheral_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 946.000 596.070 950.000 ;
    END
  END peripheral_irq[0]
  PIN peripheral_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END peripheral_irq[1]
  PIN peripheral_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 917.360 4.000 917.960 ;
    END
  END peripheral_irq[2]
  PIN peripheral_irq[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.200 4.000 926.800 ;
    END
  END peripheral_irq[3]
  PIN peripheral_irq[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END peripheral_irq[4]
  PIN peripheral_irq[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END peripheral_irq[5]
  PIN peripheral_irq[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END peripheral_irq[6]
  PIN peripheral_irq[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.720 4.000 936.320 ;
    END
  END peripheral_irq[7]
  PIN peripheral_irq[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END peripheral_irq[8]
  PIN peripheral_irq[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END peripheral_irq[9]
  PIN probe_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 78.920 600.000 79.520 ;
    END
  END probe_blink[0]
  PIN probe_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 236.680 600.000 237.280 ;
    END
  END probe_blink[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 938.640 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 938.640 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 551.520 4.000 552.120 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.680 4.000 662.280 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.800 4.000 753.400 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.920 4.000 844.520 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.960 4.000 625.560 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 4.000 780.600 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 798.360 4.000 798.960 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.720 4.000 817.320 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.800 4.000 872.400 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 938.485 ;
      LAYER met1 ;
        RECT 0.070 9.220 596.090 939.040 ;
      LAYER met2 ;
        RECT 0.100 945.720 3.490 946.290 ;
        RECT 4.330 945.720 10.850 946.290 ;
        RECT 11.690 945.720 18.670 946.290 ;
        RECT 19.510 945.720 26.490 946.290 ;
        RECT 27.330 945.720 34.310 946.290 ;
        RECT 35.150 945.720 42.130 946.290 ;
        RECT 42.970 945.720 49.950 946.290 ;
        RECT 50.790 945.720 57.770 946.290 ;
        RECT 58.610 945.720 65.590 946.290 ;
        RECT 66.430 945.720 73.410 946.290 ;
        RECT 74.250 945.720 81.230 946.290 ;
        RECT 82.070 945.720 89.050 946.290 ;
        RECT 89.890 945.720 96.870 946.290 ;
        RECT 97.710 945.720 104.690 946.290 ;
        RECT 105.530 945.720 112.510 946.290 ;
        RECT 113.350 945.720 120.330 946.290 ;
        RECT 121.170 945.720 127.690 946.290 ;
        RECT 128.530 945.720 135.510 946.290 ;
        RECT 136.350 945.720 143.330 946.290 ;
        RECT 144.170 945.720 151.150 946.290 ;
        RECT 151.990 945.720 158.970 946.290 ;
        RECT 159.810 945.720 166.790 946.290 ;
        RECT 167.630 945.720 174.610 946.290 ;
        RECT 175.450 945.720 182.430 946.290 ;
        RECT 183.270 945.720 190.250 946.290 ;
        RECT 191.090 945.720 198.070 946.290 ;
        RECT 198.910 945.720 205.890 946.290 ;
        RECT 206.730 945.720 213.710 946.290 ;
        RECT 214.550 945.720 221.530 946.290 ;
        RECT 222.370 945.720 229.350 946.290 ;
        RECT 230.190 945.720 237.170 946.290 ;
        RECT 238.010 945.720 244.530 946.290 ;
        RECT 245.370 945.720 252.350 946.290 ;
        RECT 253.190 945.720 260.170 946.290 ;
        RECT 261.010 945.720 267.990 946.290 ;
        RECT 268.830 945.720 275.810 946.290 ;
        RECT 276.650 945.720 283.630 946.290 ;
        RECT 284.470 945.720 291.450 946.290 ;
        RECT 292.290 945.720 299.270 946.290 ;
        RECT 300.110 945.720 307.090 946.290 ;
        RECT 307.930 945.720 314.910 946.290 ;
        RECT 315.750 945.720 322.730 946.290 ;
        RECT 323.570 945.720 330.550 946.290 ;
        RECT 331.390 945.720 338.370 946.290 ;
        RECT 339.210 945.720 346.190 946.290 ;
        RECT 347.030 945.720 354.010 946.290 ;
        RECT 354.850 945.720 361.830 946.290 ;
        RECT 362.670 945.720 369.190 946.290 ;
        RECT 370.030 945.720 377.010 946.290 ;
        RECT 377.850 945.720 384.830 946.290 ;
        RECT 385.670 945.720 392.650 946.290 ;
        RECT 393.490 945.720 400.470 946.290 ;
        RECT 401.310 945.720 408.290 946.290 ;
        RECT 409.130 945.720 416.110 946.290 ;
        RECT 416.950 945.720 423.930 946.290 ;
        RECT 424.770 945.720 431.750 946.290 ;
        RECT 432.590 945.720 439.570 946.290 ;
        RECT 440.410 945.720 447.390 946.290 ;
        RECT 448.230 945.720 455.210 946.290 ;
        RECT 456.050 945.720 463.030 946.290 ;
        RECT 463.870 945.720 470.850 946.290 ;
        RECT 471.690 945.720 478.670 946.290 ;
        RECT 479.510 945.720 486.030 946.290 ;
        RECT 486.870 945.720 493.850 946.290 ;
        RECT 494.690 945.720 501.670 946.290 ;
        RECT 502.510 945.720 509.490 946.290 ;
        RECT 510.330 945.720 517.310 946.290 ;
        RECT 518.150 945.720 525.130 946.290 ;
        RECT 525.970 945.720 532.950 946.290 ;
        RECT 533.790 945.720 540.770 946.290 ;
        RECT 541.610 945.720 548.590 946.290 ;
        RECT 549.430 945.720 556.410 946.290 ;
        RECT 557.250 945.720 564.230 946.290 ;
        RECT 565.070 945.720 572.050 946.290 ;
        RECT 572.890 945.720 579.870 946.290 ;
        RECT 580.710 945.720 587.690 946.290 ;
        RECT 588.530 945.720 595.510 946.290 ;
        RECT 0.100 4.280 596.060 945.720 ;
        RECT 0.100 4.000 4.410 4.280 ;
        RECT 5.250 4.000 14.070 4.280 ;
        RECT 14.910 4.000 23.730 4.280 ;
        RECT 24.570 4.000 33.850 4.280 ;
        RECT 34.690 4.000 43.510 4.280 ;
        RECT 44.350 4.000 53.170 4.280 ;
        RECT 54.010 4.000 63.290 4.280 ;
        RECT 64.130 4.000 72.950 4.280 ;
        RECT 73.790 4.000 83.070 4.280 ;
        RECT 83.910 4.000 92.730 4.280 ;
        RECT 93.570 4.000 102.390 4.280 ;
        RECT 103.230 4.000 112.510 4.280 ;
        RECT 113.350 4.000 122.170 4.280 ;
        RECT 123.010 4.000 131.830 4.280 ;
        RECT 132.670 4.000 141.950 4.280 ;
        RECT 142.790 4.000 151.610 4.280 ;
        RECT 152.450 4.000 161.730 4.280 ;
        RECT 162.570 4.000 171.390 4.280 ;
        RECT 172.230 4.000 181.050 4.280 ;
        RECT 181.890 4.000 191.170 4.280 ;
        RECT 192.010 4.000 200.830 4.280 ;
        RECT 201.670 4.000 210.490 4.280 ;
        RECT 211.330 4.000 220.610 4.280 ;
        RECT 221.450 4.000 230.270 4.280 ;
        RECT 231.110 4.000 240.390 4.280 ;
        RECT 241.230 4.000 250.050 4.280 ;
        RECT 250.890 4.000 259.710 4.280 ;
        RECT 260.550 4.000 269.830 4.280 ;
        RECT 270.670 4.000 279.490 4.280 ;
        RECT 280.330 4.000 289.150 4.280 ;
        RECT 289.990 4.000 299.270 4.280 ;
        RECT 300.110 4.000 308.930 4.280 ;
        RECT 309.770 4.000 319.050 4.280 ;
        RECT 319.890 4.000 328.710 4.280 ;
        RECT 329.550 4.000 338.370 4.280 ;
        RECT 339.210 4.000 348.490 4.280 ;
        RECT 349.330 4.000 358.150 4.280 ;
        RECT 358.990 4.000 367.810 4.280 ;
        RECT 368.650 4.000 377.930 4.280 ;
        RECT 378.770 4.000 387.590 4.280 ;
        RECT 388.430 4.000 397.710 4.280 ;
        RECT 398.550 4.000 407.370 4.280 ;
        RECT 408.210 4.000 417.030 4.280 ;
        RECT 417.870 4.000 427.150 4.280 ;
        RECT 427.990 4.000 436.810 4.280 ;
        RECT 437.650 4.000 446.470 4.280 ;
        RECT 447.310 4.000 456.590 4.280 ;
        RECT 457.430 4.000 466.250 4.280 ;
        RECT 467.090 4.000 476.370 4.280 ;
        RECT 477.210 4.000 486.030 4.280 ;
        RECT 486.870 4.000 495.690 4.280 ;
        RECT 496.530 4.000 505.810 4.280 ;
        RECT 506.650 4.000 515.470 4.280 ;
        RECT 516.310 4.000 525.130 4.280 ;
        RECT 525.970 4.000 535.250 4.280 ;
        RECT 536.090 4.000 544.910 4.280 ;
        RECT 545.750 4.000 555.030 4.280 ;
        RECT 555.870 4.000 564.690 4.280 ;
        RECT 565.530 4.000 574.350 4.280 ;
        RECT 575.190 4.000 584.470 4.280 ;
        RECT 585.310 4.000 594.130 4.280 ;
        RECT 594.970 4.000 596.060 4.280 ;
      LAYER met3 ;
        RECT 4.400 944.160 596.000 945.025 ;
        RECT 4.000 936.720 596.000 944.160 ;
        RECT 4.400 935.320 596.000 936.720 ;
        RECT 4.000 927.200 596.000 935.320 ;
        RECT 4.400 925.800 596.000 927.200 ;
        RECT 4.000 918.360 596.000 925.800 ;
        RECT 4.400 916.960 596.000 918.360 ;
        RECT 4.000 908.840 596.000 916.960 ;
        RECT 4.400 907.440 596.000 908.840 ;
        RECT 4.000 900.000 596.000 907.440 ;
        RECT 4.400 898.600 596.000 900.000 ;
        RECT 4.000 890.480 596.000 898.600 ;
        RECT 4.400 889.080 596.000 890.480 ;
        RECT 4.000 881.640 596.000 889.080 ;
        RECT 4.400 880.240 596.000 881.640 ;
        RECT 4.000 872.800 596.000 880.240 ;
        RECT 4.400 871.440 596.000 872.800 ;
        RECT 4.400 871.400 595.600 871.440 ;
        RECT 4.000 870.040 595.600 871.400 ;
        RECT 4.000 863.280 596.000 870.040 ;
        RECT 4.400 861.880 596.000 863.280 ;
        RECT 4.000 854.440 596.000 861.880 ;
        RECT 4.400 853.040 596.000 854.440 ;
        RECT 4.000 844.920 596.000 853.040 ;
        RECT 4.400 843.520 596.000 844.920 ;
        RECT 4.000 836.080 596.000 843.520 ;
        RECT 4.400 834.680 596.000 836.080 ;
        RECT 4.000 826.560 596.000 834.680 ;
        RECT 4.400 825.160 596.000 826.560 ;
        RECT 4.000 817.720 596.000 825.160 ;
        RECT 4.400 816.320 596.000 817.720 ;
        RECT 4.000 808.880 596.000 816.320 ;
        RECT 4.400 807.480 596.000 808.880 ;
        RECT 4.000 799.360 596.000 807.480 ;
        RECT 4.400 797.960 596.000 799.360 ;
        RECT 4.000 790.520 596.000 797.960 ;
        RECT 4.400 789.120 596.000 790.520 ;
        RECT 4.000 781.000 596.000 789.120 ;
        RECT 4.400 779.600 596.000 781.000 ;
        RECT 4.000 772.160 596.000 779.600 ;
        RECT 4.400 770.760 596.000 772.160 ;
        RECT 4.000 762.640 596.000 770.760 ;
        RECT 4.400 761.240 596.000 762.640 ;
        RECT 4.000 753.800 596.000 761.240 ;
        RECT 4.400 752.400 596.000 753.800 ;
        RECT 4.000 744.960 596.000 752.400 ;
        RECT 4.400 743.560 596.000 744.960 ;
        RECT 4.000 735.440 596.000 743.560 ;
        RECT 4.400 734.040 596.000 735.440 ;
        RECT 4.000 726.600 596.000 734.040 ;
        RECT 4.400 725.200 596.000 726.600 ;
        RECT 4.000 717.080 596.000 725.200 ;
        RECT 4.400 715.680 596.000 717.080 ;
        RECT 4.000 713.000 596.000 715.680 ;
        RECT 4.000 711.600 595.600 713.000 ;
        RECT 4.000 708.240 596.000 711.600 ;
        RECT 4.400 706.840 596.000 708.240 ;
        RECT 4.000 698.720 596.000 706.840 ;
        RECT 4.400 697.320 596.000 698.720 ;
        RECT 4.000 689.880 596.000 697.320 ;
        RECT 4.400 688.480 596.000 689.880 ;
        RECT 4.000 681.040 596.000 688.480 ;
        RECT 4.400 679.640 596.000 681.040 ;
        RECT 4.000 671.520 596.000 679.640 ;
        RECT 4.400 670.120 596.000 671.520 ;
        RECT 4.000 662.680 596.000 670.120 ;
        RECT 4.400 661.280 596.000 662.680 ;
        RECT 4.000 653.160 596.000 661.280 ;
        RECT 4.400 651.760 596.000 653.160 ;
        RECT 4.000 644.320 596.000 651.760 ;
        RECT 4.400 642.920 596.000 644.320 ;
        RECT 4.000 634.800 596.000 642.920 ;
        RECT 4.400 633.400 596.000 634.800 ;
        RECT 4.000 625.960 596.000 633.400 ;
        RECT 4.400 624.560 596.000 625.960 ;
        RECT 4.000 616.440 596.000 624.560 ;
        RECT 4.400 615.040 596.000 616.440 ;
        RECT 4.000 607.600 596.000 615.040 ;
        RECT 4.400 606.200 596.000 607.600 ;
        RECT 4.000 598.760 596.000 606.200 ;
        RECT 4.400 597.360 596.000 598.760 ;
        RECT 4.000 589.240 596.000 597.360 ;
        RECT 4.400 587.840 596.000 589.240 ;
        RECT 4.000 580.400 596.000 587.840 ;
        RECT 4.400 579.000 596.000 580.400 ;
        RECT 4.000 570.880 596.000 579.000 ;
        RECT 4.400 569.480 596.000 570.880 ;
        RECT 4.000 562.040 596.000 569.480 ;
        RECT 4.400 560.640 596.000 562.040 ;
        RECT 4.000 554.560 596.000 560.640 ;
        RECT 4.000 553.160 595.600 554.560 ;
        RECT 4.000 552.520 596.000 553.160 ;
        RECT 4.400 551.120 596.000 552.520 ;
        RECT 4.000 543.680 596.000 551.120 ;
        RECT 4.400 542.280 596.000 543.680 ;
        RECT 4.000 534.840 596.000 542.280 ;
        RECT 4.400 533.440 596.000 534.840 ;
        RECT 4.000 525.320 596.000 533.440 ;
        RECT 4.400 523.920 596.000 525.320 ;
        RECT 4.000 516.480 596.000 523.920 ;
        RECT 4.400 515.080 596.000 516.480 ;
        RECT 4.000 506.960 596.000 515.080 ;
        RECT 4.400 505.560 596.000 506.960 ;
        RECT 4.000 498.120 596.000 505.560 ;
        RECT 4.400 496.720 596.000 498.120 ;
        RECT 4.000 488.600 596.000 496.720 ;
        RECT 4.400 487.200 596.000 488.600 ;
        RECT 4.000 479.760 596.000 487.200 ;
        RECT 4.400 478.360 596.000 479.760 ;
        RECT 4.000 470.920 596.000 478.360 ;
        RECT 4.400 469.520 596.000 470.920 ;
        RECT 4.000 461.400 596.000 469.520 ;
        RECT 4.400 460.000 596.000 461.400 ;
        RECT 4.000 452.560 596.000 460.000 ;
        RECT 4.400 451.160 596.000 452.560 ;
        RECT 4.000 443.040 596.000 451.160 ;
        RECT 4.400 441.640 596.000 443.040 ;
        RECT 4.000 434.200 596.000 441.640 ;
        RECT 4.400 432.800 596.000 434.200 ;
        RECT 4.000 424.680 596.000 432.800 ;
        RECT 4.400 423.280 596.000 424.680 ;
        RECT 4.000 415.840 596.000 423.280 ;
        RECT 4.400 414.440 596.000 415.840 ;
        RECT 4.000 407.000 596.000 414.440 ;
        RECT 4.400 405.600 596.000 407.000 ;
        RECT 4.000 397.480 596.000 405.600 ;
        RECT 4.400 396.120 596.000 397.480 ;
        RECT 4.400 396.080 595.600 396.120 ;
        RECT 4.000 394.720 595.600 396.080 ;
        RECT 4.000 388.640 596.000 394.720 ;
        RECT 4.400 387.240 596.000 388.640 ;
        RECT 4.000 379.120 596.000 387.240 ;
        RECT 4.400 377.720 596.000 379.120 ;
        RECT 4.000 370.280 596.000 377.720 ;
        RECT 4.400 368.880 596.000 370.280 ;
        RECT 4.000 360.760 596.000 368.880 ;
        RECT 4.400 359.360 596.000 360.760 ;
        RECT 4.000 351.920 596.000 359.360 ;
        RECT 4.400 350.520 596.000 351.920 ;
        RECT 4.000 343.080 596.000 350.520 ;
        RECT 4.400 341.680 596.000 343.080 ;
        RECT 4.000 333.560 596.000 341.680 ;
        RECT 4.400 332.160 596.000 333.560 ;
        RECT 4.000 324.720 596.000 332.160 ;
        RECT 4.400 323.320 596.000 324.720 ;
        RECT 4.000 315.200 596.000 323.320 ;
        RECT 4.400 313.800 596.000 315.200 ;
        RECT 4.000 306.360 596.000 313.800 ;
        RECT 4.400 304.960 596.000 306.360 ;
        RECT 4.000 296.840 596.000 304.960 ;
        RECT 4.400 295.440 596.000 296.840 ;
        RECT 4.000 288.000 596.000 295.440 ;
        RECT 4.400 286.600 596.000 288.000 ;
        RECT 4.000 278.480 596.000 286.600 ;
        RECT 4.400 277.080 596.000 278.480 ;
        RECT 4.000 269.640 596.000 277.080 ;
        RECT 4.400 268.240 596.000 269.640 ;
        RECT 4.000 260.800 596.000 268.240 ;
        RECT 4.400 259.400 596.000 260.800 ;
        RECT 4.000 251.280 596.000 259.400 ;
        RECT 4.400 249.880 596.000 251.280 ;
        RECT 4.000 242.440 596.000 249.880 ;
        RECT 4.400 241.040 596.000 242.440 ;
        RECT 4.000 237.680 596.000 241.040 ;
        RECT 4.000 236.280 595.600 237.680 ;
        RECT 4.000 232.920 596.000 236.280 ;
        RECT 4.400 231.520 596.000 232.920 ;
        RECT 4.000 224.080 596.000 231.520 ;
        RECT 4.400 222.680 596.000 224.080 ;
        RECT 4.000 214.560 596.000 222.680 ;
        RECT 4.400 213.160 596.000 214.560 ;
        RECT 4.000 205.720 596.000 213.160 ;
        RECT 4.400 204.320 596.000 205.720 ;
        RECT 4.000 196.880 596.000 204.320 ;
        RECT 4.400 195.480 596.000 196.880 ;
        RECT 4.000 187.360 596.000 195.480 ;
        RECT 4.400 185.960 596.000 187.360 ;
        RECT 4.000 178.520 596.000 185.960 ;
        RECT 4.400 177.120 596.000 178.520 ;
        RECT 4.000 169.000 596.000 177.120 ;
        RECT 4.400 167.600 596.000 169.000 ;
        RECT 4.000 160.160 596.000 167.600 ;
        RECT 4.400 158.760 596.000 160.160 ;
        RECT 4.000 150.640 596.000 158.760 ;
        RECT 4.400 149.240 596.000 150.640 ;
        RECT 4.000 141.800 596.000 149.240 ;
        RECT 4.400 140.400 596.000 141.800 ;
        RECT 4.000 132.960 596.000 140.400 ;
        RECT 4.400 131.560 596.000 132.960 ;
        RECT 4.000 123.440 596.000 131.560 ;
        RECT 4.400 122.040 596.000 123.440 ;
        RECT 4.000 114.600 596.000 122.040 ;
        RECT 4.400 113.200 596.000 114.600 ;
        RECT 4.000 105.080 596.000 113.200 ;
        RECT 4.400 103.680 596.000 105.080 ;
        RECT 4.000 96.240 596.000 103.680 ;
        RECT 4.400 94.840 596.000 96.240 ;
        RECT 4.000 86.720 596.000 94.840 ;
        RECT 4.400 85.320 596.000 86.720 ;
        RECT 4.000 79.920 596.000 85.320 ;
        RECT 4.000 78.520 595.600 79.920 ;
        RECT 4.000 77.880 596.000 78.520 ;
        RECT 4.400 76.480 596.000 77.880 ;
        RECT 4.000 69.040 596.000 76.480 ;
        RECT 4.400 67.640 596.000 69.040 ;
        RECT 4.000 59.520 596.000 67.640 ;
        RECT 4.400 58.120 596.000 59.520 ;
        RECT 4.000 50.680 596.000 58.120 ;
        RECT 4.400 49.280 596.000 50.680 ;
        RECT 4.000 41.160 596.000 49.280 ;
        RECT 4.400 39.760 596.000 41.160 ;
        RECT 4.000 32.320 596.000 39.760 ;
        RECT 4.400 30.920 596.000 32.320 ;
        RECT 4.000 22.800 596.000 30.920 ;
        RECT 4.400 21.400 596.000 22.800 ;
        RECT 4.000 13.960 596.000 21.400 ;
        RECT 4.400 12.560 596.000 13.960 ;
        RECT 4.000 5.120 596.000 12.560 ;
        RECT 4.400 4.255 596.000 5.120 ;
      LAYER met4 ;
        RECT 9.495 13.095 20.640 934.145 ;
        RECT 23.040 13.095 97.440 934.145 ;
        RECT 99.840 13.095 174.240 934.145 ;
        RECT 176.640 13.095 251.040 934.145 ;
        RECT 253.440 13.095 327.840 934.145 ;
        RECT 330.240 13.095 404.640 934.145 ;
        RECT 407.040 13.095 481.440 934.145 ;
        RECT 483.840 13.095 558.240 934.145 ;
        RECT 560.640 13.095 580.225 934.145 ;
  END
END Peripherals
END LIBRARY

