magic
tech sky130A
magscale 1 2
timestamp 1652729090
<< nwell >>
rect 1066 97093 38862 97414
rect 1066 96005 38862 96571
rect 1066 94917 38862 95483
rect 1066 93829 38862 94395
rect 1066 92741 38862 93307
rect 1066 91653 38862 92219
rect 1066 90565 38862 91131
rect 1066 89477 38862 90043
rect 1066 88389 38862 88955
rect 1066 87301 38862 87867
rect 1066 86213 38862 86779
rect 1066 85125 38862 85691
rect 1066 84037 38862 84603
rect 1066 82949 38862 83515
rect 1066 81861 38862 82427
rect 1066 80773 38862 81339
rect 1066 79685 38862 80251
rect 1066 78597 38862 79163
rect 1066 77509 38862 78075
rect 1066 76421 38862 76987
rect 1066 75333 38862 75899
rect 1066 74245 38862 74811
rect 1066 73157 38862 73723
rect 1066 72069 38862 72635
rect 1066 70981 38862 71547
rect 1066 69893 38862 70459
rect 1066 68805 38862 69371
rect 1066 67717 38862 68283
rect 1066 66629 38862 67195
rect 1066 65541 38862 66107
rect 1066 64453 38862 65019
rect 1066 63365 38862 63931
rect 1066 62277 38862 62843
rect 1066 61189 38862 61755
rect 1066 60101 38862 60667
rect 1066 59013 38862 59579
rect 1066 57925 38862 58491
rect 1066 56837 38862 57403
rect 1066 55749 38862 56315
rect 1066 54661 38862 55227
rect 1066 53573 38862 54139
rect 1066 52485 38862 53051
rect 1066 51397 38862 51963
rect 1066 50309 38862 50875
rect 1066 49221 38862 49787
rect 1066 48133 38862 48699
rect 1066 47045 38862 47611
rect 1066 45957 38862 46523
rect 1066 44869 38862 45435
rect 1066 43781 38862 44347
rect 1066 42693 38862 43259
rect 1066 41605 38862 42171
rect 1066 40517 38862 41083
rect 1066 39429 38862 39995
rect 1066 38341 38862 38907
rect 1066 37253 38862 37819
rect 1066 36165 38862 36731
rect 1066 35077 38862 35643
rect 1066 33989 38862 34555
rect 1066 32901 38862 33467
rect 1066 31813 38862 32379
rect 1066 30725 38862 31291
rect 1066 29637 38862 30203
rect 1066 28549 38862 29115
rect 1066 27461 38862 28027
rect 1066 26373 38862 26939
rect 1066 25285 38862 25851
rect 1066 24197 38862 24763
rect 1066 23109 38862 23675
rect 1066 22021 38862 22587
rect 1066 20933 38862 21499
rect 1066 19845 38862 20411
rect 1066 18757 38862 19323
rect 1066 17669 38862 18235
rect 1066 16581 38862 17147
rect 1066 15493 38862 16059
rect 1066 14405 38862 14971
rect 1066 13317 38862 13883
rect 1066 12229 38862 12795
rect 1066 11141 38862 11707
rect 1066 10053 38862 10619
rect 1066 8965 38862 9531
rect 1066 7877 38862 8443
rect 1066 6789 38862 7355
rect 1066 5701 38862 6267
rect 1066 4613 38862 5179
rect 1066 3525 38862 4091
rect 1066 2437 38862 3003
<< obsli1 >>
rect 1104 2159 38824 97393
<< obsm1 >>
rect 1104 2128 38824 97424
<< metal2 >>
rect 2502 99200 2558 100000
rect 7470 99200 7526 100000
rect 12438 99200 12494 100000
rect 17498 99200 17554 100000
rect 22466 99200 22522 100000
rect 27434 99200 27490 100000
rect 32494 99200 32550 100000
rect 37462 99200 37518 100000
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 2614 99144 7414 99362
rect 7582 99144 12382 99362
rect 12550 99144 17442 99362
rect 17610 99144 22410 99362
rect 22578 99144 27378 99362
rect 27546 99144 32438 99362
rect 32606 99144 37406 99362
rect 37574 99144 38162 99362
rect 2558 856 38162 99144
rect 2558 439 9898 856
rect 10066 439 29862 856
rect 30030 439 38162 856
<< metal3 >>
rect 39200 99288 40000 99408
rect 39200 98336 40000 98456
rect 39200 97248 40000 97368
rect 39200 96296 40000 96416
rect 39200 95208 40000 95328
rect 39200 94256 40000 94376
rect 39200 93304 40000 93424
rect 39200 92216 40000 92336
rect 39200 91264 40000 91384
rect 39200 90176 40000 90296
rect 39200 89224 40000 89344
rect 39200 88136 40000 88256
rect 39200 87184 40000 87304
rect 39200 86232 40000 86352
rect 39200 85144 40000 85264
rect 39200 84192 40000 84312
rect 39200 83104 40000 83224
rect 39200 82152 40000 82272
rect 39200 81064 40000 81184
rect 39200 80112 40000 80232
rect 39200 79160 40000 79280
rect 39200 78072 40000 78192
rect 39200 77120 40000 77240
rect 39200 76032 40000 76152
rect 39200 75080 40000 75200
rect 39200 73992 40000 74112
rect 39200 73040 40000 73160
rect 39200 72088 40000 72208
rect 39200 71000 40000 71120
rect 39200 70048 40000 70168
rect 39200 68960 40000 69080
rect 39200 68008 40000 68128
rect 39200 67056 40000 67176
rect 39200 65968 40000 66088
rect 39200 65016 40000 65136
rect 39200 63928 40000 64048
rect 39200 62976 40000 63096
rect 39200 61888 40000 62008
rect 39200 60936 40000 61056
rect 39200 59984 40000 60104
rect 39200 58896 40000 59016
rect 39200 57944 40000 58064
rect 39200 56856 40000 56976
rect 39200 55904 40000 56024
rect 39200 54816 40000 54936
rect 39200 53864 40000 53984
rect 39200 52912 40000 53032
rect 39200 51824 40000 51944
rect 39200 50872 40000 50992
rect 39200 49784 40000 49904
rect 39200 48832 40000 48952
rect 39200 47744 40000 47864
rect 39200 46792 40000 46912
rect 39200 45840 40000 45960
rect 39200 44752 40000 44872
rect 39200 43800 40000 43920
rect 39200 42712 40000 42832
rect 39200 41760 40000 41880
rect 39200 40672 40000 40792
rect 39200 39720 40000 39840
rect 39200 38768 40000 38888
rect 39200 37680 40000 37800
rect 39200 36728 40000 36848
rect 39200 35640 40000 35760
rect 39200 34688 40000 34808
rect 39200 33736 40000 33856
rect 39200 32648 40000 32768
rect 39200 31696 40000 31816
rect 39200 30608 40000 30728
rect 39200 29656 40000 29776
rect 39200 28568 40000 28688
rect 39200 27616 40000 27736
rect 39200 26664 40000 26784
rect 39200 25576 40000 25696
rect 39200 24624 40000 24744
rect 39200 23536 40000 23656
rect 39200 22584 40000 22704
rect 39200 21496 40000 21616
rect 39200 20544 40000 20664
rect 39200 19592 40000 19712
rect 39200 18504 40000 18624
rect 39200 17552 40000 17672
rect 39200 16464 40000 16584
rect 39200 15512 40000 15632
rect 39200 14424 40000 14544
rect 39200 13472 40000 13592
rect 39200 12520 40000 12640
rect 39200 11432 40000 11552
rect 39200 10480 40000 10600
rect 39200 9392 40000 9512
rect 39200 8440 40000 8560
rect 39200 7352 40000 7472
rect 39200 6400 40000 6520
rect 39200 5448 40000 5568
rect 39200 4360 40000 4480
rect 39200 3408 40000 3528
rect 39200 2320 40000 2440
rect 39200 1368 40000 1488
rect 39200 416 40000 536
<< obsm3 >>
rect 4208 98256 39120 98429
rect 4208 97448 39200 98256
rect 4208 97168 39120 97448
rect 4208 96496 39200 97168
rect 4208 96216 39120 96496
rect 4208 95408 39200 96216
rect 4208 95128 39120 95408
rect 4208 94456 39200 95128
rect 4208 94176 39120 94456
rect 4208 93504 39200 94176
rect 4208 93224 39120 93504
rect 4208 92416 39200 93224
rect 4208 92136 39120 92416
rect 4208 91464 39200 92136
rect 4208 91184 39120 91464
rect 4208 90376 39200 91184
rect 4208 90096 39120 90376
rect 4208 89424 39200 90096
rect 4208 89144 39120 89424
rect 4208 88336 39200 89144
rect 4208 88056 39120 88336
rect 4208 87384 39200 88056
rect 4208 87104 39120 87384
rect 4208 86432 39200 87104
rect 4208 86152 39120 86432
rect 4208 85344 39200 86152
rect 4208 85064 39120 85344
rect 4208 84392 39200 85064
rect 4208 84112 39120 84392
rect 4208 83304 39200 84112
rect 4208 83024 39120 83304
rect 4208 82352 39200 83024
rect 4208 82072 39120 82352
rect 4208 81264 39200 82072
rect 4208 80984 39120 81264
rect 4208 80312 39200 80984
rect 4208 80032 39120 80312
rect 4208 79360 39200 80032
rect 4208 79080 39120 79360
rect 4208 78272 39200 79080
rect 4208 77992 39120 78272
rect 4208 77320 39200 77992
rect 4208 77040 39120 77320
rect 4208 76232 39200 77040
rect 4208 75952 39120 76232
rect 4208 75280 39200 75952
rect 4208 75000 39120 75280
rect 4208 74192 39200 75000
rect 4208 73912 39120 74192
rect 4208 73240 39200 73912
rect 4208 72960 39120 73240
rect 4208 72288 39200 72960
rect 4208 72008 39120 72288
rect 4208 71200 39200 72008
rect 4208 70920 39120 71200
rect 4208 70248 39200 70920
rect 4208 69968 39120 70248
rect 4208 69160 39200 69968
rect 4208 68880 39120 69160
rect 4208 68208 39200 68880
rect 4208 67928 39120 68208
rect 4208 67256 39200 67928
rect 4208 66976 39120 67256
rect 4208 66168 39200 66976
rect 4208 65888 39120 66168
rect 4208 65216 39200 65888
rect 4208 64936 39120 65216
rect 4208 64128 39200 64936
rect 4208 63848 39120 64128
rect 4208 63176 39200 63848
rect 4208 62896 39120 63176
rect 4208 62088 39200 62896
rect 4208 61808 39120 62088
rect 4208 61136 39200 61808
rect 4208 60856 39120 61136
rect 4208 60184 39200 60856
rect 4208 59904 39120 60184
rect 4208 59096 39200 59904
rect 4208 58816 39120 59096
rect 4208 58144 39200 58816
rect 4208 57864 39120 58144
rect 4208 57056 39200 57864
rect 4208 56776 39120 57056
rect 4208 56104 39200 56776
rect 4208 55824 39120 56104
rect 4208 55016 39200 55824
rect 4208 54736 39120 55016
rect 4208 54064 39200 54736
rect 4208 53784 39120 54064
rect 4208 53112 39200 53784
rect 4208 52832 39120 53112
rect 4208 52024 39200 52832
rect 4208 51744 39120 52024
rect 4208 51072 39200 51744
rect 4208 50792 39120 51072
rect 4208 49984 39200 50792
rect 4208 49704 39120 49984
rect 4208 49032 39200 49704
rect 4208 48752 39120 49032
rect 4208 47944 39200 48752
rect 4208 47664 39120 47944
rect 4208 46992 39200 47664
rect 4208 46712 39120 46992
rect 4208 46040 39200 46712
rect 4208 45760 39120 46040
rect 4208 44952 39200 45760
rect 4208 44672 39120 44952
rect 4208 44000 39200 44672
rect 4208 43720 39120 44000
rect 4208 42912 39200 43720
rect 4208 42632 39120 42912
rect 4208 41960 39200 42632
rect 4208 41680 39120 41960
rect 4208 40872 39200 41680
rect 4208 40592 39120 40872
rect 4208 39920 39200 40592
rect 4208 39640 39120 39920
rect 4208 38968 39200 39640
rect 4208 38688 39120 38968
rect 4208 37880 39200 38688
rect 4208 37600 39120 37880
rect 4208 36928 39200 37600
rect 4208 36648 39120 36928
rect 4208 35840 39200 36648
rect 4208 35560 39120 35840
rect 4208 34888 39200 35560
rect 4208 34608 39120 34888
rect 4208 33936 39200 34608
rect 4208 33656 39120 33936
rect 4208 32848 39200 33656
rect 4208 32568 39120 32848
rect 4208 31896 39200 32568
rect 4208 31616 39120 31896
rect 4208 30808 39200 31616
rect 4208 30528 39120 30808
rect 4208 29856 39200 30528
rect 4208 29576 39120 29856
rect 4208 28768 39200 29576
rect 4208 28488 39120 28768
rect 4208 27816 39200 28488
rect 4208 27536 39120 27816
rect 4208 26864 39200 27536
rect 4208 26584 39120 26864
rect 4208 25776 39200 26584
rect 4208 25496 39120 25776
rect 4208 24824 39200 25496
rect 4208 24544 39120 24824
rect 4208 23736 39200 24544
rect 4208 23456 39120 23736
rect 4208 22784 39200 23456
rect 4208 22504 39120 22784
rect 4208 21696 39200 22504
rect 4208 21416 39120 21696
rect 4208 20744 39200 21416
rect 4208 20464 39120 20744
rect 4208 19792 39200 20464
rect 4208 19512 39120 19792
rect 4208 18704 39200 19512
rect 4208 18424 39120 18704
rect 4208 17752 39200 18424
rect 4208 17472 39120 17752
rect 4208 16664 39200 17472
rect 4208 16384 39120 16664
rect 4208 15712 39200 16384
rect 4208 15432 39120 15712
rect 4208 14624 39200 15432
rect 4208 14344 39120 14624
rect 4208 13672 39200 14344
rect 4208 13392 39120 13672
rect 4208 12720 39200 13392
rect 4208 12440 39120 12720
rect 4208 11632 39200 12440
rect 4208 11352 39120 11632
rect 4208 10680 39200 11352
rect 4208 10400 39120 10680
rect 4208 9592 39200 10400
rect 4208 9312 39120 9592
rect 4208 8640 39200 9312
rect 4208 8360 39120 8640
rect 4208 7552 39200 8360
rect 4208 7272 39120 7552
rect 4208 6600 39200 7272
rect 4208 6320 39120 6600
rect 4208 5648 39200 6320
rect 4208 5368 39120 5648
rect 4208 4560 39200 5368
rect 4208 4280 39120 4560
rect 4208 3608 39200 4280
rect 4208 3328 39120 3608
rect 4208 2520 39200 3328
rect 4208 2240 39120 2520
rect 4208 1568 39200 2240
rect 4208 1288 39120 1568
rect 4208 616 39200 1288
rect 4208 443 39120 616
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
<< labels >>
rlabel metal2 s 9954 0 10010 800 6 clk
port 1 nsew signal input
rlabel metal3 s 39200 3408 40000 3528 6 core0Address[0]
port 2 nsew signal input
rlabel metal3 s 39200 37680 40000 37800 6 core0Address[10]
port 3 nsew signal input
rlabel metal3 s 39200 40672 40000 40792 6 core0Address[11]
port 4 nsew signal input
rlabel metal3 s 39200 43800 40000 43920 6 core0Address[12]
port 5 nsew signal input
rlabel metal3 s 39200 46792 40000 46912 6 core0Address[13]
port 6 nsew signal input
rlabel metal3 s 39200 49784 40000 49904 6 core0Address[14]
port 7 nsew signal input
rlabel metal3 s 39200 52912 40000 53032 6 core0Address[15]
port 8 nsew signal input
rlabel metal3 s 39200 55904 40000 56024 6 core0Address[16]
port 9 nsew signal input
rlabel metal3 s 39200 58896 40000 59016 6 core0Address[17]
port 10 nsew signal input
rlabel metal3 s 39200 61888 40000 62008 6 core0Address[18]
port 11 nsew signal input
rlabel metal3 s 39200 65016 40000 65136 6 core0Address[19]
port 12 nsew signal input
rlabel metal3 s 39200 7352 40000 7472 6 core0Address[1]
port 13 nsew signal input
rlabel metal3 s 39200 68008 40000 68128 6 core0Address[20]
port 14 nsew signal input
rlabel metal3 s 39200 71000 40000 71120 6 core0Address[21]
port 15 nsew signal input
rlabel metal3 s 39200 73992 40000 74112 6 core0Address[22]
port 16 nsew signal input
rlabel metal3 s 39200 77120 40000 77240 6 core0Address[23]
port 17 nsew signal input
rlabel metal3 s 39200 80112 40000 80232 6 core0Address[24]
port 18 nsew signal input
rlabel metal3 s 39200 83104 40000 83224 6 core0Address[25]
port 19 nsew signal input
rlabel metal3 s 39200 86232 40000 86352 6 core0Address[26]
port 20 nsew signal input
rlabel metal3 s 39200 89224 40000 89344 6 core0Address[27]
port 21 nsew signal input
rlabel metal3 s 39200 11432 40000 11552 6 core0Address[2]
port 22 nsew signal input
rlabel metal3 s 39200 15512 40000 15632 6 core0Address[3]
port 23 nsew signal input
rlabel metal3 s 39200 19592 40000 19712 6 core0Address[4]
port 24 nsew signal input
rlabel metal3 s 39200 22584 40000 22704 6 core0Address[5]
port 25 nsew signal input
rlabel metal3 s 39200 25576 40000 25696 6 core0Address[6]
port 26 nsew signal input
rlabel metal3 s 39200 28568 40000 28688 6 core0Address[7]
port 27 nsew signal input
rlabel metal3 s 39200 31696 40000 31816 6 core0Address[8]
port 28 nsew signal input
rlabel metal3 s 39200 34688 40000 34808 6 core0Address[9]
port 29 nsew signal input
rlabel metal3 s 39200 416 40000 536 6 core0Busy
port 30 nsew signal output
rlabel metal3 s 39200 4360 40000 4480 6 core0ByteSelect[0]
port 31 nsew signal input
rlabel metal3 s 39200 8440 40000 8560 6 core0ByteSelect[1]
port 32 nsew signal input
rlabel metal3 s 39200 12520 40000 12640 6 core0ByteSelect[2]
port 33 nsew signal input
rlabel metal3 s 39200 16464 40000 16584 6 core0ByteSelect[3]
port 34 nsew signal input
rlabel metal3 s 39200 5448 40000 5568 6 core0DataRead[0]
port 35 nsew signal output
rlabel metal3 s 39200 38768 40000 38888 6 core0DataRead[10]
port 36 nsew signal output
rlabel metal3 s 39200 41760 40000 41880 6 core0DataRead[11]
port 37 nsew signal output
rlabel metal3 s 39200 44752 40000 44872 6 core0DataRead[12]
port 38 nsew signal output
rlabel metal3 s 39200 47744 40000 47864 6 core0DataRead[13]
port 39 nsew signal output
rlabel metal3 s 39200 50872 40000 50992 6 core0DataRead[14]
port 40 nsew signal output
rlabel metal3 s 39200 53864 40000 53984 6 core0DataRead[15]
port 41 nsew signal output
rlabel metal3 s 39200 56856 40000 56976 6 core0DataRead[16]
port 42 nsew signal output
rlabel metal3 s 39200 59984 40000 60104 6 core0DataRead[17]
port 43 nsew signal output
rlabel metal3 s 39200 62976 40000 63096 6 core0DataRead[18]
port 44 nsew signal output
rlabel metal3 s 39200 65968 40000 66088 6 core0DataRead[19]
port 45 nsew signal output
rlabel metal3 s 39200 9392 40000 9512 6 core0DataRead[1]
port 46 nsew signal output
rlabel metal3 s 39200 68960 40000 69080 6 core0DataRead[20]
port 47 nsew signal output
rlabel metal3 s 39200 72088 40000 72208 6 core0DataRead[21]
port 48 nsew signal output
rlabel metal3 s 39200 75080 40000 75200 6 core0DataRead[22]
port 49 nsew signal output
rlabel metal3 s 39200 78072 40000 78192 6 core0DataRead[23]
port 50 nsew signal output
rlabel metal3 s 39200 81064 40000 81184 6 core0DataRead[24]
port 51 nsew signal output
rlabel metal3 s 39200 84192 40000 84312 6 core0DataRead[25]
port 52 nsew signal output
rlabel metal3 s 39200 87184 40000 87304 6 core0DataRead[26]
port 53 nsew signal output
rlabel metal3 s 39200 90176 40000 90296 6 core0DataRead[27]
port 54 nsew signal output
rlabel metal3 s 39200 92216 40000 92336 6 core0DataRead[28]
port 55 nsew signal output
rlabel metal3 s 39200 94256 40000 94376 6 core0DataRead[29]
port 56 nsew signal output
rlabel metal3 s 39200 13472 40000 13592 6 core0DataRead[2]
port 57 nsew signal output
rlabel metal3 s 39200 96296 40000 96416 6 core0DataRead[30]
port 58 nsew signal output
rlabel metal3 s 39200 98336 40000 98456 6 core0DataRead[31]
port 59 nsew signal output
rlabel metal3 s 39200 17552 40000 17672 6 core0DataRead[3]
port 60 nsew signal output
rlabel metal3 s 39200 20544 40000 20664 6 core0DataRead[4]
port 61 nsew signal output
rlabel metal3 s 39200 23536 40000 23656 6 core0DataRead[5]
port 62 nsew signal output
rlabel metal3 s 39200 26664 40000 26784 6 core0DataRead[6]
port 63 nsew signal output
rlabel metal3 s 39200 29656 40000 29776 6 core0DataRead[7]
port 64 nsew signal output
rlabel metal3 s 39200 32648 40000 32768 6 core0DataRead[8]
port 65 nsew signal output
rlabel metal3 s 39200 35640 40000 35760 6 core0DataRead[9]
port 66 nsew signal output
rlabel metal3 s 39200 6400 40000 6520 6 core0DataWrite[0]
port 67 nsew signal input
rlabel metal3 s 39200 39720 40000 39840 6 core0DataWrite[10]
port 68 nsew signal input
rlabel metal3 s 39200 42712 40000 42832 6 core0DataWrite[11]
port 69 nsew signal input
rlabel metal3 s 39200 45840 40000 45960 6 core0DataWrite[12]
port 70 nsew signal input
rlabel metal3 s 39200 48832 40000 48952 6 core0DataWrite[13]
port 71 nsew signal input
rlabel metal3 s 39200 51824 40000 51944 6 core0DataWrite[14]
port 72 nsew signal input
rlabel metal3 s 39200 54816 40000 54936 6 core0DataWrite[15]
port 73 nsew signal input
rlabel metal3 s 39200 57944 40000 58064 6 core0DataWrite[16]
port 74 nsew signal input
rlabel metal3 s 39200 60936 40000 61056 6 core0DataWrite[17]
port 75 nsew signal input
rlabel metal3 s 39200 63928 40000 64048 6 core0DataWrite[18]
port 76 nsew signal input
rlabel metal3 s 39200 67056 40000 67176 6 core0DataWrite[19]
port 77 nsew signal input
rlabel metal3 s 39200 10480 40000 10600 6 core0DataWrite[1]
port 78 nsew signal input
rlabel metal3 s 39200 70048 40000 70168 6 core0DataWrite[20]
port 79 nsew signal input
rlabel metal3 s 39200 73040 40000 73160 6 core0DataWrite[21]
port 80 nsew signal input
rlabel metal3 s 39200 76032 40000 76152 6 core0DataWrite[22]
port 81 nsew signal input
rlabel metal3 s 39200 79160 40000 79280 6 core0DataWrite[23]
port 82 nsew signal input
rlabel metal3 s 39200 82152 40000 82272 6 core0DataWrite[24]
port 83 nsew signal input
rlabel metal3 s 39200 85144 40000 85264 6 core0DataWrite[25]
port 84 nsew signal input
rlabel metal3 s 39200 88136 40000 88256 6 core0DataWrite[26]
port 85 nsew signal input
rlabel metal3 s 39200 91264 40000 91384 6 core0DataWrite[27]
port 86 nsew signal input
rlabel metal3 s 39200 93304 40000 93424 6 core0DataWrite[28]
port 87 nsew signal input
rlabel metal3 s 39200 95208 40000 95328 6 core0DataWrite[29]
port 88 nsew signal input
rlabel metal3 s 39200 14424 40000 14544 6 core0DataWrite[2]
port 89 nsew signal input
rlabel metal3 s 39200 97248 40000 97368 6 core0DataWrite[30]
port 90 nsew signal input
rlabel metal3 s 39200 99288 40000 99408 6 core0DataWrite[31]
port 91 nsew signal input
rlabel metal3 s 39200 18504 40000 18624 6 core0DataWrite[3]
port 92 nsew signal input
rlabel metal3 s 39200 21496 40000 21616 6 core0DataWrite[4]
port 93 nsew signal input
rlabel metal3 s 39200 24624 40000 24744 6 core0DataWrite[5]
port 94 nsew signal input
rlabel metal3 s 39200 27616 40000 27736 6 core0DataWrite[6]
port 95 nsew signal input
rlabel metal3 s 39200 30608 40000 30728 6 core0DataWrite[7]
port 96 nsew signal input
rlabel metal3 s 39200 33736 40000 33856 6 core0DataWrite[8]
port 97 nsew signal input
rlabel metal3 s 39200 36728 40000 36848 6 core0DataWrite[9]
port 98 nsew signal input
rlabel metal3 s 39200 1368 40000 1488 6 core0ReadEnable
port 99 nsew signal input
rlabel metal3 s 39200 2320 40000 2440 6 core0WriteEnable
port 100 nsew signal input
rlabel metal2 s 2502 99200 2558 100000 6 flash_csb
port 101 nsew signal output
rlabel metal2 s 7470 99200 7526 100000 6 flash_io0_read
port 102 nsew signal input
rlabel metal2 s 12438 99200 12494 100000 6 flash_io0_we
port 103 nsew signal output
rlabel metal2 s 17498 99200 17554 100000 6 flash_io0_write
port 104 nsew signal output
rlabel metal2 s 22466 99200 22522 100000 6 flash_io1_read
port 105 nsew signal input
rlabel metal2 s 27434 99200 27490 100000 6 flash_io1_we
port 106 nsew signal output
rlabel metal2 s 32494 99200 32550 100000 6 flash_io1_write
port 107 nsew signal output
rlabel metal2 s 37462 99200 37518 100000 6 flash_sck
port 108 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 rst
port 109 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 110 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 110 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 111 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1072144
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Flash/runs/Flash/results/finishing/Flash.magic.gds
string GDS_START 24096
<< end >>

