VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WBPeripheralBusInterface
  CLASS BLOCK ;
  FOREIGN WBPeripheralBusInterface ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN peripheralBus_address[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 200.000 7.440 ;
    END
  END peripheralBus_address[0]
  PIN peripheralBus_address[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.240 200.000 78.840 ;
    END
  END peripheralBus_address[10]
  PIN peripheralBus_address[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 84.360 200.000 84.960 ;
    END
  END peripheralBus_address[11]
  PIN peripheralBus_address[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 91.160 200.000 91.760 ;
    END
  END peripheralBus_address[12]
  PIN peripheralBus_address[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 97.280 200.000 97.880 ;
    END
  END peripheralBus_address[13]
  PIN peripheralBus_address[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 103.400 200.000 104.000 ;
    END
  END peripheralBus_address[14]
  PIN peripheralBus_address[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 109.520 200.000 110.120 ;
    END
  END peripheralBus_address[15]
  PIN peripheralBus_address[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 116.320 200.000 116.920 ;
    END
  END peripheralBus_address[16]
  PIN peripheralBus_address[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 122.440 200.000 123.040 ;
    END
  END peripheralBus_address[17]
  PIN peripheralBus_address[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 128.560 200.000 129.160 ;
    END
  END peripheralBus_address[18]
  PIN peripheralBus_address[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 135.360 200.000 135.960 ;
    END
  END peripheralBus_address[19]
  PIN peripheralBus_address[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 15.000 200.000 15.600 ;
    END
  END peripheralBus_address[1]
  PIN peripheralBus_address[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 141.480 200.000 142.080 ;
    END
  END peripheralBus_address[20]
  PIN peripheralBus_address[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 147.600 200.000 148.200 ;
    END
  END peripheralBus_address[21]
  PIN peripheralBus_address[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 153.720 200.000 154.320 ;
    END
  END peripheralBus_address[22]
  PIN peripheralBus_address[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 160.520 200.000 161.120 ;
    END
  END peripheralBus_address[23]
  PIN peripheralBus_address[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.840 200.000 24.440 ;
    END
  END peripheralBus_address[2]
  PIN peripheralBus_address[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 32.000 200.000 32.600 ;
    END
  END peripheralBus_address[3]
  PIN peripheralBus_address[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 40.160 200.000 40.760 ;
    END
  END peripheralBus_address[4]
  PIN peripheralBus_address[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 46.960 200.000 47.560 ;
    END
  END peripheralBus_address[5]
  PIN peripheralBus_address[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 53.080 200.000 53.680 ;
    END
  END peripheralBus_address[6]
  PIN peripheralBus_address[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 59.200 200.000 59.800 ;
    END
  END peripheralBus_address[7]
  PIN peripheralBus_address[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 65.320 200.000 65.920 ;
    END
  END peripheralBus_address[8]
  PIN peripheralBus_address[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 72.120 200.000 72.720 ;
    END
  END peripheralBus_address[9]
  PIN peripheralBus_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 0.720 200.000 1.320 ;
    END
  END peripheralBus_busy
  PIN peripheralBus_byteSelect[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 8.880 200.000 9.480 ;
    END
  END peripheralBus_byteSelect[0]
  PIN peripheralBus_byteSelect[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 17.040 200.000 17.640 ;
    END
  END peripheralBus_byteSelect[1]
  PIN peripheralBus_byteSelect[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 25.880 200.000 26.480 ;
    END
  END peripheralBus_byteSelect[2]
  PIN peripheralBus_byteSelect[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.040 200.000 34.640 ;
    END
  END peripheralBus_byteSelect[3]
  PIN peripheralBus_dataRead[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 10.920 200.000 11.520 ;
    END
  END peripheralBus_dataRead[0]
  PIN peripheralBus_dataRead[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 80.280 200.000 80.880 ;
    END
  END peripheralBus_dataRead[10]
  PIN peripheralBus_dataRead[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 86.400 200.000 87.000 ;
    END
  END peripheralBus_dataRead[11]
  PIN peripheralBus_dataRead[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 93.200 200.000 93.800 ;
    END
  END peripheralBus_dataRead[12]
  PIN peripheralBus_dataRead[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 99.320 200.000 99.920 ;
    END
  END peripheralBus_dataRead[13]
  PIN peripheralBus_dataRead[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 105.440 200.000 106.040 ;
    END
  END peripheralBus_dataRead[14]
  PIN peripheralBus_dataRead[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 200.000 112.840 ;
    END
  END peripheralBus_dataRead[15]
  PIN peripheralBus_dataRead[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 118.360 200.000 118.960 ;
    END
  END peripheralBus_dataRead[16]
  PIN peripheralBus_dataRead[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 124.480 200.000 125.080 ;
    END
  END peripheralBus_dataRead[17]
  PIN peripheralBus_dataRead[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 130.600 200.000 131.200 ;
    END
  END peripheralBus_dataRead[18]
  PIN peripheralBus_dataRead[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 137.400 200.000 138.000 ;
    END
  END peripheralBus_dataRead[19]
  PIN peripheralBus_dataRead[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 19.080 200.000 19.680 ;
    END
  END peripheralBus_dataRead[1]
  PIN peripheralBus_dataRead[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 143.520 200.000 144.120 ;
    END
  END peripheralBus_dataRead[20]
  PIN peripheralBus_dataRead[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 149.640 200.000 150.240 ;
    END
  END peripheralBus_dataRead[21]
  PIN peripheralBus_dataRead[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 156.440 200.000 157.040 ;
    END
  END peripheralBus_dataRead[22]
  PIN peripheralBus_dataRead[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 162.560 200.000 163.160 ;
    END
  END peripheralBus_dataRead[23]
  PIN peripheralBus_dataRead[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 166.640 200.000 167.240 ;
    END
  END peripheralBus_dataRead[24]
  PIN peripheralBus_dataRead[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.720 200.000 171.320 ;
    END
  END peripheralBus_dataRead[25]
  PIN peripheralBus_dataRead[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 174.800 200.000 175.400 ;
    END
  END peripheralBus_dataRead[26]
  PIN peripheralBus_dataRead[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 179.560 200.000 180.160 ;
    END
  END peripheralBus_dataRead[27]
  PIN peripheralBus_dataRead[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 183.640 200.000 184.240 ;
    END
  END peripheralBus_dataRead[28]
  PIN peripheralBus_dataRead[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.720 200.000 188.320 ;
    END
  END peripheralBus_dataRead[29]
  PIN peripheralBus_dataRead[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 27.920 200.000 28.520 ;
    END
  END peripheralBus_dataRead[2]
  PIN peripheralBus_dataRead[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 191.800 200.000 192.400 ;
    END
  END peripheralBus_dataRead[30]
  PIN peripheralBus_dataRead[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 195.880 200.000 196.480 ;
    END
  END peripheralBus_dataRead[31]
  PIN peripheralBus_dataRead[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 36.080 200.000 36.680 ;
    END
  END peripheralBus_dataRead[3]
  PIN peripheralBus_dataRead[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 42.200 200.000 42.800 ;
    END
  END peripheralBus_dataRead[4]
  PIN peripheralBus_dataRead[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 49.000 200.000 49.600 ;
    END
  END peripheralBus_dataRead[5]
  PIN peripheralBus_dataRead[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 55.120 200.000 55.720 ;
    END
  END peripheralBus_dataRead[6]
  PIN peripheralBus_dataRead[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END peripheralBus_dataRead[7]
  PIN peripheralBus_dataRead[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 68.040 200.000 68.640 ;
    END
  END peripheralBus_dataRead[8]
  PIN peripheralBus_dataRead[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.160 200.000 74.760 ;
    END
  END peripheralBus_dataRead[9]
  PIN peripheralBus_dataWrite[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 12.960 200.000 13.560 ;
    END
  END peripheralBus_dataWrite[0]
  PIN peripheralBus_dataWrite[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 82.320 200.000 82.920 ;
    END
  END peripheralBus_dataWrite[10]
  PIN peripheralBus_dataWrite[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 200.000 89.040 ;
    END
  END peripheralBus_dataWrite[11]
  PIN peripheralBus_dataWrite[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END peripheralBus_dataWrite[12]
  PIN peripheralBus_dataWrite[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 101.360 200.000 101.960 ;
    END
  END peripheralBus_dataWrite[13]
  PIN peripheralBus_dataWrite[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 107.480 200.000 108.080 ;
    END
  END peripheralBus_dataWrite[14]
  PIN peripheralBus_dataWrite[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 114.280 200.000 114.880 ;
    END
  END peripheralBus_dataWrite[15]
  PIN peripheralBus_dataWrite[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 120.400 200.000 121.000 ;
    END
  END peripheralBus_dataWrite[16]
  PIN peripheralBus_dataWrite[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 126.520 200.000 127.120 ;
    END
  END peripheralBus_dataWrite[17]
  PIN peripheralBus_dataWrite[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 132.640 200.000 133.240 ;
    END
  END peripheralBus_dataWrite[18]
  PIN peripheralBus_dataWrite[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 139.440 200.000 140.040 ;
    END
  END peripheralBus_dataWrite[19]
  PIN peripheralBus_dataWrite[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 21.120 200.000 21.720 ;
    END
  END peripheralBus_dataWrite[1]
  PIN peripheralBus_dataWrite[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 145.560 200.000 146.160 ;
    END
  END peripheralBus_dataWrite[20]
  PIN peripheralBus_dataWrite[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 151.680 200.000 152.280 ;
    END
  END peripheralBus_dataWrite[21]
  PIN peripheralBus_dataWrite[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 158.480 200.000 159.080 ;
    END
  END peripheralBus_dataWrite[22]
  PIN peripheralBus_dataWrite[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 164.600 200.000 165.200 ;
    END
  END peripheralBus_dataWrite[23]
  PIN peripheralBus_dataWrite[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END peripheralBus_dataWrite[24]
  PIN peripheralBus_dataWrite[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 172.760 200.000 173.360 ;
    END
  END peripheralBus_dataWrite[25]
  PIN peripheralBus_dataWrite[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 200.000 177.440 ;
    END
  END peripheralBus_dataWrite[26]
  PIN peripheralBus_dataWrite[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 181.600 200.000 182.200 ;
    END
  END peripheralBus_dataWrite[27]
  PIN peripheralBus_dataWrite[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 185.680 200.000 186.280 ;
    END
  END peripheralBus_dataWrite[28]
  PIN peripheralBus_dataWrite[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 189.760 200.000 190.360 ;
    END
  END peripheralBus_dataWrite[29]
  PIN peripheralBus_dataWrite[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.960 200.000 30.560 ;
    END
  END peripheralBus_dataWrite[2]
  PIN peripheralBus_dataWrite[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.840 200.000 194.440 ;
    END
  END peripheralBus_dataWrite[30]
  PIN peripheralBus_dataWrite[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 197.920 200.000 198.520 ;
    END
  END peripheralBus_dataWrite[31]
  PIN peripheralBus_dataWrite[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 38.120 200.000 38.720 ;
    END
  END peripheralBus_dataWrite[3]
  PIN peripheralBus_dataWrite[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 44.240 200.000 44.840 ;
    END
  END peripheralBus_dataWrite[4]
  PIN peripheralBus_dataWrite[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.040 200.000 51.640 ;
    END
  END peripheralBus_dataWrite[5]
  PIN peripheralBus_dataWrite[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 57.160 200.000 57.760 ;
    END
  END peripheralBus_dataWrite[6]
  PIN peripheralBus_dataWrite[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 63.280 200.000 63.880 ;
    END
  END peripheralBus_dataWrite[7]
  PIN peripheralBus_dataWrite[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 70.080 200.000 70.680 ;
    END
  END peripheralBus_dataWrite[8]
  PIN peripheralBus_dataWrite[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 76.200 200.000 76.800 ;
    END
  END peripheralBus_dataWrite[9]
  PIN peripheralBus_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2.760 200.000 3.360 ;
    END
  END peripheralBus_oe
  PIN peripheralBus_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 4.800 200.000 5.400 ;
    END
  END peripheralBus_we
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END wb_data_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 6.500 194.120 187.920 ;
      LAYER met2 ;
        RECT 6.990 0.835 190.810 199.085 ;
      LAYER met3 ;
        RECT 4.400 198.920 196.000 199.065 ;
        RECT 4.400 198.200 195.600 198.920 ;
        RECT 4.000 197.560 195.600 198.200 ;
        RECT 4.400 197.520 195.600 197.560 ;
        RECT 4.400 196.880 196.000 197.520 ;
        RECT 4.400 196.160 195.600 196.880 ;
        RECT 4.000 195.520 195.600 196.160 ;
        RECT 4.400 195.480 195.600 195.520 ;
        RECT 4.400 194.840 196.000 195.480 ;
        RECT 4.400 194.120 195.600 194.840 ;
        RECT 4.000 193.480 195.600 194.120 ;
        RECT 4.400 193.440 195.600 193.480 ;
        RECT 4.400 192.800 196.000 193.440 ;
        RECT 4.400 192.080 195.600 192.800 ;
        RECT 4.000 191.440 195.600 192.080 ;
        RECT 4.400 191.400 195.600 191.440 ;
        RECT 4.400 190.760 196.000 191.400 ;
        RECT 4.400 190.040 195.600 190.760 ;
        RECT 4.000 189.400 195.600 190.040 ;
        RECT 4.400 189.360 195.600 189.400 ;
        RECT 4.400 188.720 196.000 189.360 ;
        RECT 4.400 188.000 195.600 188.720 ;
        RECT 4.000 187.360 195.600 188.000 ;
        RECT 4.400 187.320 195.600 187.360 ;
        RECT 4.400 186.680 196.000 187.320 ;
        RECT 4.400 185.960 195.600 186.680 ;
        RECT 4.000 185.320 195.600 185.960 ;
        RECT 4.400 185.280 195.600 185.320 ;
        RECT 4.400 184.640 196.000 185.280 ;
        RECT 4.400 183.920 195.600 184.640 ;
        RECT 4.000 183.280 195.600 183.920 ;
        RECT 4.400 183.240 195.600 183.280 ;
        RECT 4.400 182.600 196.000 183.240 ;
        RECT 4.400 181.880 195.600 182.600 ;
        RECT 4.000 181.240 195.600 181.880 ;
        RECT 4.400 181.200 195.600 181.240 ;
        RECT 4.400 180.560 196.000 181.200 ;
        RECT 4.400 179.840 195.600 180.560 ;
        RECT 4.000 179.200 195.600 179.840 ;
        RECT 4.400 179.160 195.600 179.200 ;
        RECT 4.400 177.840 196.000 179.160 ;
        RECT 4.400 177.800 195.600 177.840 ;
        RECT 4.000 177.160 195.600 177.800 ;
        RECT 4.400 176.440 195.600 177.160 ;
        RECT 4.400 175.800 196.000 176.440 ;
        RECT 4.400 175.760 195.600 175.800 ;
        RECT 4.000 175.120 195.600 175.760 ;
        RECT 4.400 174.400 195.600 175.120 ;
        RECT 4.400 173.760 196.000 174.400 ;
        RECT 4.400 173.720 195.600 173.760 ;
        RECT 4.000 173.080 195.600 173.720 ;
        RECT 4.400 172.360 195.600 173.080 ;
        RECT 4.400 171.720 196.000 172.360 ;
        RECT 4.400 171.680 195.600 171.720 ;
        RECT 4.000 171.040 195.600 171.680 ;
        RECT 4.400 170.320 195.600 171.040 ;
        RECT 4.400 169.680 196.000 170.320 ;
        RECT 4.400 169.640 195.600 169.680 ;
        RECT 4.000 169.000 195.600 169.640 ;
        RECT 4.400 168.280 195.600 169.000 ;
        RECT 4.400 167.640 196.000 168.280 ;
        RECT 4.400 167.600 195.600 167.640 ;
        RECT 4.000 166.960 195.600 167.600 ;
        RECT 4.400 166.240 195.600 166.960 ;
        RECT 4.400 165.600 196.000 166.240 ;
        RECT 4.400 165.560 195.600 165.600 ;
        RECT 4.000 164.920 195.600 165.560 ;
        RECT 4.400 164.200 195.600 164.920 ;
        RECT 4.400 163.560 196.000 164.200 ;
        RECT 4.400 163.520 195.600 163.560 ;
        RECT 4.000 162.880 195.600 163.520 ;
        RECT 4.400 162.160 195.600 162.880 ;
        RECT 4.400 161.520 196.000 162.160 ;
        RECT 4.400 161.480 195.600 161.520 ;
        RECT 4.000 160.840 195.600 161.480 ;
        RECT 4.400 160.120 195.600 160.840 ;
        RECT 4.400 159.480 196.000 160.120 ;
        RECT 4.400 159.440 195.600 159.480 ;
        RECT 4.000 158.800 195.600 159.440 ;
        RECT 4.400 158.080 195.600 158.800 ;
        RECT 4.400 157.440 196.000 158.080 ;
        RECT 4.400 157.400 195.600 157.440 ;
        RECT 4.000 156.760 195.600 157.400 ;
        RECT 4.400 156.040 195.600 156.760 ;
        RECT 4.400 155.360 196.000 156.040 ;
        RECT 4.000 154.720 196.000 155.360 ;
        RECT 4.400 153.320 195.600 154.720 ;
        RECT 4.000 152.680 196.000 153.320 ;
        RECT 4.400 151.280 195.600 152.680 ;
        RECT 4.000 150.640 196.000 151.280 ;
        RECT 4.400 149.240 195.600 150.640 ;
        RECT 4.000 148.600 196.000 149.240 ;
        RECT 4.400 147.200 195.600 148.600 ;
        RECT 4.000 146.560 196.000 147.200 ;
        RECT 4.400 145.160 195.600 146.560 ;
        RECT 4.000 144.520 196.000 145.160 ;
        RECT 4.400 143.120 195.600 144.520 ;
        RECT 4.000 142.480 196.000 143.120 ;
        RECT 4.400 141.080 195.600 142.480 ;
        RECT 4.000 140.440 196.000 141.080 ;
        RECT 4.400 139.040 195.600 140.440 ;
        RECT 4.000 138.400 196.000 139.040 ;
        RECT 4.400 137.000 195.600 138.400 ;
        RECT 4.000 136.360 196.000 137.000 ;
        RECT 4.400 134.960 195.600 136.360 ;
        RECT 4.400 133.640 196.000 134.960 ;
        RECT 4.400 133.600 195.600 133.640 ;
        RECT 4.000 132.960 195.600 133.600 ;
        RECT 4.400 132.240 195.600 132.960 ;
        RECT 4.400 131.600 196.000 132.240 ;
        RECT 4.400 131.560 195.600 131.600 ;
        RECT 4.000 130.920 195.600 131.560 ;
        RECT 4.400 130.200 195.600 130.920 ;
        RECT 4.400 129.560 196.000 130.200 ;
        RECT 4.400 129.520 195.600 129.560 ;
        RECT 4.000 128.880 195.600 129.520 ;
        RECT 4.400 128.160 195.600 128.880 ;
        RECT 4.400 127.520 196.000 128.160 ;
        RECT 4.400 127.480 195.600 127.520 ;
        RECT 4.000 126.840 195.600 127.480 ;
        RECT 4.400 126.120 195.600 126.840 ;
        RECT 4.400 125.480 196.000 126.120 ;
        RECT 4.400 125.440 195.600 125.480 ;
        RECT 4.000 124.800 195.600 125.440 ;
        RECT 4.400 124.080 195.600 124.800 ;
        RECT 4.400 123.440 196.000 124.080 ;
        RECT 4.400 123.400 195.600 123.440 ;
        RECT 4.000 122.760 195.600 123.400 ;
        RECT 4.400 122.040 195.600 122.760 ;
        RECT 4.400 121.400 196.000 122.040 ;
        RECT 4.400 121.360 195.600 121.400 ;
        RECT 4.000 120.720 195.600 121.360 ;
        RECT 4.400 120.000 195.600 120.720 ;
        RECT 4.400 119.360 196.000 120.000 ;
        RECT 4.400 119.320 195.600 119.360 ;
        RECT 4.000 118.680 195.600 119.320 ;
        RECT 4.400 117.960 195.600 118.680 ;
        RECT 4.400 117.320 196.000 117.960 ;
        RECT 4.400 117.280 195.600 117.320 ;
        RECT 4.000 116.640 195.600 117.280 ;
        RECT 4.400 115.920 195.600 116.640 ;
        RECT 4.400 115.280 196.000 115.920 ;
        RECT 4.400 115.240 195.600 115.280 ;
        RECT 4.000 114.600 195.600 115.240 ;
        RECT 4.400 113.880 195.600 114.600 ;
        RECT 4.400 113.240 196.000 113.880 ;
        RECT 4.400 113.200 195.600 113.240 ;
        RECT 4.000 112.560 195.600 113.200 ;
        RECT 4.400 111.840 195.600 112.560 ;
        RECT 4.400 111.160 196.000 111.840 ;
        RECT 4.000 110.520 196.000 111.160 ;
        RECT 4.400 109.120 195.600 110.520 ;
        RECT 4.000 108.480 196.000 109.120 ;
        RECT 4.400 107.080 195.600 108.480 ;
        RECT 4.000 106.440 196.000 107.080 ;
        RECT 4.400 105.040 195.600 106.440 ;
        RECT 4.000 104.400 196.000 105.040 ;
        RECT 4.400 103.000 195.600 104.400 ;
        RECT 4.000 102.360 196.000 103.000 ;
        RECT 4.400 100.960 195.600 102.360 ;
        RECT 4.000 100.320 196.000 100.960 ;
        RECT 4.400 98.920 195.600 100.320 ;
        RECT 4.000 98.280 196.000 98.920 ;
        RECT 4.400 96.880 195.600 98.280 ;
        RECT 4.000 96.240 196.000 96.880 ;
        RECT 4.400 94.840 195.600 96.240 ;
        RECT 4.000 94.200 196.000 94.840 ;
        RECT 4.400 92.800 195.600 94.200 ;
        RECT 4.000 92.160 196.000 92.800 ;
        RECT 4.400 90.760 195.600 92.160 ;
        RECT 4.000 90.120 196.000 90.760 ;
        RECT 4.400 89.440 196.000 90.120 ;
        RECT 4.400 88.720 195.600 89.440 ;
        RECT 4.000 88.080 195.600 88.720 ;
        RECT 4.400 88.040 195.600 88.080 ;
        RECT 4.400 87.400 196.000 88.040 ;
        RECT 4.400 86.680 195.600 87.400 ;
        RECT 4.000 86.040 195.600 86.680 ;
        RECT 4.400 86.000 195.600 86.040 ;
        RECT 4.400 85.360 196.000 86.000 ;
        RECT 4.400 84.640 195.600 85.360 ;
        RECT 4.000 84.000 195.600 84.640 ;
        RECT 4.400 83.960 195.600 84.000 ;
        RECT 4.400 83.320 196.000 83.960 ;
        RECT 4.400 82.600 195.600 83.320 ;
        RECT 4.000 81.960 195.600 82.600 ;
        RECT 4.400 81.920 195.600 81.960 ;
        RECT 4.400 81.280 196.000 81.920 ;
        RECT 4.400 80.560 195.600 81.280 ;
        RECT 4.000 79.920 195.600 80.560 ;
        RECT 4.400 79.880 195.600 79.920 ;
        RECT 4.400 79.240 196.000 79.880 ;
        RECT 4.400 78.520 195.600 79.240 ;
        RECT 4.000 77.880 195.600 78.520 ;
        RECT 4.400 77.840 195.600 77.880 ;
        RECT 4.400 77.200 196.000 77.840 ;
        RECT 4.400 76.480 195.600 77.200 ;
        RECT 4.000 75.840 195.600 76.480 ;
        RECT 4.400 75.800 195.600 75.840 ;
        RECT 4.400 75.160 196.000 75.800 ;
        RECT 4.400 74.440 195.600 75.160 ;
        RECT 4.000 73.800 195.600 74.440 ;
        RECT 4.400 73.760 195.600 73.800 ;
        RECT 4.400 73.120 196.000 73.760 ;
        RECT 4.400 72.400 195.600 73.120 ;
        RECT 4.000 71.760 195.600 72.400 ;
        RECT 4.400 71.720 195.600 71.760 ;
        RECT 4.400 71.080 196.000 71.720 ;
        RECT 4.400 70.360 195.600 71.080 ;
        RECT 4.000 69.720 195.600 70.360 ;
        RECT 4.400 69.680 195.600 69.720 ;
        RECT 4.400 69.040 196.000 69.680 ;
        RECT 4.400 67.640 195.600 69.040 ;
        RECT 4.400 66.960 196.000 67.640 ;
        RECT 4.000 66.320 196.000 66.960 ;
        RECT 4.400 64.920 195.600 66.320 ;
        RECT 4.000 64.280 196.000 64.920 ;
        RECT 4.400 62.880 195.600 64.280 ;
        RECT 4.000 62.240 196.000 62.880 ;
        RECT 4.400 60.840 195.600 62.240 ;
        RECT 4.000 60.200 196.000 60.840 ;
        RECT 4.400 58.800 195.600 60.200 ;
        RECT 4.000 58.160 196.000 58.800 ;
        RECT 4.400 56.760 195.600 58.160 ;
        RECT 4.000 56.120 196.000 56.760 ;
        RECT 4.400 54.720 195.600 56.120 ;
        RECT 4.000 54.080 196.000 54.720 ;
        RECT 4.400 52.680 195.600 54.080 ;
        RECT 4.000 52.040 196.000 52.680 ;
        RECT 4.400 50.640 195.600 52.040 ;
        RECT 4.000 50.000 196.000 50.640 ;
        RECT 4.400 48.600 195.600 50.000 ;
        RECT 4.000 47.960 196.000 48.600 ;
        RECT 4.400 46.560 195.600 47.960 ;
        RECT 4.000 45.920 196.000 46.560 ;
        RECT 4.400 45.240 196.000 45.920 ;
        RECT 4.400 44.520 195.600 45.240 ;
        RECT 4.000 43.880 195.600 44.520 ;
        RECT 4.400 43.840 195.600 43.880 ;
        RECT 4.400 43.200 196.000 43.840 ;
        RECT 4.400 42.480 195.600 43.200 ;
        RECT 4.000 41.840 195.600 42.480 ;
        RECT 4.400 41.800 195.600 41.840 ;
        RECT 4.400 41.160 196.000 41.800 ;
        RECT 4.400 40.440 195.600 41.160 ;
        RECT 4.000 39.800 195.600 40.440 ;
        RECT 4.400 39.760 195.600 39.800 ;
        RECT 4.400 39.120 196.000 39.760 ;
        RECT 4.400 38.400 195.600 39.120 ;
        RECT 4.000 37.760 195.600 38.400 ;
        RECT 4.400 37.720 195.600 37.760 ;
        RECT 4.400 37.080 196.000 37.720 ;
        RECT 4.400 36.360 195.600 37.080 ;
        RECT 4.000 35.720 195.600 36.360 ;
        RECT 4.400 35.680 195.600 35.720 ;
        RECT 4.400 35.040 196.000 35.680 ;
        RECT 4.400 34.320 195.600 35.040 ;
        RECT 4.000 33.680 195.600 34.320 ;
        RECT 4.400 33.640 195.600 33.680 ;
        RECT 4.400 33.000 196.000 33.640 ;
        RECT 4.400 32.280 195.600 33.000 ;
        RECT 4.000 31.640 195.600 32.280 ;
        RECT 4.400 31.600 195.600 31.640 ;
        RECT 4.400 30.960 196.000 31.600 ;
        RECT 4.400 30.240 195.600 30.960 ;
        RECT 4.000 29.600 195.600 30.240 ;
        RECT 4.400 29.560 195.600 29.600 ;
        RECT 4.400 28.920 196.000 29.560 ;
        RECT 4.400 28.200 195.600 28.920 ;
        RECT 4.000 27.560 195.600 28.200 ;
        RECT 4.400 27.520 195.600 27.560 ;
        RECT 4.400 26.880 196.000 27.520 ;
        RECT 4.400 26.160 195.600 26.880 ;
        RECT 4.000 25.520 195.600 26.160 ;
        RECT 4.400 25.480 195.600 25.520 ;
        RECT 4.400 24.840 196.000 25.480 ;
        RECT 4.400 24.120 195.600 24.840 ;
        RECT 4.000 23.480 195.600 24.120 ;
        RECT 4.400 23.440 195.600 23.480 ;
        RECT 4.400 22.120 196.000 23.440 ;
        RECT 4.400 22.080 195.600 22.120 ;
        RECT 4.000 21.440 195.600 22.080 ;
        RECT 4.400 20.720 195.600 21.440 ;
        RECT 4.400 20.080 196.000 20.720 ;
        RECT 4.400 20.040 195.600 20.080 ;
        RECT 4.000 19.400 195.600 20.040 ;
        RECT 4.400 18.680 195.600 19.400 ;
        RECT 4.400 18.040 196.000 18.680 ;
        RECT 4.400 18.000 195.600 18.040 ;
        RECT 4.000 17.360 195.600 18.000 ;
        RECT 4.400 16.640 195.600 17.360 ;
        RECT 4.400 16.000 196.000 16.640 ;
        RECT 4.400 15.960 195.600 16.000 ;
        RECT 4.000 15.320 195.600 15.960 ;
        RECT 4.400 14.600 195.600 15.320 ;
        RECT 4.400 13.960 196.000 14.600 ;
        RECT 4.400 13.920 195.600 13.960 ;
        RECT 4.000 13.280 195.600 13.920 ;
        RECT 4.400 12.560 195.600 13.280 ;
        RECT 4.400 11.920 196.000 12.560 ;
        RECT 4.400 11.880 195.600 11.920 ;
        RECT 4.000 11.240 195.600 11.880 ;
        RECT 4.400 10.520 195.600 11.240 ;
        RECT 4.400 9.880 196.000 10.520 ;
        RECT 4.400 9.840 195.600 9.880 ;
        RECT 4.000 9.200 195.600 9.840 ;
        RECT 4.400 8.480 195.600 9.200 ;
        RECT 4.400 7.840 196.000 8.480 ;
        RECT 4.400 7.800 195.600 7.840 ;
        RECT 4.000 7.160 195.600 7.800 ;
        RECT 4.400 6.440 195.600 7.160 ;
        RECT 4.400 5.800 196.000 6.440 ;
        RECT 4.400 5.760 195.600 5.800 ;
        RECT 4.000 5.120 195.600 5.760 ;
        RECT 4.400 4.400 195.600 5.120 ;
        RECT 4.400 3.760 196.000 4.400 ;
        RECT 4.400 3.720 195.600 3.760 ;
        RECT 4.000 3.080 195.600 3.720 ;
        RECT 4.400 2.360 195.600 3.080 ;
        RECT 4.400 1.720 196.000 2.360 ;
        RECT 4.400 0.855 195.600 1.720 ;
  END
END WBPeripheralBusInterface
END LIBRARY

