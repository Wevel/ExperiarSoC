magic
tech sky130A
magscale 1 2
timestamp 1652994636
<< obsli1 >>
rect 1104 2159 118864 37553
<< obsm1 >>
rect 382 1368 119586 37584
<< metal2 >>
rect 1766 39200 1822 40000
rect 5262 39200 5318 40000
rect 8758 39200 8814 40000
rect 12346 39200 12402 40000
rect 15842 39200 15898 40000
rect 19338 39200 19394 40000
rect 22926 39200 22982 40000
rect 26422 39200 26478 40000
rect 29918 39200 29974 40000
rect 33506 39200 33562 40000
rect 37002 39200 37058 40000
rect 40498 39200 40554 40000
rect 44086 39200 44142 40000
rect 47582 39200 47638 40000
rect 51078 39200 51134 40000
rect 54666 39200 54722 40000
rect 58162 39200 58218 40000
rect 61750 39200 61806 40000
rect 65246 39200 65302 40000
rect 68742 39200 68798 40000
rect 72330 39200 72386 40000
rect 75826 39200 75882 40000
rect 79322 39200 79378 40000
rect 82910 39200 82966 40000
rect 86406 39200 86462 40000
rect 89902 39200 89958 40000
rect 93490 39200 93546 40000
rect 96986 39200 97042 40000
rect 100482 39200 100538 40000
rect 104070 39200 104126 40000
rect 107566 39200 107622 40000
rect 111062 39200 111118 40000
rect 114650 39200 114706 40000
rect 118146 39200 118202 40000
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2778 0 2834 800
rect 3606 0 3662 800
rect 4434 0 4490 800
rect 5262 0 5318 800
rect 6090 0 6146 800
rect 6918 0 6974 800
rect 7746 0 7802 800
rect 8574 0 8630 800
rect 9402 0 9458 800
rect 10230 0 10286 800
rect 11058 0 11114 800
rect 11886 0 11942 800
rect 12622 0 12678 800
rect 13450 0 13506 800
rect 14278 0 14334 800
rect 15106 0 15162 800
rect 15934 0 15990 800
rect 16762 0 16818 800
rect 17590 0 17646 800
rect 18418 0 18474 800
rect 19246 0 19302 800
rect 20074 0 20130 800
rect 20902 0 20958 800
rect 21730 0 21786 800
rect 22558 0 22614 800
rect 23386 0 23442 800
rect 24214 0 24270 800
rect 24950 0 25006 800
rect 25778 0 25834 800
rect 26606 0 26662 800
rect 27434 0 27490 800
rect 28262 0 28318 800
rect 29090 0 29146 800
rect 29918 0 29974 800
rect 30746 0 30802 800
rect 31574 0 31630 800
rect 32402 0 32458 800
rect 33230 0 33286 800
rect 34058 0 34114 800
rect 34886 0 34942 800
rect 35714 0 35770 800
rect 36450 0 36506 800
rect 37278 0 37334 800
rect 38106 0 38162 800
rect 38934 0 38990 800
rect 39762 0 39818 800
rect 40590 0 40646 800
rect 41418 0 41474 800
rect 42246 0 42302 800
rect 43074 0 43130 800
rect 43902 0 43958 800
rect 44730 0 44786 800
rect 45558 0 45614 800
rect 46386 0 46442 800
rect 47214 0 47270 800
rect 48042 0 48098 800
rect 48778 0 48834 800
rect 49606 0 49662 800
rect 50434 0 50490 800
rect 51262 0 51318 800
rect 52090 0 52146 800
rect 52918 0 52974 800
rect 53746 0 53802 800
rect 54574 0 54630 800
rect 55402 0 55458 800
rect 56230 0 56286 800
rect 57058 0 57114 800
rect 57886 0 57942 800
rect 58714 0 58770 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61106 0 61162 800
rect 61934 0 61990 800
rect 62762 0 62818 800
rect 63590 0 63646 800
rect 64418 0 64474 800
rect 65246 0 65302 800
rect 66074 0 66130 800
rect 66902 0 66958 800
rect 67730 0 67786 800
rect 68558 0 68614 800
rect 69386 0 69442 800
rect 70214 0 70270 800
rect 71042 0 71098 800
rect 71870 0 71926 800
rect 72606 0 72662 800
rect 73434 0 73490 800
rect 74262 0 74318 800
rect 75090 0 75146 800
rect 75918 0 75974 800
rect 76746 0 76802 800
rect 77574 0 77630 800
rect 78402 0 78458 800
rect 79230 0 79286 800
rect 80058 0 80114 800
rect 80886 0 80942 800
rect 81714 0 81770 800
rect 82542 0 82598 800
rect 83370 0 83426 800
rect 84198 0 84254 800
rect 84934 0 84990 800
rect 85762 0 85818 800
rect 86590 0 86646 800
rect 87418 0 87474 800
rect 88246 0 88302 800
rect 89074 0 89130 800
rect 89902 0 89958 800
rect 90730 0 90786 800
rect 91558 0 91614 800
rect 92386 0 92442 800
rect 93214 0 93270 800
rect 94042 0 94098 800
rect 94870 0 94926 800
rect 95698 0 95754 800
rect 96434 0 96490 800
rect 97262 0 97318 800
rect 98090 0 98146 800
rect 98918 0 98974 800
rect 99746 0 99802 800
rect 100574 0 100630 800
rect 101402 0 101458 800
rect 102230 0 102286 800
rect 103058 0 103114 800
rect 103886 0 103942 800
rect 104714 0 104770 800
rect 105542 0 105598 800
rect 106370 0 106426 800
rect 107198 0 107254 800
rect 108026 0 108082 800
rect 108762 0 108818 800
rect 109590 0 109646 800
rect 110418 0 110474 800
rect 111246 0 111302 800
rect 112074 0 112130 800
rect 112902 0 112958 800
rect 113730 0 113786 800
rect 114558 0 114614 800
rect 115386 0 115442 800
rect 116214 0 116270 800
rect 117042 0 117098 800
rect 117870 0 117926 800
rect 118698 0 118754 800
rect 119526 0 119582 800
<< obsm2 >>
rect 388 39144 1710 39273
rect 1878 39144 5206 39273
rect 5374 39144 8702 39273
rect 8870 39144 12290 39273
rect 12458 39144 15786 39273
rect 15954 39144 19282 39273
rect 19450 39144 22870 39273
rect 23038 39144 26366 39273
rect 26534 39144 29862 39273
rect 30030 39144 33450 39273
rect 33618 39144 36946 39273
rect 37114 39144 40442 39273
rect 40610 39144 44030 39273
rect 44198 39144 47526 39273
rect 47694 39144 51022 39273
rect 51190 39144 54610 39273
rect 54778 39144 58106 39273
rect 58274 39144 61694 39273
rect 61862 39144 65190 39273
rect 65358 39144 68686 39273
rect 68854 39144 72274 39273
rect 72442 39144 75770 39273
rect 75938 39144 79266 39273
rect 79434 39144 82854 39273
rect 83022 39144 86350 39273
rect 86518 39144 89846 39273
rect 90014 39144 93434 39273
rect 93602 39144 96930 39273
rect 97098 39144 100426 39273
rect 100594 39144 104014 39273
rect 104182 39144 107510 39273
rect 107678 39144 111006 39273
rect 111174 39144 114594 39273
rect 114762 39144 118090 39273
rect 118258 39144 119580 39273
rect 388 856 119580 39144
rect 498 575 1066 856
rect 1234 575 1894 856
rect 2062 575 2722 856
rect 2890 575 3550 856
rect 3718 575 4378 856
rect 4546 575 5206 856
rect 5374 575 6034 856
rect 6202 575 6862 856
rect 7030 575 7690 856
rect 7858 575 8518 856
rect 8686 575 9346 856
rect 9514 575 10174 856
rect 10342 575 11002 856
rect 11170 575 11830 856
rect 11998 575 12566 856
rect 12734 575 13394 856
rect 13562 575 14222 856
rect 14390 575 15050 856
rect 15218 575 15878 856
rect 16046 575 16706 856
rect 16874 575 17534 856
rect 17702 575 18362 856
rect 18530 575 19190 856
rect 19358 575 20018 856
rect 20186 575 20846 856
rect 21014 575 21674 856
rect 21842 575 22502 856
rect 22670 575 23330 856
rect 23498 575 24158 856
rect 24326 575 24894 856
rect 25062 575 25722 856
rect 25890 575 26550 856
rect 26718 575 27378 856
rect 27546 575 28206 856
rect 28374 575 29034 856
rect 29202 575 29862 856
rect 30030 575 30690 856
rect 30858 575 31518 856
rect 31686 575 32346 856
rect 32514 575 33174 856
rect 33342 575 34002 856
rect 34170 575 34830 856
rect 34998 575 35658 856
rect 35826 575 36394 856
rect 36562 575 37222 856
rect 37390 575 38050 856
rect 38218 575 38878 856
rect 39046 575 39706 856
rect 39874 575 40534 856
rect 40702 575 41362 856
rect 41530 575 42190 856
rect 42358 575 43018 856
rect 43186 575 43846 856
rect 44014 575 44674 856
rect 44842 575 45502 856
rect 45670 575 46330 856
rect 46498 575 47158 856
rect 47326 575 47986 856
rect 48154 575 48722 856
rect 48890 575 49550 856
rect 49718 575 50378 856
rect 50546 575 51206 856
rect 51374 575 52034 856
rect 52202 575 52862 856
rect 53030 575 53690 856
rect 53858 575 54518 856
rect 54686 575 55346 856
rect 55514 575 56174 856
rect 56342 575 57002 856
rect 57170 575 57830 856
rect 57998 575 58658 856
rect 58826 575 59486 856
rect 59654 575 60314 856
rect 60482 575 61050 856
rect 61218 575 61878 856
rect 62046 575 62706 856
rect 62874 575 63534 856
rect 63702 575 64362 856
rect 64530 575 65190 856
rect 65358 575 66018 856
rect 66186 575 66846 856
rect 67014 575 67674 856
rect 67842 575 68502 856
rect 68670 575 69330 856
rect 69498 575 70158 856
rect 70326 575 70986 856
rect 71154 575 71814 856
rect 71982 575 72550 856
rect 72718 575 73378 856
rect 73546 575 74206 856
rect 74374 575 75034 856
rect 75202 575 75862 856
rect 76030 575 76690 856
rect 76858 575 77518 856
rect 77686 575 78346 856
rect 78514 575 79174 856
rect 79342 575 80002 856
rect 80170 575 80830 856
rect 80998 575 81658 856
rect 81826 575 82486 856
rect 82654 575 83314 856
rect 83482 575 84142 856
rect 84310 575 84878 856
rect 85046 575 85706 856
rect 85874 575 86534 856
rect 86702 575 87362 856
rect 87530 575 88190 856
rect 88358 575 89018 856
rect 89186 575 89846 856
rect 90014 575 90674 856
rect 90842 575 91502 856
rect 91670 575 92330 856
rect 92498 575 93158 856
rect 93326 575 93986 856
rect 94154 575 94814 856
rect 94982 575 95642 856
rect 95810 575 96378 856
rect 96546 575 97206 856
rect 97374 575 98034 856
rect 98202 575 98862 856
rect 99030 575 99690 856
rect 99858 575 100518 856
rect 100686 575 101346 856
rect 101514 575 102174 856
rect 102342 575 103002 856
rect 103170 575 103830 856
rect 103998 575 104658 856
rect 104826 575 105486 856
rect 105654 575 106314 856
rect 106482 575 107142 856
rect 107310 575 107970 856
rect 108138 575 108706 856
rect 108874 575 109534 856
rect 109702 575 110362 856
rect 110530 575 111190 856
rect 111358 575 112018 856
rect 112186 575 112846 856
rect 113014 575 113674 856
rect 113842 575 114502 856
rect 114670 575 115330 856
rect 115498 575 116158 856
rect 116326 575 116986 856
rect 117154 575 117814 856
rect 117982 575 118642 856
rect 118810 575 119470 856
<< metal3 >>
rect 0 39040 800 39160
rect 119200 39176 120000 39296
rect 119200 37816 120000 37936
rect 0 37136 800 37256
rect 119200 36456 120000 36576
rect 0 35232 800 35352
rect 119200 35096 120000 35216
rect 119200 33872 120000 33992
rect 0 33328 800 33448
rect 119200 32512 120000 32632
rect 0 31424 800 31544
rect 119200 31152 120000 31272
rect 119200 29792 120000 29912
rect 0 29520 800 29640
rect 119200 28432 120000 28552
rect 0 27616 800 27736
rect 119200 27208 120000 27328
rect 0 25712 800 25832
rect 119200 25848 120000 25968
rect 119200 24488 120000 24608
rect 0 23808 800 23928
rect 119200 23128 120000 23248
rect 0 21904 800 22024
rect 119200 21768 120000 21888
rect 119200 20544 120000 20664
rect 0 20000 800 20120
rect 119200 19184 120000 19304
rect 0 18096 800 18216
rect 119200 17824 120000 17944
rect 119200 16464 120000 16584
rect 0 16192 800 16312
rect 119200 15104 120000 15224
rect 0 14288 800 14408
rect 119200 13880 120000 14000
rect 0 12384 800 12504
rect 119200 12520 120000 12640
rect 119200 11160 120000 11280
rect 0 10480 800 10600
rect 119200 9800 120000 9920
rect 0 8576 800 8696
rect 119200 8440 120000 8560
rect 119200 7216 120000 7336
rect 0 6672 800 6792
rect 119200 5856 120000 5976
rect 0 4768 800 4888
rect 119200 4496 120000 4616
rect 119200 3136 120000 3256
rect 0 2864 800 2984
rect 119200 1776 120000 1896
rect 0 960 800 1080
rect 119200 552 120000 672
<< obsm3 >>
rect 800 39240 119120 39269
rect 880 39096 119120 39240
rect 880 38960 119200 39096
rect 800 38016 119200 38960
rect 800 37736 119120 38016
rect 800 37336 119200 37736
rect 880 37056 119200 37336
rect 800 36656 119200 37056
rect 800 36376 119120 36656
rect 800 35432 119200 36376
rect 880 35296 119200 35432
rect 880 35152 119120 35296
rect 800 35016 119120 35152
rect 800 34072 119200 35016
rect 800 33792 119120 34072
rect 800 33528 119200 33792
rect 880 33248 119200 33528
rect 800 32712 119200 33248
rect 800 32432 119120 32712
rect 800 31624 119200 32432
rect 880 31352 119200 31624
rect 880 31344 119120 31352
rect 800 31072 119120 31344
rect 800 29992 119200 31072
rect 800 29720 119120 29992
rect 880 29712 119120 29720
rect 880 29440 119200 29712
rect 800 28632 119200 29440
rect 800 28352 119120 28632
rect 800 27816 119200 28352
rect 880 27536 119200 27816
rect 800 27408 119200 27536
rect 800 27128 119120 27408
rect 800 26048 119200 27128
rect 800 25912 119120 26048
rect 880 25768 119120 25912
rect 880 25632 119200 25768
rect 800 24688 119200 25632
rect 800 24408 119120 24688
rect 800 24008 119200 24408
rect 880 23728 119200 24008
rect 800 23328 119200 23728
rect 800 23048 119120 23328
rect 800 22104 119200 23048
rect 880 21968 119200 22104
rect 880 21824 119120 21968
rect 800 21688 119120 21824
rect 800 20744 119200 21688
rect 800 20464 119120 20744
rect 800 20200 119200 20464
rect 880 19920 119200 20200
rect 800 19384 119200 19920
rect 800 19104 119120 19384
rect 800 18296 119200 19104
rect 880 18024 119200 18296
rect 880 18016 119120 18024
rect 800 17744 119120 18016
rect 800 16664 119200 17744
rect 800 16392 119120 16664
rect 880 16384 119120 16392
rect 880 16112 119200 16384
rect 800 15304 119200 16112
rect 800 15024 119120 15304
rect 800 14488 119200 15024
rect 880 14208 119200 14488
rect 800 14080 119200 14208
rect 800 13800 119120 14080
rect 800 12720 119200 13800
rect 800 12584 119120 12720
rect 880 12440 119120 12584
rect 880 12304 119200 12440
rect 800 11360 119200 12304
rect 800 11080 119120 11360
rect 800 10680 119200 11080
rect 880 10400 119200 10680
rect 800 10000 119200 10400
rect 800 9720 119120 10000
rect 800 8776 119200 9720
rect 880 8640 119200 8776
rect 880 8496 119120 8640
rect 800 8360 119120 8496
rect 800 7416 119200 8360
rect 800 7136 119120 7416
rect 800 6872 119200 7136
rect 880 6592 119200 6872
rect 800 6056 119200 6592
rect 800 5776 119120 6056
rect 800 4968 119200 5776
rect 880 4696 119200 4968
rect 880 4688 119120 4696
rect 800 4416 119120 4688
rect 800 3336 119200 4416
rect 800 3064 119120 3336
rect 880 3056 119120 3064
rect 880 2784 119200 3056
rect 800 1976 119200 2784
rect 800 1696 119120 1976
rect 800 1160 119200 1696
rect 880 880 119200 1160
rect 800 752 119200 880
rect 800 579 119120 752
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
rect 65648 2128 65968 37584
rect 81008 2128 81328 37584
rect 96368 2128 96688 37584
rect 111728 2128 112048 37584
<< labels >>
rlabel metal2 s 1766 39200 1822 40000 6 flash_csb
port 1 nsew signal output
rlabel metal2 s 5262 39200 5318 40000 6 flash_io0_read
port 2 nsew signal input
rlabel metal2 s 8758 39200 8814 40000 6 flash_io0_we
port 3 nsew signal output
rlabel metal2 s 12346 39200 12402 40000 6 flash_io0_write
port 4 nsew signal output
rlabel metal2 s 15842 39200 15898 40000 6 flash_io1_read
port 5 nsew signal input
rlabel metal2 s 19338 39200 19394 40000 6 flash_io1_we
port 6 nsew signal output
rlabel metal2 s 22926 39200 22982 40000 6 flash_io1_write
port 7 nsew signal output
rlabel metal2 s 26422 39200 26478 40000 6 flash_sck
port 8 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 sram_addr0[0]
port 9 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 sram_addr0[1]
port 10 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 sram_addr0[2]
port 11 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 sram_addr0[3]
port 12 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 sram_addr0[4]
port 13 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 sram_addr0[5]
port 14 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 sram_addr0[6]
port 15 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 sram_addr0[7]
port 16 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 sram_addr0[8]
port 17 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 sram_addr1[0]
port 18 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 sram_addr1[1]
port 19 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 sram_addr1[2]
port 20 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 sram_addr1[3]
port 21 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 sram_addr1[4]
port 22 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 sram_addr1[5]
port 23 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 sram_addr1[6]
port 24 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 sram_addr1[7]
port 25 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 sram_addr1[8]
port 26 nsew signal output
rlabel metal2 s 386 0 442 800 6 sram_clk0
port 27 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 sram_clk1
port 28 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 sram_csb0
port 29 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 sram_csb1
port 30 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 sram_din0[0]
port 31 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 sram_din0[10]
port 32 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 sram_din0[11]
port 33 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 sram_din0[12]
port 34 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 sram_din0[13]
port 35 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 sram_din0[14]
port 36 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 sram_din0[15]
port 37 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 sram_din0[16]
port 38 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 sram_din0[17]
port 39 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 sram_din0[18]
port 40 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 sram_din0[19]
port 41 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 sram_din0[1]
port 42 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 sram_din0[20]
port 43 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 sram_din0[21]
port 44 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 sram_din0[22]
port 45 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 sram_din0[23]
port 46 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 sram_din0[24]
port 47 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 sram_din0[25]
port 48 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 sram_din0[26]
port 49 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 sram_din0[27]
port 50 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 sram_din0[28]
port 51 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 sram_din0[29]
port 52 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 sram_din0[2]
port 53 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 sram_din0[30]
port 54 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 sram_din0[31]
port 55 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 sram_din0[3]
port 56 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 sram_din0[4]
port 57 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 sram_din0[5]
port 58 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 sram_din0[6]
port 59 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 sram_din0[7]
port 60 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 sram_din0[8]
port 61 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 sram_din0[9]
port 62 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 sram_dout0[0]
port 63 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 sram_dout0[10]
port 64 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 sram_dout0[11]
port 65 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 sram_dout0[12]
port 66 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 sram_dout0[13]
port 67 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 sram_dout0[14]
port 68 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 sram_dout0[15]
port 69 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 sram_dout0[16]
port 70 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 sram_dout0[17]
port 71 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 sram_dout0[18]
port 72 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 sram_dout0[19]
port 73 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 sram_dout0[1]
port 74 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 sram_dout0[20]
port 75 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 sram_dout0[21]
port 76 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 sram_dout0[22]
port 77 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 sram_dout0[23]
port 78 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 sram_dout0[24]
port 79 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 sram_dout0[25]
port 80 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 sram_dout0[26]
port 81 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 sram_dout0[27]
port 82 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 sram_dout0[28]
port 83 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 sram_dout0[29]
port 84 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 sram_dout0[2]
port 85 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 sram_dout0[30]
port 86 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 sram_dout0[31]
port 87 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 sram_dout0[3]
port 88 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 sram_dout0[4]
port 89 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 sram_dout0[5]
port 90 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 sram_dout0[6]
port 91 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 sram_dout0[7]
port 92 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 sram_dout0[8]
port 93 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 sram_dout0[9]
port 94 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 sram_dout1[0]
port 95 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 sram_dout1[10]
port 96 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 sram_dout1[11]
port 97 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 sram_dout1[12]
port 98 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 sram_dout1[13]
port 99 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 sram_dout1[14]
port 100 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 sram_dout1[15]
port 101 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 sram_dout1[16]
port 102 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 sram_dout1[17]
port 103 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 sram_dout1[18]
port 104 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 sram_dout1[19]
port 105 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 sram_dout1[1]
port 106 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 sram_dout1[20]
port 107 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 sram_dout1[21]
port 108 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 sram_dout1[22]
port 109 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 sram_dout1[23]
port 110 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 sram_dout1[24]
port 111 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 sram_dout1[25]
port 112 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 sram_dout1[26]
port 113 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 sram_dout1[27]
port 114 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 sram_dout1[28]
port 115 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 sram_dout1[29]
port 116 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 sram_dout1[2]
port 117 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 sram_dout1[30]
port 118 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 sram_dout1[31]
port 119 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 sram_dout1[3]
port 120 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 sram_dout1[4]
port 121 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 sram_dout1[5]
port 122 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 sram_dout1[6]
port 123 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 sram_dout1[7]
port 124 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 sram_dout1[8]
port 125 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 sram_dout1[9]
port 126 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 sram_web0
port 127 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 sram_wmask0[0]
port 128 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 sram_wmask0[1]
port 129 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 sram_wmask0[2]
port 130 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 sram_wmask0[3]
port 131 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 132 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 37584 6 vssd1
port 133 nsew ground bidirectional
rlabel metal2 s 101402 0 101458 800 6 wb_ack_o
port 134 nsew signal output
rlabel metal3 s 0 960 800 1080 6 wb_adr_i[0]
port 135 nsew signal input
rlabel metal3 s 119200 19184 120000 19304 6 wb_adr_i[10]
port 136 nsew signal input
rlabel metal2 s 79322 39200 79378 40000 6 wb_adr_i[11]
port 137 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 wb_adr_i[12]
port 138 nsew signal input
rlabel metal3 s 119200 20544 120000 20664 6 wb_adr_i[13]
port 139 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wb_adr_i[14]
port 140 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 wb_adr_i[15]
port 141 nsew signal input
rlabel metal2 s 89902 39200 89958 40000 6 wb_adr_i[16]
port 142 nsew signal input
rlabel metal2 s 96986 39200 97042 40000 6 wb_adr_i[17]
port 143 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 wb_adr_i[18]
port 144 nsew signal input
rlabel metal3 s 119200 25848 120000 25968 6 wb_adr_i[19]
port 145 nsew signal input
rlabel metal3 s 119200 5856 120000 5976 6 wb_adr_i[1]
port 146 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 wb_adr_i[20]
port 147 nsew signal input
rlabel metal2 s 107566 39200 107622 40000 6 wb_adr_i[21]
port 148 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 wb_adr_i[22]
port 149 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 wb_adr_i[23]
port 150 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 wb_adr_i[2]
port 151 nsew signal input
rlabel metal3 s 119200 12520 120000 12640 6 wb_adr_i[3]
port 152 nsew signal input
rlabel metal2 s 47582 39200 47638 40000 6 wb_adr_i[4]
port 153 nsew signal input
rlabel metal2 s 54666 39200 54722 40000 6 wb_adr_i[5]
port 154 nsew signal input
rlabel metal2 s 58162 39200 58218 40000 6 wb_adr_i[6]
port 155 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 wb_adr_i[7]
port 156 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 wb_adr_i[8]
port 157 nsew signal input
rlabel metal2 s 72330 39200 72386 40000 6 wb_adr_i[9]
port 158 nsew signal input
rlabel metal2 s 29918 39200 29974 40000 6 wb_clk_i
port 159 nsew signal input
rlabel metal3 s 119200 552 120000 672 6 wb_cyc_i
port 160 nsew signal input
rlabel metal2 s 37002 39200 37058 40000 6 wb_data_i[0]
port 161 nsew signal input
rlabel metal2 s 75826 39200 75882 40000 6 wb_data_i[10]
port 162 nsew signal input
rlabel metal2 s 82910 39200 82966 40000 6 wb_data_i[11]
port 163 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 wb_data_i[12]
port 164 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 wb_data_i[13]
port 165 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 wb_data_i[14]
port 166 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 wb_data_i[15]
port 167 nsew signal input
rlabel metal2 s 93490 39200 93546 40000 6 wb_data_i[16]
port 168 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[17]
port 169 nsew signal input
rlabel metal3 s 119200 24488 120000 24608 6 wb_data_i[18]
port 170 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_data_i[19]
port 171 nsew signal input
rlabel metal3 s 119200 7216 120000 7336 6 wb_data_i[1]
port 172 nsew signal input
rlabel metal2 s 104070 39200 104126 40000 6 wb_data_i[20]
port 173 nsew signal input
rlabel metal2 s 111062 39200 111118 40000 6 wb_data_i[21]
port 174 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wb_data_i[22]
port 175 nsew signal input
rlabel metal3 s 119200 28432 120000 28552 6 wb_data_i[23]
port 176 nsew signal input
rlabel metal3 s 119200 29792 120000 29912 6 wb_data_i[24]
port 177 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 wb_data_i[25]
port 178 nsew signal input
rlabel metal2 s 118146 39200 118202 40000 6 wb_data_i[26]
port 179 nsew signal input
rlabel metal3 s 119200 33872 120000 33992 6 wb_data_i[27]
port 180 nsew signal input
rlabel metal3 s 119200 36456 120000 36576 6 wb_data_i[28]
port 181 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 wb_data_i[29]
port 182 nsew signal input
rlabel metal3 s 119200 9800 120000 9920 6 wb_data_i[2]
port 183 nsew signal input
rlabel metal3 s 0 37136 800 37256 6 wb_data_i[30]
port 184 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 wb_data_i[31]
port 185 nsew signal input
rlabel metal2 s 40498 39200 40554 40000 6 wb_data_i[3]
port 186 nsew signal input
rlabel metal2 s 51078 39200 51134 40000 6 wb_data_i[4]
port 187 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 wb_data_i[5]
port 188 nsew signal input
rlabel metal2 s 61750 39200 61806 40000 6 wb_data_i[6]
port 189 nsew signal input
rlabel metal2 s 65246 39200 65302 40000 6 wb_data_i[7]
port 190 nsew signal input
rlabel metal3 s 119200 15104 120000 15224 6 wb_data_i[8]
port 191 nsew signal input
rlabel metal3 s 119200 17824 120000 17944 6 wb_data_i[9]
port 192 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 wb_data_o[0]
port 193 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 wb_data_o[10]
port 194 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 wb_data_o[11]
port 195 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 wb_data_o[12]
port 196 nsew signal output
rlabel metal3 s 119200 21768 120000 21888 6 wb_data_o[13]
port 197 nsew signal output
rlabel metal3 s 119200 23128 120000 23248 6 wb_data_o[14]
port 198 nsew signal output
rlabel metal2 s 86406 39200 86462 40000 6 wb_data_o[15]
port 199 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 wb_data_o[16]
port 200 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 wb_data_o[17]
port 201 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 wb_data_o[18]
port 202 nsew signal output
rlabel metal2 s 100482 39200 100538 40000 6 wb_data_o[19]
port 203 nsew signal output
rlabel metal3 s 119200 8440 120000 8560 6 wb_data_o[1]
port 204 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 wb_data_o[20]
port 205 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 wb_data_o[21]
port 206 nsew signal output
rlabel metal3 s 119200 27208 120000 27328 6 wb_data_o[22]
port 207 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 wb_data_o[23]
port 208 nsew signal output
rlabel metal3 s 119200 31152 120000 31272 6 wb_data_o[24]
port 209 nsew signal output
rlabel metal2 s 114650 39200 114706 40000 6 wb_data_o[25]
port 210 nsew signal output
rlabel metal3 s 119200 32512 120000 32632 6 wb_data_o[26]
port 211 nsew signal output
rlabel metal3 s 119200 35096 120000 35216 6 wb_data_o[27]
port 212 nsew signal output
rlabel metal3 s 119200 37816 120000 37936 6 wb_data_o[28]
port 213 nsew signal output
rlabel metal3 s 119200 39176 120000 39296 6 wb_data_o[29]
port 214 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 wb_data_o[2]
port 215 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 wb_data_o[30]
port 216 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 wb_data_o[31]
port 217 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 wb_data_o[3]
port 218 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 wb_data_o[4]
port 219 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 wb_data_o[5]
port 220 nsew signal output
rlabel metal3 s 119200 13880 120000 14000 6 wb_data_o[6]
port 221 nsew signal output
rlabel metal2 s 68742 39200 68798 40000 6 wb_data_o[7]
port 222 nsew signal output
rlabel metal3 s 119200 16464 120000 16584 6 wb_data_o[8]
port 223 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 wb_data_o[9]
port 224 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 wb_error_o
port 225 nsew signal output
rlabel metal3 s 119200 1776 120000 1896 6 wb_rst_i
port 226 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 wb_sel_i[0]
port 227 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wb_sel_i[1]
port 228 nsew signal input
rlabel metal3 s 119200 11160 120000 11280 6 wb_sel_i[2]
port 229 nsew signal input
rlabel metal2 s 44086 39200 44142 40000 6 wb_sel_i[3]
port 230 nsew signal input
rlabel metal3 s 119200 3136 120000 3256 6 wb_stall_o
port 231 nsew signal output
rlabel metal3 s 119200 4496 120000 4616 6 wb_stb_i
port 232 nsew signal input
rlabel metal2 s 33506 39200 33562 40000 6 wb_we_i
port 233 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1817668
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Flash/runs/Flash/results/signoff/Flash.magic.gds
string GDS_START 176410
<< end >>

