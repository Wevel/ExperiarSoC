* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_sram_2kbyte_1rw1r_32x512_8 abstract view
.subckt sky130_sram_2kbyte_1rw1r_32x512_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr1[0]
+ addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] addr1[8] csb0 csb1
+ web0 clk0 clk1 wmask0[0] wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4]
+ dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13]
+ dout1[14] dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21]
+ dout1[22] dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29]
+ dout1[30] dout1[31] vccd1 vssd1
.ends

* Black-box entry subcircuit for Art abstract view
.subckt Art vccd1 vssd1
.ends

* Black-box entry subcircuit for ExperiarCore abstract view
.subckt ExperiarCore addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] addr0[8] addr1[0] addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6]
+ addr1[7] addr1[8] clk0 clk1 coreIndex[0] coreIndex[1] coreIndex[2] coreIndex[3]
+ coreIndex[4] coreIndex[5] coreIndex[6] coreIndex[7] core_wb_ack_i core_wb_adr_o[0]
+ core_wb_adr_o[10] core_wb_adr_o[11] core_wb_adr_o[12] core_wb_adr_o[13] core_wb_adr_o[14]
+ core_wb_adr_o[15] core_wb_adr_o[16] core_wb_adr_o[17] core_wb_adr_o[18] core_wb_adr_o[19]
+ core_wb_adr_o[1] core_wb_adr_o[20] core_wb_adr_o[21] core_wb_adr_o[22] core_wb_adr_o[23]
+ core_wb_adr_o[24] core_wb_adr_o[25] core_wb_adr_o[26] core_wb_adr_o[27] core_wb_adr_o[2]
+ core_wb_adr_o[3] core_wb_adr_o[4] core_wb_adr_o[5] core_wb_adr_o[6] core_wb_adr_o[7]
+ core_wb_adr_o[8] core_wb_adr_o[9] core_wb_cyc_o core_wb_data_i[0] core_wb_data_i[10]
+ core_wb_data_i[11] core_wb_data_i[12] core_wb_data_i[13] core_wb_data_i[14] core_wb_data_i[15]
+ core_wb_data_i[16] core_wb_data_i[17] core_wb_data_i[18] core_wb_data_i[19] core_wb_data_i[1]
+ core_wb_data_i[20] core_wb_data_i[21] core_wb_data_i[22] core_wb_data_i[23] core_wb_data_i[24]
+ core_wb_data_i[25] core_wb_data_i[26] core_wb_data_i[27] core_wb_data_i[28] core_wb_data_i[29]
+ core_wb_data_i[2] core_wb_data_i[30] core_wb_data_i[31] core_wb_data_i[3] core_wb_data_i[4]
+ core_wb_data_i[5] core_wb_data_i[6] core_wb_data_i[7] core_wb_data_i[8] core_wb_data_i[9]
+ core_wb_data_o[0] core_wb_data_o[10] core_wb_data_o[11] core_wb_data_o[12] core_wb_data_o[13]
+ core_wb_data_o[14] core_wb_data_o[15] core_wb_data_o[16] core_wb_data_o[17] core_wb_data_o[18]
+ core_wb_data_o[19] core_wb_data_o[1] core_wb_data_o[20] core_wb_data_o[21] core_wb_data_o[22]
+ core_wb_data_o[23] core_wb_data_o[24] core_wb_data_o[25] core_wb_data_o[26] core_wb_data_o[27]
+ core_wb_data_o[28] core_wb_data_o[29] core_wb_data_o[2] core_wb_data_o[30] core_wb_data_o[31]
+ core_wb_data_o[3] core_wb_data_o[4] core_wb_data_o[5] core_wb_data_o[6] core_wb_data_o[7]
+ core_wb_data_o[8] core_wb_data_o[9] core_wb_error_i core_wb_sel_o[0] core_wb_sel_o[1]
+ core_wb_sel_o[2] core_wb_sel_o[3] core_wb_stall_i core_wb_stb_o core_wb_we_o csb0[0]
+ csb0[1] csb1[0] csb1[1] din0[0] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[1] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[2] din0[30] din0[31]
+ din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] dout0[0] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[1] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[2] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35]
+ dout0[36] dout0[37] dout0[38] dout0[39] dout0[3] dout0[40] dout0[41] dout0[42] dout0[43]
+ dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[4] dout0[50] dout0[51]
+ dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59]
+ dout0[5] dout0[60] dout0[61] dout0[62] dout0[63] dout0[6] dout0[7] dout0[8] dout0[9]
+ dout1[0] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16] dout1[17]
+ dout1[18] dout1[19] dout1[1] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24] dout1[25]
+ dout1[26] dout1[27] dout1[28] dout1[29] dout1[2] dout1[30] dout1[31] dout1[32] dout1[33]
+ dout1[34] dout1[35] dout1[36] dout1[37] dout1[38] dout1[39] dout1[3] dout1[40] dout1[41]
+ dout1[42] dout1[43] dout1[44] dout1[45] dout1[46] dout1[47] dout1[48] dout1[49]
+ dout1[4] dout1[50] dout1[51] dout1[52] dout1[53] dout1[54] dout1[55] dout1[56] dout1[57]
+ dout1[58] dout1[59] dout1[5] dout1[60] dout1[61] dout1[62] dout1[63] dout1[6] dout1[7]
+ dout1[8] dout1[9] irq[0] irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[1]
+ irq[2] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] jtag_tck jtag_tdi jtag_tdo
+ jtag_tms localMemory_wb_ack_o localMemory_wb_adr_i[0] localMemory_wb_adr_i[10] localMemory_wb_adr_i[11]
+ localMemory_wb_adr_i[12] localMemory_wb_adr_i[13] localMemory_wb_adr_i[14] localMemory_wb_adr_i[15]
+ localMemory_wb_adr_i[16] localMemory_wb_adr_i[17] localMemory_wb_adr_i[18] localMemory_wb_adr_i[19]
+ localMemory_wb_adr_i[1] localMemory_wb_adr_i[20] localMemory_wb_adr_i[21] localMemory_wb_adr_i[22]
+ localMemory_wb_adr_i[23] localMemory_wb_adr_i[2] localMemory_wb_adr_i[3] localMemory_wb_adr_i[4]
+ localMemory_wb_adr_i[5] localMemory_wb_adr_i[6] localMemory_wb_adr_i[7] localMemory_wb_adr_i[8]
+ localMemory_wb_adr_i[9] localMemory_wb_cyc_i localMemory_wb_data_i[0] localMemory_wb_data_i[10]
+ localMemory_wb_data_i[11] localMemory_wb_data_i[12] localMemory_wb_data_i[13] localMemory_wb_data_i[14]
+ localMemory_wb_data_i[15] localMemory_wb_data_i[16] localMemory_wb_data_i[17] localMemory_wb_data_i[18]
+ localMemory_wb_data_i[19] localMemory_wb_data_i[1] localMemory_wb_data_i[20] localMemory_wb_data_i[21]
+ localMemory_wb_data_i[22] localMemory_wb_data_i[23] localMemory_wb_data_i[24] localMemory_wb_data_i[25]
+ localMemory_wb_data_i[26] localMemory_wb_data_i[27] localMemory_wb_data_i[28] localMemory_wb_data_i[29]
+ localMemory_wb_data_i[2] localMemory_wb_data_i[30] localMemory_wb_data_i[31] localMemory_wb_data_i[3]
+ localMemory_wb_data_i[4] localMemory_wb_data_i[5] localMemory_wb_data_i[6] localMemory_wb_data_i[7]
+ localMemory_wb_data_i[8] localMemory_wb_data_i[9] localMemory_wb_data_o[0] localMemory_wb_data_o[10]
+ localMemory_wb_data_o[11] localMemory_wb_data_o[12] localMemory_wb_data_o[13] localMemory_wb_data_o[14]
+ localMemory_wb_data_o[15] localMemory_wb_data_o[16] localMemory_wb_data_o[17] localMemory_wb_data_o[18]
+ localMemory_wb_data_o[19] localMemory_wb_data_o[1] localMemory_wb_data_o[20] localMemory_wb_data_o[21]
+ localMemory_wb_data_o[22] localMemory_wb_data_o[23] localMemory_wb_data_o[24] localMemory_wb_data_o[25]
+ localMemory_wb_data_o[26] localMemory_wb_data_o[27] localMemory_wb_data_o[28] localMemory_wb_data_o[29]
+ localMemory_wb_data_o[2] localMemory_wb_data_o[30] localMemory_wb_data_o[31] localMemory_wb_data_o[3]
+ localMemory_wb_data_o[4] localMemory_wb_data_o[5] localMemory_wb_data_o[6] localMemory_wb_data_o[7]
+ localMemory_wb_data_o[8] localMemory_wb_data_o[9] localMemory_wb_error_o localMemory_wb_sel_i[0]
+ localMemory_wb_sel_i[1] localMemory_wb_sel_i[2] localMemory_wb_sel_i[3] localMemory_wb_stall_o
+ localMemory_wb_stb_i localMemory_wb_we_i manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] probe_env[0] probe_env[1] probe_errorCode[0]
+ probe_errorCode[1] probe_isBranch probe_isCompressed probe_isLoad probe_isStore
+ probe_jtagInstruction[0] probe_jtagInstruction[1] probe_jtagInstruction[2] probe_jtagInstruction[3]
+ probe_jtagInstruction[4] probe_opcode[0] probe_opcode[1] probe_opcode[2] probe_opcode[3]
+ probe_opcode[4] probe_opcode[5] probe_opcode[6] probe_programCounter[0] probe_programCounter[10]
+ probe_programCounter[11] probe_programCounter[12] probe_programCounter[13] probe_programCounter[14]
+ probe_programCounter[15] probe_programCounter[16] probe_programCounter[17] probe_programCounter[18]
+ probe_programCounter[19] probe_programCounter[1] probe_programCounter[20] probe_programCounter[21]
+ probe_programCounter[22] probe_programCounter[23] probe_programCounter[24] probe_programCounter[25]
+ probe_programCounter[26] probe_programCounter[27] probe_programCounter[28] probe_programCounter[29]
+ probe_programCounter[2] probe_programCounter[30] probe_programCounter[31] probe_programCounter[3]
+ probe_programCounter[4] probe_programCounter[5] probe_programCounter[6] probe_programCounter[7]
+ probe_programCounter[8] probe_programCounter[9] probe_state[0] probe_state[1] probe_takeBranch
+ vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i
+ web0 wmask0[0] wmask0[1] wmask0[2] wmask0[3]
.ends

* Black-box entry subcircuit for Peripherals abstract view
.subckt Peripherals flash_csb flash_io0_read flash_io0_we flash_io0_write flash_io1_read
+ flash_io1_we flash_io1_write flash_sck internal_uart_rx internal_uart_tx io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] jtag_tck jtag_tdi jtag_tdo
+ jtag_tms peripheral_irq[0] peripheral_irq[1] peripheral_irq[2] peripheral_irq[3]
+ peripheral_irq[4] peripheral_irq[5] peripheral_irq[6] peripheral_irq[7] peripheral_irq[8]
+ peripheral_irq[9] probe_blink[0] probe_blink[1] vccd1 vga_b[0] vga_b[1] vga_g[0]
+ vga_g[1] vga_hsync vga_r[0] vga_r[1] vga_vsync vssd1 wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[2] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8]
+ wb_adr_i[9] wb_clk_i wb_cyc_i wb_data_i[0] wb_data_i[10] wb_data_i[11] wb_data_i[12]
+ wb_data_i[13] wb_data_i[14] wb_data_i[15] wb_data_i[16] wb_data_i[17] wb_data_i[18]
+ wb_data_i[19] wb_data_i[1] wb_data_i[20] wb_data_i[21] wb_data_i[22] wb_data_i[23]
+ wb_data_i[24] wb_data_i[25] wb_data_i[26] wb_data_i[27] wb_data_i[28] wb_data_i[29]
+ wb_data_i[2] wb_data_i[30] wb_data_i[31] wb_data_i[3] wb_data_i[4] wb_data_i[5]
+ wb_data_i[6] wb_data_i[7] wb_data_i[8] wb_data_i[9] wb_data_o[0] wb_data_o[10] wb_data_o[11]
+ wb_data_o[12] wb_data_o[13] wb_data_o[14] wb_data_o[15] wb_data_o[16] wb_data_o[17]
+ wb_data_o[18] wb_data_o[19] wb_data_o[1] wb_data_o[20] wb_data_o[21] wb_data_o[22]
+ wb_data_o[23] wb_data_o[24] wb_data_o[25] wb_data_o[26] wb_data_o[27] wb_data_o[28]
+ wb_data_o[29] wb_data_o[2] wb_data_o[30] wb_data_o[31] wb_data_o[3] wb_data_o[4]
+ wb_data_o[5] wb_data_o[6] wb_data_o[7] wb_data_o[8] wb_data_o[9] wb_error_o wb_rst_i
+ wb_sel_i[0] wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stall_o wb_stb_i wb_we_i
.ends

* Black-box entry subcircuit for WishboneInterconnect abstract view
.subckt WishboneInterconnect master0_wb_ack_i master0_wb_adr_o[0] master0_wb_adr_o[10]
+ master0_wb_adr_o[11] master0_wb_adr_o[12] master0_wb_adr_o[13] master0_wb_adr_o[14]
+ master0_wb_adr_o[15] master0_wb_adr_o[16] master0_wb_adr_o[17] master0_wb_adr_o[18]
+ master0_wb_adr_o[19] master0_wb_adr_o[1] master0_wb_adr_o[20] master0_wb_adr_o[21]
+ master0_wb_adr_o[22] master0_wb_adr_o[23] master0_wb_adr_o[24] master0_wb_adr_o[25]
+ master0_wb_adr_o[26] master0_wb_adr_o[27] master0_wb_adr_o[2] master0_wb_adr_o[3]
+ master0_wb_adr_o[4] master0_wb_adr_o[5] master0_wb_adr_o[6] master0_wb_adr_o[7]
+ master0_wb_adr_o[8] master0_wb_adr_o[9] master0_wb_cyc_o master0_wb_data_i[0] master0_wb_data_i[10]
+ master0_wb_data_i[11] master0_wb_data_i[12] master0_wb_data_i[13] master0_wb_data_i[14]
+ master0_wb_data_i[15] master0_wb_data_i[16] master0_wb_data_i[17] master0_wb_data_i[18]
+ master0_wb_data_i[19] master0_wb_data_i[1] master0_wb_data_i[20] master0_wb_data_i[21]
+ master0_wb_data_i[22] master0_wb_data_i[23] master0_wb_data_i[24] master0_wb_data_i[25]
+ master0_wb_data_i[26] master0_wb_data_i[27] master0_wb_data_i[28] master0_wb_data_i[29]
+ master0_wb_data_i[2] master0_wb_data_i[30] master0_wb_data_i[31] master0_wb_data_i[3]
+ master0_wb_data_i[4] master0_wb_data_i[5] master0_wb_data_i[6] master0_wb_data_i[7]
+ master0_wb_data_i[8] master0_wb_data_i[9] master0_wb_data_o[0] master0_wb_data_o[10]
+ master0_wb_data_o[11] master0_wb_data_o[12] master0_wb_data_o[13] master0_wb_data_o[14]
+ master0_wb_data_o[15] master0_wb_data_o[16] master0_wb_data_o[17] master0_wb_data_o[18]
+ master0_wb_data_o[19] master0_wb_data_o[1] master0_wb_data_o[20] master0_wb_data_o[21]
+ master0_wb_data_o[22] master0_wb_data_o[23] master0_wb_data_o[24] master0_wb_data_o[25]
+ master0_wb_data_o[26] master0_wb_data_o[27] master0_wb_data_o[28] master0_wb_data_o[29]
+ master0_wb_data_o[2] master0_wb_data_o[30] master0_wb_data_o[31] master0_wb_data_o[3]
+ master0_wb_data_o[4] master0_wb_data_o[5] master0_wb_data_o[6] master0_wb_data_o[7]
+ master0_wb_data_o[8] master0_wb_data_o[9] master0_wb_error_i master0_wb_sel_o[0]
+ master0_wb_sel_o[1] master0_wb_sel_o[2] master0_wb_sel_o[3] master0_wb_stall_i master0_wb_stb_o
+ master0_wb_we_o master1_wb_ack_i master1_wb_adr_o[0] master1_wb_adr_o[10] master1_wb_adr_o[11]
+ master1_wb_adr_o[12] master1_wb_adr_o[13] master1_wb_adr_o[14] master1_wb_adr_o[15]
+ master1_wb_adr_o[16] master1_wb_adr_o[17] master1_wb_adr_o[18] master1_wb_adr_o[19]
+ master1_wb_adr_o[1] master1_wb_adr_o[20] master1_wb_adr_o[21] master1_wb_adr_o[22]
+ master1_wb_adr_o[23] master1_wb_adr_o[24] master1_wb_adr_o[25] master1_wb_adr_o[26]
+ master1_wb_adr_o[27] master1_wb_adr_o[2] master1_wb_adr_o[3] master1_wb_adr_o[4]
+ master1_wb_adr_o[5] master1_wb_adr_o[6] master1_wb_adr_o[7] master1_wb_adr_o[8]
+ master1_wb_adr_o[9] master1_wb_cyc_o master1_wb_data_i[0] master1_wb_data_i[10]
+ master1_wb_data_i[11] master1_wb_data_i[12] master1_wb_data_i[13] master1_wb_data_i[14]
+ master1_wb_data_i[15] master1_wb_data_i[16] master1_wb_data_i[17] master1_wb_data_i[18]
+ master1_wb_data_i[19] master1_wb_data_i[1] master1_wb_data_i[20] master1_wb_data_i[21]
+ master1_wb_data_i[22] master1_wb_data_i[23] master1_wb_data_i[24] master1_wb_data_i[25]
+ master1_wb_data_i[26] master1_wb_data_i[27] master1_wb_data_i[28] master1_wb_data_i[29]
+ master1_wb_data_i[2] master1_wb_data_i[30] master1_wb_data_i[31] master1_wb_data_i[3]
+ master1_wb_data_i[4] master1_wb_data_i[5] master1_wb_data_i[6] master1_wb_data_i[7]
+ master1_wb_data_i[8] master1_wb_data_i[9] master1_wb_data_o[0] master1_wb_data_o[10]
+ master1_wb_data_o[11] master1_wb_data_o[12] master1_wb_data_o[13] master1_wb_data_o[14]
+ master1_wb_data_o[15] master1_wb_data_o[16] master1_wb_data_o[17] master1_wb_data_o[18]
+ master1_wb_data_o[19] master1_wb_data_o[1] master1_wb_data_o[20] master1_wb_data_o[21]
+ master1_wb_data_o[22] master1_wb_data_o[23] master1_wb_data_o[24] master1_wb_data_o[25]
+ master1_wb_data_o[26] master1_wb_data_o[27] master1_wb_data_o[28] master1_wb_data_o[29]
+ master1_wb_data_o[2] master1_wb_data_o[30] master1_wb_data_o[31] master1_wb_data_o[3]
+ master1_wb_data_o[4] master1_wb_data_o[5] master1_wb_data_o[6] master1_wb_data_o[7]
+ master1_wb_data_o[8] master1_wb_data_o[9] master1_wb_error_i master1_wb_sel_o[0]
+ master1_wb_sel_o[1] master1_wb_sel_o[2] master1_wb_sel_o[3] master1_wb_stall_i master1_wb_stb_o
+ master1_wb_we_o master2_wb_ack_i master2_wb_adr_o[0] master2_wb_adr_o[10] master2_wb_adr_o[11]
+ master2_wb_adr_o[12] master2_wb_adr_o[13] master2_wb_adr_o[14] master2_wb_adr_o[15]
+ master2_wb_adr_o[16] master2_wb_adr_o[17] master2_wb_adr_o[18] master2_wb_adr_o[19]
+ master2_wb_adr_o[1] master2_wb_adr_o[20] master2_wb_adr_o[21] master2_wb_adr_o[22]
+ master2_wb_adr_o[23] master2_wb_adr_o[24] master2_wb_adr_o[25] master2_wb_adr_o[26]
+ master2_wb_adr_o[27] master2_wb_adr_o[2] master2_wb_adr_o[3] master2_wb_adr_o[4]
+ master2_wb_adr_o[5] master2_wb_adr_o[6] master2_wb_adr_o[7] master2_wb_adr_o[8]
+ master2_wb_adr_o[9] master2_wb_cyc_o master2_wb_data_i[0] master2_wb_data_i[10]
+ master2_wb_data_i[11] master2_wb_data_i[12] master2_wb_data_i[13] master2_wb_data_i[14]
+ master2_wb_data_i[15] master2_wb_data_i[16] master2_wb_data_i[17] master2_wb_data_i[18]
+ master2_wb_data_i[19] master2_wb_data_i[1] master2_wb_data_i[20] master2_wb_data_i[21]
+ master2_wb_data_i[22] master2_wb_data_i[23] master2_wb_data_i[24] master2_wb_data_i[25]
+ master2_wb_data_i[26] master2_wb_data_i[27] master2_wb_data_i[28] master2_wb_data_i[29]
+ master2_wb_data_i[2] master2_wb_data_i[30] master2_wb_data_i[31] master2_wb_data_i[3]
+ master2_wb_data_i[4] master2_wb_data_i[5] master2_wb_data_i[6] master2_wb_data_i[7]
+ master2_wb_data_i[8] master2_wb_data_i[9] master2_wb_data_o[0] master2_wb_data_o[10]
+ master2_wb_data_o[11] master2_wb_data_o[12] master2_wb_data_o[13] master2_wb_data_o[14]
+ master2_wb_data_o[15] master2_wb_data_o[16] master2_wb_data_o[17] master2_wb_data_o[18]
+ master2_wb_data_o[19] master2_wb_data_o[1] master2_wb_data_o[20] master2_wb_data_o[21]
+ master2_wb_data_o[22] master2_wb_data_o[23] master2_wb_data_o[24] master2_wb_data_o[25]
+ master2_wb_data_o[26] master2_wb_data_o[27] master2_wb_data_o[28] master2_wb_data_o[29]
+ master2_wb_data_o[2] master2_wb_data_o[30] master2_wb_data_o[31] master2_wb_data_o[3]
+ master2_wb_data_o[4] master2_wb_data_o[5] master2_wb_data_o[6] master2_wb_data_o[7]
+ master2_wb_data_o[8] master2_wb_data_o[9] master2_wb_error_i master2_wb_sel_o[0]
+ master2_wb_sel_o[1] master2_wb_sel_o[2] master2_wb_sel_o[3] master2_wb_stall_i master2_wb_stb_o
+ master2_wb_we_o probe_master0_currentSlave[0] probe_master0_currentSlave[1] probe_master1_currentSlave[0]
+ probe_master1_currentSlave[1] probe_master2_currentSlave[0] probe_master2_currentSlave[1]
+ probe_master3_currentSlave[0] probe_master3_currentSlave[1] probe_slave0_currentMaster[0]
+ probe_slave0_currentMaster[1] probe_slave1_currentMaster[0] probe_slave1_currentMaster[1]
+ probe_slave2_currentMaster[0] probe_slave2_currentMaster[1] probe_slave3_currentMaster[0]
+ probe_slave3_currentMaster[1] slave0_wb_ack_o slave0_wb_adr_i[0] slave0_wb_adr_i[10]
+ slave0_wb_adr_i[11] slave0_wb_adr_i[12] slave0_wb_adr_i[13] slave0_wb_adr_i[14]
+ slave0_wb_adr_i[15] slave0_wb_adr_i[16] slave0_wb_adr_i[17] slave0_wb_adr_i[18]
+ slave0_wb_adr_i[19] slave0_wb_adr_i[1] slave0_wb_adr_i[20] slave0_wb_adr_i[21] slave0_wb_adr_i[22]
+ slave0_wb_adr_i[23] slave0_wb_adr_i[2] slave0_wb_adr_i[3] slave0_wb_adr_i[4] slave0_wb_adr_i[5]
+ slave0_wb_adr_i[6] slave0_wb_adr_i[7] slave0_wb_adr_i[8] slave0_wb_adr_i[9] slave0_wb_cyc_i
+ slave0_wb_data_i[0] slave0_wb_data_i[10] slave0_wb_data_i[11] slave0_wb_data_i[12]
+ slave0_wb_data_i[13] slave0_wb_data_i[14] slave0_wb_data_i[15] slave0_wb_data_i[16]
+ slave0_wb_data_i[17] slave0_wb_data_i[18] slave0_wb_data_i[19] slave0_wb_data_i[1]
+ slave0_wb_data_i[20] slave0_wb_data_i[21] slave0_wb_data_i[22] slave0_wb_data_i[23]
+ slave0_wb_data_i[24] slave0_wb_data_i[25] slave0_wb_data_i[26] slave0_wb_data_i[27]
+ slave0_wb_data_i[28] slave0_wb_data_i[29] slave0_wb_data_i[2] slave0_wb_data_i[30]
+ slave0_wb_data_i[31] slave0_wb_data_i[3] slave0_wb_data_i[4] slave0_wb_data_i[5]
+ slave0_wb_data_i[6] slave0_wb_data_i[7] slave0_wb_data_i[8] slave0_wb_data_i[9]
+ slave0_wb_data_o[0] slave0_wb_data_o[10] slave0_wb_data_o[11] slave0_wb_data_o[12]
+ slave0_wb_data_o[13] slave0_wb_data_o[14] slave0_wb_data_o[15] slave0_wb_data_o[16]
+ slave0_wb_data_o[17] slave0_wb_data_o[18] slave0_wb_data_o[19] slave0_wb_data_o[1]
+ slave0_wb_data_o[20] slave0_wb_data_o[21] slave0_wb_data_o[22] slave0_wb_data_o[23]
+ slave0_wb_data_o[24] slave0_wb_data_o[25] slave0_wb_data_o[26] slave0_wb_data_o[27]
+ slave0_wb_data_o[28] slave0_wb_data_o[29] slave0_wb_data_o[2] slave0_wb_data_o[30]
+ slave0_wb_data_o[31] slave0_wb_data_o[3] slave0_wb_data_o[4] slave0_wb_data_o[5]
+ slave0_wb_data_o[6] slave0_wb_data_o[7] slave0_wb_data_o[8] slave0_wb_data_o[9]
+ slave0_wb_error_o slave0_wb_sel_i[0] slave0_wb_sel_i[1] slave0_wb_sel_i[2] slave0_wb_sel_i[3]
+ slave0_wb_stall_o slave0_wb_stb_i slave0_wb_we_i slave1_wb_ack_o slave1_wb_adr_i[0]
+ slave1_wb_adr_i[10] slave1_wb_adr_i[11] slave1_wb_adr_i[12] slave1_wb_adr_i[13]
+ slave1_wb_adr_i[14] slave1_wb_adr_i[15] slave1_wb_adr_i[16] slave1_wb_adr_i[17]
+ slave1_wb_adr_i[18] slave1_wb_adr_i[19] slave1_wb_adr_i[1] slave1_wb_adr_i[20] slave1_wb_adr_i[21]
+ slave1_wb_adr_i[22] slave1_wb_adr_i[23] slave1_wb_adr_i[2] slave1_wb_adr_i[3] slave1_wb_adr_i[4]
+ slave1_wb_adr_i[5] slave1_wb_adr_i[6] slave1_wb_adr_i[7] slave1_wb_adr_i[8] slave1_wb_adr_i[9]
+ slave1_wb_cyc_i slave1_wb_data_i[0] slave1_wb_data_i[10] slave1_wb_data_i[11] slave1_wb_data_i[12]
+ slave1_wb_data_i[13] slave1_wb_data_i[14] slave1_wb_data_i[15] slave1_wb_data_i[16]
+ slave1_wb_data_i[17] slave1_wb_data_i[18] slave1_wb_data_i[19] slave1_wb_data_i[1]
+ slave1_wb_data_i[20] slave1_wb_data_i[21] slave1_wb_data_i[22] slave1_wb_data_i[23]
+ slave1_wb_data_i[24] slave1_wb_data_i[25] slave1_wb_data_i[26] slave1_wb_data_i[27]
+ slave1_wb_data_i[28] slave1_wb_data_i[29] slave1_wb_data_i[2] slave1_wb_data_i[30]
+ slave1_wb_data_i[31] slave1_wb_data_i[3] slave1_wb_data_i[4] slave1_wb_data_i[5]
+ slave1_wb_data_i[6] slave1_wb_data_i[7] slave1_wb_data_i[8] slave1_wb_data_i[9]
+ slave1_wb_data_o[0] slave1_wb_data_o[10] slave1_wb_data_o[11] slave1_wb_data_o[12]
+ slave1_wb_data_o[13] slave1_wb_data_o[14] slave1_wb_data_o[15] slave1_wb_data_o[16]
+ slave1_wb_data_o[17] slave1_wb_data_o[18] slave1_wb_data_o[19] slave1_wb_data_o[1]
+ slave1_wb_data_o[20] slave1_wb_data_o[21] slave1_wb_data_o[22] slave1_wb_data_o[23]
+ slave1_wb_data_o[24] slave1_wb_data_o[25] slave1_wb_data_o[26] slave1_wb_data_o[27]
+ slave1_wb_data_o[28] slave1_wb_data_o[29] slave1_wb_data_o[2] slave1_wb_data_o[30]
+ slave1_wb_data_o[31] slave1_wb_data_o[3] slave1_wb_data_o[4] slave1_wb_data_o[5]
+ slave1_wb_data_o[6] slave1_wb_data_o[7] slave1_wb_data_o[8] slave1_wb_data_o[9]
+ slave1_wb_error_o slave1_wb_sel_i[0] slave1_wb_sel_i[1] slave1_wb_sel_i[2] slave1_wb_sel_i[3]
+ slave1_wb_stall_o slave1_wb_stb_i slave1_wb_we_i slave2_wb_ack_o slave2_wb_adr_i[0]
+ slave2_wb_adr_i[10] slave2_wb_adr_i[11] slave2_wb_adr_i[12] slave2_wb_adr_i[13]
+ slave2_wb_adr_i[14] slave2_wb_adr_i[15] slave2_wb_adr_i[16] slave2_wb_adr_i[17]
+ slave2_wb_adr_i[18] slave2_wb_adr_i[19] slave2_wb_adr_i[1] slave2_wb_adr_i[20] slave2_wb_adr_i[21]
+ slave2_wb_adr_i[22] slave2_wb_adr_i[23] slave2_wb_adr_i[2] slave2_wb_adr_i[3] slave2_wb_adr_i[4]
+ slave2_wb_adr_i[5] slave2_wb_adr_i[6] slave2_wb_adr_i[7] slave2_wb_adr_i[8] slave2_wb_adr_i[9]
+ slave2_wb_cyc_i slave2_wb_data_i[0] slave2_wb_data_i[10] slave2_wb_data_i[11] slave2_wb_data_i[12]
+ slave2_wb_data_i[13] slave2_wb_data_i[14] slave2_wb_data_i[15] slave2_wb_data_i[16]
+ slave2_wb_data_i[17] slave2_wb_data_i[18] slave2_wb_data_i[19] slave2_wb_data_i[1]
+ slave2_wb_data_i[20] slave2_wb_data_i[21] slave2_wb_data_i[22] slave2_wb_data_i[23]
+ slave2_wb_data_i[24] slave2_wb_data_i[25] slave2_wb_data_i[26] slave2_wb_data_i[27]
+ slave2_wb_data_i[28] slave2_wb_data_i[29] slave2_wb_data_i[2] slave2_wb_data_i[30]
+ slave2_wb_data_i[31] slave2_wb_data_i[3] slave2_wb_data_i[4] slave2_wb_data_i[5]
+ slave2_wb_data_i[6] slave2_wb_data_i[7] slave2_wb_data_i[8] slave2_wb_data_i[9]
+ slave2_wb_data_o[0] slave2_wb_data_o[10] slave2_wb_data_o[11] slave2_wb_data_o[12]
+ slave2_wb_data_o[13] slave2_wb_data_o[14] slave2_wb_data_o[15] slave2_wb_data_o[16]
+ slave2_wb_data_o[17] slave2_wb_data_o[18] slave2_wb_data_o[19] slave2_wb_data_o[1]
+ slave2_wb_data_o[20] slave2_wb_data_o[21] slave2_wb_data_o[22] slave2_wb_data_o[23]
+ slave2_wb_data_o[24] slave2_wb_data_o[25] slave2_wb_data_o[26] slave2_wb_data_o[27]
+ slave2_wb_data_o[28] slave2_wb_data_o[29] slave2_wb_data_o[2] slave2_wb_data_o[30]
+ slave2_wb_data_o[31] slave2_wb_data_o[3] slave2_wb_data_o[4] slave2_wb_data_o[5]
+ slave2_wb_data_o[6] slave2_wb_data_o[7] slave2_wb_data_o[8] slave2_wb_data_o[9]
+ slave2_wb_error_o slave2_wb_sel_i[0] slave2_wb_sel_i[1] slave2_wb_sel_i[2] slave2_wb_sel_i[3]
+ slave2_wb_stall_o slave2_wb_stb_i slave2_wb_we_i slave3_wb_ack_o slave3_wb_adr_i[0]
+ slave3_wb_adr_i[10] slave3_wb_adr_i[11] slave3_wb_adr_i[12] slave3_wb_adr_i[13]
+ slave3_wb_adr_i[14] slave3_wb_adr_i[15] slave3_wb_adr_i[16] slave3_wb_adr_i[17]
+ slave3_wb_adr_i[18] slave3_wb_adr_i[19] slave3_wb_adr_i[1] slave3_wb_adr_i[20] slave3_wb_adr_i[21]
+ slave3_wb_adr_i[22] slave3_wb_adr_i[23] slave3_wb_adr_i[2] slave3_wb_adr_i[3] slave3_wb_adr_i[4]
+ slave3_wb_adr_i[5] slave3_wb_adr_i[6] slave3_wb_adr_i[7] slave3_wb_adr_i[8] slave3_wb_adr_i[9]
+ slave3_wb_cyc_i slave3_wb_data_i[0] slave3_wb_data_i[10] slave3_wb_data_i[11] slave3_wb_data_i[12]
+ slave3_wb_data_i[13] slave3_wb_data_i[14] slave3_wb_data_i[15] slave3_wb_data_i[16]
+ slave3_wb_data_i[17] slave3_wb_data_i[18] slave3_wb_data_i[19] slave3_wb_data_i[1]
+ slave3_wb_data_i[20] slave3_wb_data_i[21] slave3_wb_data_i[22] slave3_wb_data_i[23]
+ slave3_wb_data_i[24] slave3_wb_data_i[25] slave3_wb_data_i[26] slave3_wb_data_i[27]
+ slave3_wb_data_i[28] slave3_wb_data_i[29] slave3_wb_data_i[2] slave3_wb_data_i[30]
+ slave3_wb_data_i[31] slave3_wb_data_i[3] slave3_wb_data_i[4] slave3_wb_data_i[5]
+ slave3_wb_data_i[6] slave3_wb_data_i[7] slave3_wb_data_i[8] slave3_wb_data_i[9]
+ slave3_wb_data_o[0] slave3_wb_data_o[10] slave3_wb_data_o[11] slave3_wb_data_o[12]
+ slave3_wb_data_o[13] slave3_wb_data_o[14] slave3_wb_data_o[15] slave3_wb_data_o[16]
+ slave3_wb_data_o[17] slave3_wb_data_o[18] slave3_wb_data_o[19] slave3_wb_data_o[1]
+ slave3_wb_data_o[20] slave3_wb_data_o[21] slave3_wb_data_o[22] slave3_wb_data_o[23]
+ slave3_wb_data_o[24] slave3_wb_data_o[25] slave3_wb_data_o[26] slave3_wb_data_o[27]
+ slave3_wb_data_o[28] slave3_wb_data_o[29] slave3_wb_data_o[2] slave3_wb_data_o[30]
+ slave3_wb_data_o[31] slave3_wb_data_o[3] slave3_wb_data_o[4] slave3_wb_data_o[5]
+ slave3_wb_data_o[6] slave3_wb_data_o[7] slave3_wb_data_o[8] slave3_wb_data_o[9]
+ slave3_wb_error_o slave3_wb_sel_i[0] slave3_wb_sel_i[1] slave3_wb_sel_i[2] slave3_wb_sel_i[3]
+ slave3_wb_stall_o slave3_wb_stb_i slave3_wb_we_i slave4_wb_ack_o slave4_wb_adr_i[0]
+ slave4_wb_adr_i[10] slave4_wb_adr_i[11] slave4_wb_adr_i[12] slave4_wb_adr_i[13]
+ slave4_wb_adr_i[14] slave4_wb_adr_i[15] slave4_wb_adr_i[16] slave4_wb_adr_i[17]
+ slave4_wb_adr_i[18] slave4_wb_adr_i[19] slave4_wb_adr_i[1] slave4_wb_adr_i[20] slave4_wb_adr_i[21]
+ slave4_wb_adr_i[22] slave4_wb_adr_i[23] slave4_wb_adr_i[2] slave4_wb_adr_i[3] slave4_wb_adr_i[4]
+ slave4_wb_adr_i[5] slave4_wb_adr_i[6] slave4_wb_adr_i[7] slave4_wb_adr_i[8] slave4_wb_adr_i[9]
+ slave4_wb_cyc_i slave4_wb_data_i[0] slave4_wb_data_i[10] slave4_wb_data_i[11] slave4_wb_data_i[12]
+ slave4_wb_data_i[13] slave4_wb_data_i[14] slave4_wb_data_i[15] slave4_wb_data_i[16]
+ slave4_wb_data_i[17] slave4_wb_data_i[18] slave4_wb_data_i[19] slave4_wb_data_i[1]
+ slave4_wb_data_i[20] slave4_wb_data_i[21] slave4_wb_data_i[22] slave4_wb_data_i[23]
+ slave4_wb_data_i[24] slave4_wb_data_i[25] slave4_wb_data_i[26] slave4_wb_data_i[27]
+ slave4_wb_data_i[28] slave4_wb_data_i[29] slave4_wb_data_i[2] slave4_wb_data_i[30]
+ slave4_wb_data_i[31] slave4_wb_data_i[3] slave4_wb_data_i[4] slave4_wb_data_i[5]
+ slave4_wb_data_i[6] slave4_wb_data_i[7] slave4_wb_data_i[8] slave4_wb_data_i[9]
+ slave4_wb_data_o[0] slave4_wb_data_o[10] slave4_wb_data_o[11] slave4_wb_data_o[12]
+ slave4_wb_data_o[13] slave4_wb_data_o[14] slave4_wb_data_o[15] slave4_wb_data_o[16]
+ slave4_wb_data_o[17] slave4_wb_data_o[18] slave4_wb_data_o[19] slave4_wb_data_o[1]
+ slave4_wb_data_o[20] slave4_wb_data_o[21] slave4_wb_data_o[22] slave4_wb_data_o[23]
+ slave4_wb_data_o[24] slave4_wb_data_o[25] slave4_wb_data_o[26] slave4_wb_data_o[27]
+ slave4_wb_data_o[28] slave4_wb_data_o[29] slave4_wb_data_o[2] slave4_wb_data_o[30]
+ slave4_wb_data_o[31] slave4_wb_data_o[3] slave4_wb_data_o[4] slave4_wb_data_o[5]
+ slave4_wb_data_o[6] slave4_wb_data_o[7] slave4_wb_data_o[8] slave4_wb_data_o[9]
+ slave4_wb_error_o slave4_wb_sel_i[0] slave4_wb_sel_i[1] slave4_wb_sel_i[2] slave4_wb_sel_i[3]
+ slave4_wb_stall_o slave4_wb_stb_i slave4_wb_we_i vccd1 vssd1 wb_clk_i wb_rst_i
.ends

* Black-box entry subcircuit for CaravelHost abstract view
.subckt CaravelHost caravel_irq[0] caravel_irq[1] caravel_irq[2] caravel_irq[3] caravel_uart_rx
+ caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0] caravel_wb_adr_o[10] caravel_wb_adr_o[11]
+ caravel_wb_adr_o[12] caravel_wb_adr_o[13] caravel_wb_adr_o[14] caravel_wb_adr_o[15]
+ caravel_wb_adr_o[16] caravel_wb_adr_o[17] caravel_wb_adr_o[18] caravel_wb_adr_o[19]
+ caravel_wb_adr_o[1] caravel_wb_adr_o[20] caravel_wb_adr_o[21] caravel_wb_adr_o[22]
+ caravel_wb_adr_o[23] caravel_wb_adr_o[24] caravel_wb_adr_o[25] caravel_wb_adr_o[26]
+ caravel_wb_adr_o[27] caravel_wb_adr_o[2] caravel_wb_adr_o[3] caravel_wb_adr_o[4]
+ caravel_wb_adr_o[5] caravel_wb_adr_o[6] caravel_wb_adr_o[7] caravel_wb_adr_o[8]
+ caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0] caravel_wb_data_i[10]
+ caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13] caravel_wb_data_i[14]
+ caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17] caravel_wb_data_i[18]
+ caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20] caravel_wb_data_i[21]
+ caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24] caravel_wb_data_i[25]
+ caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28] caravel_wb_data_i[29]
+ caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31] caravel_wb_data_i[3]
+ caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6] caravel_wb_data_i[7]
+ caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0] caravel_wb_data_o[10]
+ caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13] caravel_wb_data_o[14]
+ caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17] caravel_wb_data_o[18]
+ caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20] caravel_wb_data_o[21]
+ caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24] caravel_wb_data_o[25]
+ caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28] caravel_wb_data_o[29]
+ caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31] caravel_wb_data_o[3]
+ caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6] caravel_wb_data_o[7]
+ caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i caravel_wb_sel_o[0]
+ caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3] caravel_wb_stall_i caravel_wb_stb_o
+ caravel_wb_we_o core0Index[0] core0Index[1] core0Index[2] core0Index[3] core0Index[4]
+ core0Index[5] core0Index[6] core0Index[7] core1Index[0] core1Index[1] core1Index[2]
+ core1Index[3] core1Index[4] core1Index[5] core1Index[6] core1Index[7] manufacturerID[0]
+ manufacturerID[10] manufacturerID[1] manufacturerID[2] manufacturerID[3] manufacturerID[4]
+ manufacturerID[5] manufacturerID[6] manufacturerID[7] manufacturerID[8] manufacturerID[9]
+ partID[0] partID[10] partID[11] partID[12] partID[13] partID[14] partID[15] partID[1]
+ partID[2] partID[3] partID[4] partID[5] partID[6] partID[7] partID[8] partID[9]
+ vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12]
+ wbs_data_i[13] wbs_data_i[14] wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18]
+ wbs_data_i[19] wbs_data_i[1] wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23]
+ wbs_data_i[24] wbs_data_i[25] wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29]
+ wbs_data_i[2] wbs_data_i[30] wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5]
+ wbs_data_i[6] wbs_data_i[7] wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10]
+ wbs_data_o[11] wbs_data_o[12] wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16]
+ wbs_data_o[17] wbs_data_o[18] wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21]
+ wbs_data_o[22] wbs_data_o[23] wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27]
+ wbs_data_o[28] wbs_data_o[29] wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3]
+ wbs_data_o[4] wbs_data_o[5] wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for Video abstract view
.subckt Video sram0_addr0[0] sram0_addr0[1] sram0_addr0[2] sram0_addr0[3] sram0_addr0[4]
+ sram0_addr0[5] sram0_addr0[6] sram0_addr0[7] sram0_addr0[8] sram0_addr1[0] sram0_addr1[1]
+ sram0_addr1[2] sram0_addr1[3] sram0_addr1[4] sram0_addr1[5] sram0_addr1[6] sram0_addr1[7]
+ sram0_addr1[8] sram0_clk0 sram0_clk1 sram0_csb0[0] sram0_csb0[1] sram0_csb1[0] sram0_csb1[1]
+ sram0_din0[0] sram0_din0[10] sram0_din0[11] sram0_din0[12] sram0_din0[13] sram0_din0[14]
+ sram0_din0[15] sram0_din0[16] sram0_din0[17] sram0_din0[18] sram0_din0[19] sram0_din0[1]
+ sram0_din0[20] sram0_din0[21] sram0_din0[22] sram0_din0[23] sram0_din0[24] sram0_din0[25]
+ sram0_din0[26] sram0_din0[27] sram0_din0[28] sram0_din0[29] sram0_din0[2] sram0_din0[30]
+ sram0_din0[31] sram0_din0[3] sram0_din0[4] sram0_din0[5] sram0_din0[6] sram0_din0[7]
+ sram0_din0[8] sram0_din0[9] sram0_dout0[0] sram0_dout0[10] sram0_dout0[11] sram0_dout0[12]
+ sram0_dout0[13] sram0_dout0[14] sram0_dout0[15] sram0_dout0[16] sram0_dout0[17]
+ sram0_dout0[18] sram0_dout0[19] sram0_dout0[1] sram0_dout0[20] sram0_dout0[21] sram0_dout0[22]
+ sram0_dout0[23] sram0_dout0[24] sram0_dout0[25] sram0_dout0[26] sram0_dout0[27]
+ sram0_dout0[28] sram0_dout0[29] sram0_dout0[2] sram0_dout0[30] sram0_dout0[31] sram0_dout0[32]
+ sram0_dout0[33] sram0_dout0[34] sram0_dout0[35] sram0_dout0[36] sram0_dout0[37]
+ sram0_dout0[38] sram0_dout0[39] sram0_dout0[3] sram0_dout0[40] sram0_dout0[41] sram0_dout0[42]
+ sram0_dout0[43] sram0_dout0[44] sram0_dout0[45] sram0_dout0[46] sram0_dout0[47]
+ sram0_dout0[48] sram0_dout0[49] sram0_dout0[4] sram0_dout0[50] sram0_dout0[51] sram0_dout0[52]
+ sram0_dout0[53] sram0_dout0[54] sram0_dout0[55] sram0_dout0[56] sram0_dout0[57]
+ sram0_dout0[58] sram0_dout0[59] sram0_dout0[5] sram0_dout0[60] sram0_dout0[61] sram0_dout0[62]
+ sram0_dout0[63] sram0_dout0[6] sram0_dout0[7] sram0_dout0[8] sram0_dout0[9] sram0_dout1[0]
+ sram0_dout1[10] sram0_dout1[11] sram0_dout1[12] sram0_dout1[13] sram0_dout1[14]
+ sram0_dout1[15] sram0_dout1[16] sram0_dout1[17] sram0_dout1[18] sram0_dout1[19]
+ sram0_dout1[1] sram0_dout1[20] sram0_dout1[21] sram0_dout1[22] sram0_dout1[23] sram0_dout1[24]
+ sram0_dout1[25] sram0_dout1[26] sram0_dout1[27] sram0_dout1[28] sram0_dout1[29]
+ sram0_dout1[2] sram0_dout1[30] sram0_dout1[31] sram0_dout1[32] sram0_dout1[33] sram0_dout1[34]
+ sram0_dout1[35] sram0_dout1[36] sram0_dout1[37] sram0_dout1[38] sram0_dout1[39]
+ sram0_dout1[3] sram0_dout1[40] sram0_dout1[41] sram0_dout1[42] sram0_dout1[43] sram0_dout1[44]
+ sram0_dout1[45] sram0_dout1[46] sram0_dout1[47] sram0_dout1[48] sram0_dout1[49]
+ sram0_dout1[4] sram0_dout1[50] sram0_dout1[51] sram0_dout1[52] sram0_dout1[53] sram0_dout1[54]
+ sram0_dout1[55] sram0_dout1[56] sram0_dout1[57] sram0_dout1[58] sram0_dout1[59]
+ sram0_dout1[5] sram0_dout1[60] sram0_dout1[61] sram0_dout1[62] sram0_dout1[63] sram0_dout1[6]
+ sram0_dout1[7] sram0_dout1[8] sram0_dout1[9] sram0_web0 sram0_wmask0[0] sram0_wmask0[1]
+ sram0_wmask0[2] sram0_wmask0[3] sram1_addr0[0] sram1_addr0[1] sram1_addr0[2] sram1_addr0[3]
+ sram1_addr0[4] sram1_addr0[5] sram1_addr0[6] sram1_addr0[7] sram1_addr0[8] sram1_addr1[0]
+ sram1_addr1[1] sram1_addr1[2] sram1_addr1[3] sram1_addr1[4] sram1_addr1[5] sram1_addr1[6]
+ sram1_addr1[7] sram1_addr1[8] sram1_clk0 sram1_clk1 sram1_csb0[0] sram1_csb0[1]
+ sram1_csb1[0] sram1_csb1[1] sram1_din0[0] sram1_din0[10] sram1_din0[11] sram1_din0[12]
+ sram1_din0[13] sram1_din0[14] sram1_din0[15] sram1_din0[16] sram1_din0[17] sram1_din0[18]
+ sram1_din0[19] sram1_din0[1] sram1_din0[20] sram1_din0[21] sram1_din0[22] sram1_din0[23]
+ sram1_din0[24] sram1_din0[25] sram1_din0[26] sram1_din0[27] sram1_din0[28] sram1_din0[29]
+ sram1_din0[2] sram1_din0[30] sram1_din0[31] sram1_din0[3] sram1_din0[4] sram1_din0[5]
+ sram1_din0[6] sram1_din0[7] sram1_din0[8] sram1_din0[9] sram1_dout0[0] sram1_dout0[10]
+ sram1_dout0[11] sram1_dout0[12] sram1_dout0[13] sram1_dout0[14] sram1_dout0[15]
+ sram1_dout0[16] sram1_dout0[17] sram1_dout0[18] sram1_dout0[19] sram1_dout0[1] sram1_dout0[20]
+ sram1_dout0[21] sram1_dout0[22] sram1_dout0[23] sram1_dout0[24] sram1_dout0[25]
+ sram1_dout0[26] sram1_dout0[27] sram1_dout0[28] sram1_dout0[29] sram1_dout0[2] sram1_dout0[30]
+ sram1_dout0[31] sram1_dout0[32] sram1_dout0[33] sram1_dout0[34] sram1_dout0[35]
+ sram1_dout0[36] sram1_dout0[37] sram1_dout0[38] sram1_dout0[39] sram1_dout0[3] sram1_dout0[40]
+ sram1_dout0[41] sram1_dout0[42] sram1_dout0[43] sram1_dout0[44] sram1_dout0[45]
+ sram1_dout0[46] sram1_dout0[47] sram1_dout0[48] sram1_dout0[49] sram1_dout0[4] sram1_dout0[50]
+ sram1_dout0[51] sram1_dout0[52] sram1_dout0[53] sram1_dout0[54] sram1_dout0[55]
+ sram1_dout0[56] sram1_dout0[57] sram1_dout0[58] sram1_dout0[59] sram1_dout0[5] sram1_dout0[60]
+ sram1_dout0[61] sram1_dout0[62] sram1_dout0[63] sram1_dout0[6] sram1_dout0[7] sram1_dout0[8]
+ sram1_dout0[9] sram1_dout1[0] sram1_dout1[10] sram1_dout1[11] sram1_dout1[12] sram1_dout1[13]
+ sram1_dout1[14] sram1_dout1[15] sram1_dout1[16] sram1_dout1[17] sram1_dout1[18]
+ sram1_dout1[19] sram1_dout1[1] sram1_dout1[20] sram1_dout1[21] sram1_dout1[22] sram1_dout1[23]
+ sram1_dout1[24] sram1_dout1[25] sram1_dout1[26] sram1_dout1[27] sram1_dout1[28]
+ sram1_dout1[29] sram1_dout1[2] sram1_dout1[30] sram1_dout1[31] sram1_dout1[32] sram1_dout1[33]
+ sram1_dout1[34] sram1_dout1[35] sram1_dout1[36] sram1_dout1[37] sram1_dout1[38]
+ sram1_dout1[39] sram1_dout1[3] sram1_dout1[40] sram1_dout1[41] sram1_dout1[42] sram1_dout1[43]
+ sram1_dout1[44] sram1_dout1[45] sram1_dout1[46] sram1_dout1[47] sram1_dout1[48]
+ sram1_dout1[49] sram1_dout1[4] sram1_dout1[50] sram1_dout1[51] sram1_dout1[52] sram1_dout1[53]
+ sram1_dout1[54] sram1_dout1[55] sram1_dout1[56] sram1_dout1[57] sram1_dout1[58]
+ sram1_dout1[59] sram1_dout1[5] sram1_dout1[60] sram1_dout1[61] sram1_dout1[62] sram1_dout1[63]
+ sram1_dout1[6] sram1_dout1[7] sram1_dout1[8] sram1_dout1[9] sram1_web0 sram1_wmask0[0]
+ sram1_wmask0[1] sram1_wmask0[2] sram1_wmask0[3] vccd1 vga_b[0] vga_b[1] vga_g[0]
+ vga_g[1] vga_hsync vga_r[0] vga_r[1] vga_vsync video_irq[0] video_irq[1] vssd1 wb_ack_o
+ wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15]
+ wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21]
+ wb_adr_i[22] wb_adr_i[23] wb_adr_i[2] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6]
+ wb_adr_i[7] wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_data_i[0] wb_data_i[10]
+ wb_data_i[11] wb_data_i[12] wb_data_i[13] wb_data_i[14] wb_data_i[15] wb_data_i[16]
+ wb_data_i[17] wb_data_i[18] wb_data_i[19] wb_data_i[1] wb_data_i[20] wb_data_i[21]
+ wb_data_i[22] wb_data_i[23] wb_data_i[24] wb_data_i[25] wb_data_i[26] wb_data_i[27]
+ wb_data_i[28] wb_data_i[29] wb_data_i[2] wb_data_i[30] wb_data_i[31] wb_data_i[3]
+ wb_data_i[4] wb_data_i[5] wb_data_i[6] wb_data_i[7] wb_data_i[8] wb_data_i[9] wb_data_o[0]
+ wb_data_o[10] wb_data_o[11] wb_data_o[12] wb_data_o[13] wb_data_o[14] wb_data_o[15]
+ wb_data_o[16] wb_data_o[17] wb_data_o[18] wb_data_o[19] wb_data_o[1] wb_data_o[20]
+ wb_data_o[21] wb_data_o[22] wb_data_o[23] wb_data_o[24] wb_data_o[25] wb_data_o[26]
+ wb_data_o[27] wb_data_o[28] wb_data_o[29] wb_data_o[2] wb_data_o[30] wb_data_o[31]
+ wb_data_o[3] wb_data_o[4] wb_data_o[5] wb_data_o[6] wb_data_o[7] wb_data_o[8] wb_data_o[9]
+ wb_error_o wb_rst_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stall_o wb_stb_i
+ wb_we_i
.ends

* Black-box entry subcircuit for Flash abstract view
.subckt Flash flash_csb flash_io0_read flash_io0_we flash_io0_write flash_io1_read
+ flash_io1_we flash_io1_write flash_sck sram_addr0[0] sram_addr0[1] sram_addr0[2]
+ sram_addr0[3] sram_addr0[4] sram_addr0[5] sram_addr0[6] sram_addr0[7] sram_addr0[8]
+ sram_addr1[0] sram_addr1[1] sram_addr1[2] sram_addr1[3] sram_addr1[4] sram_addr1[5]
+ sram_addr1[6] sram_addr1[7] sram_addr1[8] sram_clk0 sram_clk1 sram_csb0 sram_csb1
+ sram_din0[0] sram_din0[10] sram_din0[11] sram_din0[12] sram_din0[13] sram_din0[14]
+ sram_din0[15] sram_din0[16] sram_din0[17] sram_din0[18] sram_din0[19] sram_din0[1]
+ sram_din0[20] sram_din0[21] sram_din0[22] sram_din0[23] sram_din0[24] sram_din0[25]
+ sram_din0[26] sram_din0[27] sram_din0[28] sram_din0[29] sram_din0[2] sram_din0[30]
+ sram_din0[31] sram_din0[3] sram_din0[4] sram_din0[5] sram_din0[6] sram_din0[7] sram_din0[8]
+ sram_din0[9] sram_dout0[0] sram_dout0[10] sram_dout0[11] sram_dout0[12] sram_dout0[13]
+ sram_dout0[14] sram_dout0[15] sram_dout0[16] sram_dout0[17] sram_dout0[18] sram_dout0[19]
+ sram_dout0[1] sram_dout0[20] sram_dout0[21] sram_dout0[22] sram_dout0[23] sram_dout0[24]
+ sram_dout0[25] sram_dout0[26] sram_dout0[27] sram_dout0[28] sram_dout0[29] sram_dout0[2]
+ sram_dout0[30] sram_dout0[31] sram_dout0[3] sram_dout0[4] sram_dout0[5] sram_dout0[6]
+ sram_dout0[7] sram_dout0[8] sram_dout0[9] sram_dout1[0] sram_dout1[10] sram_dout1[11]
+ sram_dout1[12] sram_dout1[13] sram_dout1[14] sram_dout1[15] sram_dout1[16] sram_dout1[17]
+ sram_dout1[18] sram_dout1[19] sram_dout1[1] sram_dout1[20] sram_dout1[21] sram_dout1[22]
+ sram_dout1[23] sram_dout1[24] sram_dout1[25] sram_dout1[26] sram_dout1[27] sram_dout1[28]
+ sram_dout1[29] sram_dout1[2] sram_dout1[30] sram_dout1[31] sram_dout1[3] sram_dout1[4]
+ sram_dout1[5] sram_dout1[6] sram_dout1[7] sram_dout1[8] sram_dout1[9] sram_web0
+ sram_wmask0[0] sram_wmask0[1] sram_wmask0[2] sram_wmask0[3] vccd1 vssd1 wb_ack_o
+ wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15]
+ wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21]
+ wb_adr_i[22] wb_adr_i[23] wb_adr_i[2] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6]
+ wb_adr_i[7] wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_data_i[0] wb_data_i[10]
+ wb_data_i[11] wb_data_i[12] wb_data_i[13] wb_data_i[14] wb_data_i[15] wb_data_i[16]
+ wb_data_i[17] wb_data_i[18] wb_data_i[19] wb_data_i[1] wb_data_i[20] wb_data_i[21]
+ wb_data_i[22] wb_data_i[23] wb_data_i[24] wb_data_i[25] wb_data_i[26] wb_data_i[27]
+ wb_data_i[28] wb_data_i[29] wb_data_i[2] wb_data_i[30] wb_data_i[31] wb_data_i[3]
+ wb_data_i[4] wb_data_i[5] wb_data_i[6] wb_data_i[7] wb_data_i[8] wb_data_i[9] wb_data_o[0]
+ wb_data_o[10] wb_data_o[11] wb_data_o[12] wb_data_o[13] wb_data_o[14] wb_data_o[15]
+ wb_data_o[16] wb_data_o[17] wb_data_o[18] wb_data_o[19] wb_data_o[1] wb_data_o[20]
+ wb_data_o[21] wb_data_o[22] wb_data_o[23] wb_data_o[24] wb_data_o[25] wb_data_o[26]
+ wb_data_o[27] wb_data_o[28] wb_data_o[29] wb_data_o[2] wb_data_o[30] wb_data_o[31]
+ wb_data_o[3] wb_data_o[4] wb_data_o[5] wb_data_o[6] wb_data_o[7] wb_data_o[8] wb_data_o[9]
+ wb_error_o wb_rst_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stall_o wb_stb_i
+ wb_we_i
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XexperiarSoC_videoSRAM0 experiarSoC_videoSRAM1/din0[0] experiarSoC_videoSRAM1/din0[1]
+ experiarSoC_videoSRAM1/din0[2] experiarSoC_videoSRAM1/din0[3] experiarSoC_videoSRAM1/din0[4]
+ experiarSoC_videoSRAM1/din0[5] experiarSoC_videoSRAM1/din0[6] experiarSoC_videoSRAM1/din0[7]
+ experiarSoC_videoSRAM1/din0[8] experiarSoC_videoSRAM1/din0[9] experiarSoC_videoSRAM1/din0[10]
+ experiarSoC_videoSRAM1/din0[11] experiarSoC_videoSRAM1/din0[12] experiarSoC_videoSRAM1/din0[13]
+ experiarSoC_videoSRAM1/din0[14] experiarSoC_videoSRAM1/din0[15] experiarSoC_videoSRAM1/din0[16]
+ experiarSoC_videoSRAM1/din0[17] experiarSoC_videoSRAM1/din0[18] experiarSoC_videoSRAM1/din0[19]
+ experiarSoC_videoSRAM1/din0[20] experiarSoC_videoSRAM1/din0[21] experiarSoC_videoSRAM1/din0[22]
+ experiarSoC_videoSRAM1/din0[23] experiarSoC_videoSRAM1/din0[24] experiarSoC_videoSRAM1/din0[25]
+ experiarSoC_videoSRAM1/din0[26] experiarSoC_videoSRAM1/din0[27] experiarSoC_videoSRAM1/din0[28]
+ experiarSoC_videoSRAM1/din0[29] experiarSoC_videoSRAM1/din0[30] experiarSoC_videoSRAM1/din0[31]
+ experiarSoC_videoSRAM1/addr0[0] experiarSoC_videoSRAM1/addr0[1] experiarSoC_videoSRAM1/addr0[2]
+ experiarSoC_videoSRAM1/addr0[3] experiarSoC_videoSRAM1/addr0[4] experiarSoC_videoSRAM1/addr0[5]
+ experiarSoC_videoSRAM1/addr0[6] experiarSoC_videoSRAM1/addr0[7] experiarSoC_videoSRAM1/addr0[8]
+ experiarSoC_videoSRAM1/addr1[0] experiarSoC_videoSRAM1/addr1[1] experiarSoC_videoSRAM1/addr1[2]
+ experiarSoC_videoSRAM1/addr1[3] experiarSoC_videoSRAM1/addr1[4] experiarSoC_videoSRAM1/addr1[5]
+ experiarSoC_videoSRAM1/addr1[6] experiarSoC_videoSRAM1/addr1[7] experiarSoC_videoSRAM1/addr1[8]
+ experiarSoC_videoSRAM0/csb0 experiarSoC_videoSRAM0/csb1 experiarSoC_videoSRAM1/web0
+ experiarSoC_videoSRAM1/clk0 experiarSoC_videoSRAM1/clk1 experiarSoC_videoSRAM1/wmask0[0]
+ experiarSoC_videoSRAM1/wmask0[1] experiarSoC_videoSRAM1/wmask0[2] experiarSoC_videoSRAM1/wmask0[3]
+ experiarSoC_videoSRAM0/dout0[0] experiarSoC_videoSRAM0/dout0[1] experiarSoC_videoSRAM0/dout0[2]
+ experiarSoC_videoSRAM0/dout0[3] experiarSoC_videoSRAM0/dout0[4] experiarSoC_videoSRAM0/dout0[5]
+ experiarSoC_videoSRAM0/dout0[6] experiarSoC_videoSRAM0/dout0[7] experiarSoC_videoSRAM0/dout0[8]
+ experiarSoC_videoSRAM0/dout0[9] experiarSoC_videoSRAM0/dout0[10] experiarSoC_videoSRAM0/dout0[11]
+ experiarSoC_videoSRAM0/dout0[12] experiarSoC_videoSRAM0/dout0[13] experiarSoC_videoSRAM0/dout0[14]
+ experiarSoC_videoSRAM0/dout0[15] experiarSoC_videoSRAM0/dout0[16] experiarSoC_videoSRAM0/dout0[17]
+ experiarSoC_videoSRAM0/dout0[18] experiarSoC_videoSRAM0/dout0[19] experiarSoC_videoSRAM0/dout0[20]
+ experiarSoC_videoSRAM0/dout0[21] experiarSoC_videoSRAM0/dout0[22] experiarSoC_videoSRAM0/dout0[23]
+ experiarSoC_videoSRAM0/dout0[24] experiarSoC_videoSRAM0/dout0[25] experiarSoC_videoSRAM0/dout0[26]
+ experiarSoC_videoSRAM0/dout0[27] experiarSoC_videoSRAM0/dout0[28] experiarSoC_videoSRAM0/dout0[29]
+ experiarSoC_videoSRAM0/dout0[30] experiarSoC_videoSRAM0/dout0[31] experiarSoC_videoSRAM0/dout1[0]
+ experiarSoC_videoSRAM0/dout1[1] experiarSoC_videoSRAM0/dout1[2] experiarSoC_videoSRAM0/dout1[3]
+ experiarSoC_videoSRAM0/dout1[4] experiarSoC_videoSRAM0/dout1[5] experiarSoC_videoSRAM0/dout1[6]
+ experiarSoC_videoSRAM0/dout1[7] experiarSoC_videoSRAM0/dout1[8] experiarSoC_videoSRAM0/dout1[9]
+ experiarSoC_videoSRAM0/dout1[10] experiarSoC_videoSRAM0/dout1[11] experiarSoC_videoSRAM0/dout1[12]
+ experiarSoC_videoSRAM0/dout1[13] experiarSoC_videoSRAM0/dout1[14] experiarSoC_videoSRAM0/dout1[15]
+ experiarSoC_videoSRAM0/dout1[16] experiarSoC_videoSRAM0/dout1[17] experiarSoC_videoSRAM0/dout1[18]
+ experiarSoC_videoSRAM0/dout1[19] experiarSoC_videoSRAM0/dout1[20] experiarSoC_videoSRAM0/dout1[21]
+ experiarSoC_videoSRAM0/dout1[22] experiarSoC_videoSRAM0/dout1[23] experiarSoC_videoSRAM0/dout1[24]
+ experiarSoC_videoSRAM0/dout1[25] experiarSoC_videoSRAM0/dout1[26] experiarSoC_videoSRAM0/dout1[27]
+ experiarSoC_videoSRAM0/dout1[28] experiarSoC_videoSRAM0/dout1[29] experiarSoC_videoSRAM0/dout1[30]
+ experiarSoC_videoSRAM0/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_videoSRAM1 experiarSoC_videoSRAM1/din0[0] experiarSoC_videoSRAM1/din0[1]
+ experiarSoC_videoSRAM1/din0[2] experiarSoC_videoSRAM1/din0[3] experiarSoC_videoSRAM1/din0[4]
+ experiarSoC_videoSRAM1/din0[5] experiarSoC_videoSRAM1/din0[6] experiarSoC_videoSRAM1/din0[7]
+ experiarSoC_videoSRAM1/din0[8] experiarSoC_videoSRAM1/din0[9] experiarSoC_videoSRAM1/din0[10]
+ experiarSoC_videoSRAM1/din0[11] experiarSoC_videoSRAM1/din0[12] experiarSoC_videoSRAM1/din0[13]
+ experiarSoC_videoSRAM1/din0[14] experiarSoC_videoSRAM1/din0[15] experiarSoC_videoSRAM1/din0[16]
+ experiarSoC_videoSRAM1/din0[17] experiarSoC_videoSRAM1/din0[18] experiarSoC_videoSRAM1/din0[19]
+ experiarSoC_videoSRAM1/din0[20] experiarSoC_videoSRAM1/din0[21] experiarSoC_videoSRAM1/din0[22]
+ experiarSoC_videoSRAM1/din0[23] experiarSoC_videoSRAM1/din0[24] experiarSoC_videoSRAM1/din0[25]
+ experiarSoC_videoSRAM1/din0[26] experiarSoC_videoSRAM1/din0[27] experiarSoC_videoSRAM1/din0[28]
+ experiarSoC_videoSRAM1/din0[29] experiarSoC_videoSRAM1/din0[30] experiarSoC_videoSRAM1/din0[31]
+ experiarSoC_videoSRAM1/addr0[0] experiarSoC_videoSRAM1/addr0[1] experiarSoC_videoSRAM1/addr0[2]
+ experiarSoC_videoSRAM1/addr0[3] experiarSoC_videoSRAM1/addr0[4] experiarSoC_videoSRAM1/addr0[5]
+ experiarSoC_videoSRAM1/addr0[6] experiarSoC_videoSRAM1/addr0[7] experiarSoC_videoSRAM1/addr0[8]
+ experiarSoC_videoSRAM1/addr1[0] experiarSoC_videoSRAM1/addr1[1] experiarSoC_videoSRAM1/addr1[2]
+ experiarSoC_videoSRAM1/addr1[3] experiarSoC_videoSRAM1/addr1[4] experiarSoC_videoSRAM1/addr1[5]
+ experiarSoC_videoSRAM1/addr1[6] experiarSoC_videoSRAM1/addr1[7] experiarSoC_videoSRAM1/addr1[8]
+ experiarSoC_videoSRAM1/csb0 experiarSoC_videoSRAM1/csb1 experiarSoC_videoSRAM1/web0
+ experiarSoC_videoSRAM1/clk0 experiarSoC_videoSRAM1/clk1 experiarSoC_videoSRAM1/wmask0[0]
+ experiarSoC_videoSRAM1/wmask0[1] experiarSoC_videoSRAM1/wmask0[2] experiarSoC_videoSRAM1/wmask0[3]
+ experiarSoC_videoSRAM1/dout0[0] experiarSoC_videoSRAM1/dout0[1] experiarSoC_videoSRAM1/dout0[2]
+ experiarSoC_videoSRAM1/dout0[3] experiarSoC_videoSRAM1/dout0[4] experiarSoC_videoSRAM1/dout0[5]
+ experiarSoC_videoSRAM1/dout0[6] experiarSoC_videoSRAM1/dout0[7] experiarSoC_videoSRAM1/dout0[8]
+ experiarSoC_videoSRAM1/dout0[9] experiarSoC_videoSRAM1/dout0[10] experiarSoC_videoSRAM1/dout0[11]
+ experiarSoC_videoSRAM1/dout0[12] experiarSoC_videoSRAM1/dout0[13] experiarSoC_videoSRAM1/dout0[14]
+ experiarSoC_videoSRAM1/dout0[15] experiarSoC_videoSRAM1/dout0[16] experiarSoC_videoSRAM1/dout0[17]
+ experiarSoC_videoSRAM1/dout0[18] experiarSoC_videoSRAM1/dout0[19] experiarSoC_videoSRAM1/dout0[20]
+ experiarSoC_videoSRAM1/dout0[21] experiarSoC_videoSRAM1/dout0[22] experiarSoC_videoSRAM1/dout0[23]
+ experiarSoC_videoSRAM1/dout0[24] experiarSoC_videoSRAM1/dout0[25] experiarSoC_videoSRAM1/dout0[26]
+ experiarSoC_videoSRAM1/dout0[27] experiarSoC_videoSRAM1/dout0[28] experiarSoC_videoSRAM1/dout0[29]
+ experiarSoC_videoSRAM1/dout0[30] experiarSoC_videoSRAM1/dout0[31] experiarSoC_videoSRAM1/dout1[0]
+ experiarSoC_videoSRAM1/dout1[1] experiarSoC_videoSRAM1/dout1[2] experiarSoC_videoSRAM1/dout1[3]
+ experiarSoC_videoSRAM1/dout1[4] experiarSoC_videoSRAM1/dout1[5] experiarSoC_videoSRAM1/dout1[6]
+ experiarSoC_videoSRAM1/dout1[7] experiarSoC_videoSRAM1/dout1[8] experiarSoC_videoSRAM1/dout1[9]
+ experiarSoC_videoSRAM1/dout1[10] experiarSoC_videoSRAM1/dout1[11] experiarSoC_videoSRAM1/dout1[12]
+ experiarSoC_videoSRAM1/dout1[13] experiarSoC_videoSRAM1/dout1[14] experiarSoC_videoSRAM1/dout1[15]
+ experiarSoC_videoSRAM1/dout1[16] experiarSoC_videoSRAM1/dout1[17] experiarSoC_videoSRAM1/dout1[18]
+ experiarSoC_videoSRAM1/dout1[19] experiarSoC_videoSRAM1/dout1[20] experiarSoC_videoSRAM1/dout1[21]
+ experiarSoC_videoSRAM1/dout1[22] experiarSoC_videoSRAM1/dout1[23] experiarSoC_videoSRAM1/dout1[24]
+ experiarSoC_videoSRAM1/dout1[25] experiarSoC_videoSRAM1/dout1[26] experiarSoC_videoSRAM1/dout1[27]
+ experiarSoC_videoSRAM1/dout1[28] experiarSoC_videoSRAM1/dout1[29] experiarSoC_videoSRAM1/dout1[30]
+ experiarSoC_videoSRAM1/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_videoSRAM2 experiarSoC_videoSRAM3/din0[0] experiarSoC_videoSRAM3/din0[1]
+ experiarSoC_videoSRAM3/din0[2] experiarSoC_videoSRAM3/din0[3] experiarSoC_videoSRAM3/din0[4]
+ experiarSoC_videoSRAM3/din0[5] experiarSoC_videoSRAM3/din0[6] experiarSoC_videoSRAM3/din0[7]
+ experiarSoC_videoSRAM3/din0[8] experiarSoC_videoSRAM3/din0[9] experiarSoC_videoSRAM3/din0[10]
+ experiarSoC_videoSRAM3/din0[11] experiarSoC_videoSRAM3/din0[12] experiarSoC_videoSRAM3/din0[13]
+ experiarSoC_videoSRAM3/din0[14] experiarSoC_videoSRAM3/din0[15] experiarSoC_videoSRAM3/din0[16]
+ experiarSoC_videoSRAM3/din0[17] experiarSoC_videoSRAM3/din0[18] experiarSoC_videoSRAM3/din0[19]
+ experiarSoC_videoSRAM3/din0[20] experiarSoC_videoSRAM3/din0[21] experiarSoC_videoSRAM3/din0[22]
+ experiarSoC_videoSRAM3/din0[23] experiarSoC_videoSRAM3/din0[24] experiarSoC_videoSRAM3/din0[25]
+ experiarSoC_videoSRAM3/din0[26] experiarSoC_videoSRAM3/din0[27] experiarSoC_videoSRAM3/din0[28]
+ experiarSoC_videoSRAM3/din0[29] experiarSoC_videoSRAM3/din0[30] experiarSoC_videoSRAM3/din0[31]
+ experiarSoC_videoSRAM3/addr0[0] experiarSoC_videoSRAM3/addr0[1] experiarSoC_videoSRAM3/addr0[2]
+ experiarSoC_videoSRAM3/addr0[3] experiarSoC_videoSRAM3/addr0[4] experiarSoC_videoSRAM3/addr0[5]
+ experiarSoC_videoSRAM3/addr0[6] experiarSoC_videoSRAM3/addr0[7] experiarSoC_videoSRAM3/addr0[8]
+ experiarSoC_videoSRAM3/addr1[0] experiarSoC_videoSRAM3/addr1[1] experiarSoC_videoSRAM3/addr1[2]
+ experiarSoC_videoSRAM3/addr1[3] experiarSoC_videoSRAM3/addr1[4] experiarSoC_videoSRAM3/addr1[5]
+ experiarSoC_videoSRAM3/addr1[6] experiarSoC_videoSRAM3/addr1[7] experiarSoC_videoSRAM3/addr1[8]
+ experiarSoC_videoSRAM2/csb0 experiarSoC_videoSRAM2/csb1 experiarSoC_videoSRAM3/web0
+ experiarSoC_videoSRAM3/clk0 experiarSoC_videoSRAM3/clk1 experiarSoC_videoSRAM3/wmask0[0]
+ experiarSoC_videoSRAM3/wmask0[1] experiarSoC_videoSRAM3/wmask0[2] experiarSoC_videoSRAM3/wmask0[3]
+ experiarSoC_videoSRAM2/dout0[0] experiarSoC_videoSRAM2/dout0[1] experiarSoC_videoSRAM2/dout0[2]
+ experiarSoC_videoSRAM2/dout0[3] experiarSoC_videoSRAM2/dout0[4] experiarSoC_videoSRAM2/dout0[5]
+ experiarSoC_videoSRAM2/dout0[6] experiarSoC_videoSRAM2/dout0[7] experiarSoC_videoSRAM2/dout0[8]
+ experiarSoC_videoSRAM2/dout0[9] experiarSoC_videoSRAM2/dout0[10] experiarSoC_videoSRAM2/dout0[11]
+ experiarSoC_videoSRAM2/dout0[12] experiarSoC_videoSRAM2/dout0[13] experiarSoC_videoSRAM2/dout0[14]
+ experiarSoC_videoSRAM2/dout0[15] experiarSoC_videoSRAM2/dout0[16] experiarSoC_videoSRAM2/dout0[17]
+ experiarSoC_videoSRAM2/dout0[18] experiarSoC_videoSRAM2/dout0[19] experiarSoC_videoSRAM2/dout0[20]
+ experiarSoC_videoSRAM2/dout0[21] experiarSoC_videoSRAM2/dout0[22] experiarSoC_videoSRAM2/dout0[23]
+ experiarSoC_videoSRAM2/dout0[24] experiarSoC_videoSRAM2/dout0[25] experiarSoC_videoSRAM2/dout0[26]
+ experiarSoC_videoSRAM2/dout0[27] experiarSoC_videoSRAM2/dout0[28] experiarSoC_videoSRAM2/dout0[29]
+ experiarSoC_videoSRAM2/dout0[30] experiarSoC_videoSRAM2/dout0[31] experiarSoC_videoSRAM2/dout1[0]
+ experiarSoC_videoSRAM2/dout1[1] experiarSoC_videoSRAM2/dout1[2] experiarSoC_videoSRAM2/dout1[3]
+ experiarSoC_videoSRAM2/dout1[4] experiarSoC_videoSRAM2/dout1[5] experiarSoC_videoSRAM2/dout1[6]
+ experiarSoC_videoSRAM2/dout1[7] experiarSoC_videoSRAM2/dout1[8] experiarSoC_videoSRAM2/dout1[9]
+ experiarSoC_videoSRAM2/dout1[10] experiarSoC_videoSRAM2/dout1[11] experiarSoC_videoSRAM2/dout1[12]
+ experiarSoC_videoSRAM2/dout1[13] experiarSoC_videoSRAM2/dout1[14] experiarSoC_videoSRAM2/dout1[15]
+ experiarSoC_videoSRAM2/dout1[16] experiarSoC_videoSRAM2/dout1[17] experiarSoC_videoSRAM2/dout1[18]
+ experiarSoC_videoSRAM2/dout1[19] experiarSoC_videoSRAM2/dout1[20] experiarSoC_videoSRAM2/dout1[21]
+ experiarSoC_videoSRAM2/dout1[22] experiarSoC_videoSRAM2/dout1[23] experiarSoC_videoSRAM2/dout1[24]
+ experiarSoC_videoSRAM2/dout1[25] experiarSoC_videoSRAM2/dout1[26] experiarSoC_videoSRAM2/dout1[27]
+ experiarSoC_videoSRAM2/dout1[28] experiarSoC_videoSRAM2/dout1[29] experiarSoC_videoSRAM2/dout1[30]
+ experiarSoC_videoSRAM2/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_videoSRAM3 experiarSoC_videoSRAM3/din0[0] experiarSoC_videoSRAM3/din0[1]
+ experiarSoC_videoSRAM3/din0[2] experiarSoC_videoSRAM3/din0[3] experiarSoC_videoSRAM3/din0[4]
+ experiarSoC_videoSRAM3/din0[5] experiarSoC_videoSRAM3/din0[6] experiarSoC_videoSRAM3/din0[7]
+ experiarSoC_videoSRAM3/din0[8] experiarSoC_videoSRAM3/din0[9] experiarSoC_videoSRAM3/din0[10]
+ experiarSoC_videoSRAM3/din0[11] experiarSoC_videoSRAM3/din0[12] experiarSoC_videoSRAM3/din0[13]
+ experiarSoC_videoSRAM3/din0[14] experiarSoC_videoSRAM3/din0[15] experiarSoC_videoSRAM3/din0[16]
+ experiarSoC_videoSRAM3/din0[17] experiarSoC_videoSRAM3/din0[18] experiarSoC_videoSRAM3/din0[19]
+ experiarSoC_videoSRAM3/din0[20] experiarSoC_videoSRAM3/din0[21] experiarSoC_videoSRAM3/din0[22]
+ experiarSoC_videoSRAM3/din0[23] experiarSoC_videoSRAM3/din0[24] experiarSoC_videoSRAM3/din0[25]
+ experiarSoC_videoSRAM3/din0[26] experiarSoC_videoSRAM3/din0[27] experiarSoC_videoSRAM3/din0[28]
+ experiarSoC_videoSRAM3/din0[29] experiarSoC_videoSRAM3/din0[30] experiarSoC_videoSRAM3/din0[31]
+ experiarSoC_videoSRAM3/addr0[0] experiarSoC_videoSRAM3/addr0[1] experiarSoC_videoSRAM3/addr0[2]
+ experiarSoC_videoSRAM3/addr0[3] experiarSoC_videoSRAM3/addr0[4] experiarSoC_videoSRAM3/addr0[5]
+ experiarSoC_videoSRAM3/addr0[6] experiarSoC_videoSRAM3/addr0[7] experiarSoC_videoSRAM3/addr0[8]
+ experiarSoC_videoSRAM3/addr1[0] experiarSoC_videoSRAM3/addr1[1] experiarSoC_videoSRAM3/addr1[2]
+ experiarSoC_videoSRAM3/addr1[3] experiarSoC_videoSRAM3/addr1[4] experiarSoC_videoSRAM3/addr1[5]
+ experiarSoC_videoSRAM3/addr1[6] experiarSoC_videoSRAM3/addr1[7] experiarSoC_videoSRAM3/addr1[8]
+ experiarSoC_videoSRAM3/csb0 experiarSoC_videoSRAM3/csb1 experiarSoC_videoSRAM3/web0
+ experiarSoC_videoSRAM3/clk0 experiarSoC_videoSRAM3/clk1 experiarSoC_videoSRAM3/wmask0[0]
+ experiarSoC_videoSRAM3/wmask0[1] experiarSoC_videoSRAM3/wmask0[2] experiarSoC_videoSRAM3/wmask0[3]
+ experiarSoC_videoSRAM3/dout0[0] experiarSoC_videoSRAM3/dout0[1] experiarSoC_videoSRAM3/dout0[2]
+ experiarSoC_videoSRAM3/dout0[3] experiarSoC_videoSRAM3/dout0[4] experiarSoC_videoSRAM3/dout0[5]
+ experiarSoC_videoSRAM3/dout0[6] experiarSoC_videoSRAM3/dout0[7] experiarSoC_videoSRAM3/dout0[8]
+ experiarSoC_videoSRAM3/dout0[9] experiarSoC_videoSRAM3/dout0[10] experiarSoC_videoSRAM3/dout0[11]
+ experiarSoC_videoSRAM3/dout0[12] experiarSoC_videoSRAM3/dout0[13] experiarSoC_videoSRAM3/dout0[14]
+ experiarSoC_videoSRAM3/dout0[15] experiarSoC_videoSRAM3/dout0[16] experiarSoC_videoSRAM3/dout0[17]
+ experiarSoC_videoSRAM3/dout0[18] experiarSoC_videoSRAM3/dout0[19] experiarSoC_videoSRAM3/dout0[20]
+ experiarSoC_videoSRAM3/dout0[21] experiarSoC_videoSRAM3/dout0[22] experiarSoC_videoSRAM3/dout0[23]
+ experiarSoC_videoSRAM3/dout0[24] experiarSoC_videoSRAM3/dout0[25] experiarSoC_videoSRAM3/dout0[26]
+ experiarSoC_videoSRAM3/dout0[27] experiarSoC_videoSRAM3/dout0[28] experiarSoC_videoSRAM3/dout0[29]
+ experiarSoC_videoSRAM3/dout0[30] experiarSoC_videoSRAM3/dout0[31] experiarSoC_videoSRAM3/dout1[0]
+ experiarSoC_videoSRAM3/dout1[1] experiarSoC_videoSRAM3/dout1[2] experiarSoC_videoSRAM3/dout1[3]
+ experiarSoC_videoSRAM3/dout1[4] experiarSoC_videoSRAM3/dout1[5] experiarSoC_videoSRAM3/dout1[6]
+ experiarSoC_videoSRAM3/dout1[7] experiarSoC_videoSRAM3/dout1[8] experiarSoC_videoSRAM3/dout1[9]
+ experiarSoC_videoSRAM3/dout1[10] experiarSoC_videoSRAM3/dout1[11] experiarSoC_videoSRAM3/dout1[12]
+ experiarSoC_videoSRAM3/dout1[13] experiarSoC_videoSRAM3/dout1[14] experiarSoC_videoSRAM3/dout1[15]
+ experiarSoC_videoSRAM3/dout1[16] experiarSoC_videoSRAM3/dout1[17] experiarSoC_videoSRAM3/dout1[18]
+ experiarSoC_videoSRAM3/dout1[19] experiarSoC_videoSRAM3/dout1[20] experiarSoC_videoSRAM3/dout1[21]
+ experiarSoC_videoSRAM3/dout1[22] experiarSoC_videoSRAM3/dout1[23] experiarSoC_videoSRAM3/dout1[24]
+ experiarSoC_videoSRAM3/dout1[25] experiarSoC_videoSRAM3/dout1[26] experiarSoC_videoSRAM3/dout1[27]
+ experiarSoC_videoSRAM3/dout1[28] experiarSoC_videoSRAM3/dout1[29] experiarSoC_videoSRAM3/dout1[30]
+ experiarSoC_videoSRAM3/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_core0SRAM0 experiarSoC_core0/din0[0] experiarSoC_core0/din0[1] experiarSoC_core0/din0[2]
+ experiarSoC_core0/din0[3] experiarSoC_core0/din0[4] experiarSoC_core0/din0[5] experiarSoC_core0/din0[6]
+ experiarSoC_core0/din0[7] experiarSoC_core0/din0[8] experiarSoC_core0/din0[9] experiarSoC_core0/din0[10]
+ experiarSoC_core0/din0[11] experiarSoC_core0/din0[12] experiarSoC_core0/din0[13]
+ experiarSoC_core0/din0[14] experiarSoC_core0/din0[15] experiarSoC_core0/din0[16]
+ experiarSoC_core0/din0[17] experiarSoC_core0/din0[18] experiarSoC_core0/din0[19]
+ experiarSoC_core0/din0[20] experiarSoC_core0/din0[21] experiarSoC_core0/din0[22]
+ experiarSoC_core0/din0[23] experiarSoC_core0/din0[24] experiarSoC_core0/din0[25]
+ experiarSoC_core0/din0[26] experiarSoC_core0/din0[27] experiarSoC_core0/din0[28]
+ experiarSoC_core0/din0[29] experiarSoC_core0/din0[30] experiarSoC_core0/din0[31]
+ experiarSoC_core0/addr0[0] experiarSoC_core0/addr0[1] experiarSoC_core0/addr0[2]
+ experiarSoC_core0/addr0[3] experiarSoC_core0/addr0[4] experiarSoC_core0/addr0[5]
+ experiarSoC_core0/addr0[6] experiarSoC_core0/addr0[7] experiarSoC_core0/addr0[8]
+ experiarSoC_core0/addr1[0] experiarSoC_core0/addr1[1] experiarSoC_core0/addr1[2]
+ experiarSoC_core0/addr1[3] experiarSoC_core0/addr1[4] experiarSoC_core0/addr1[5]
+ experiarSoC_core0/addr1[6] experiarSoC_core0/addr1[7] experiarSoC_core0/addr1[8]
+ experiarSoC_core0/csb0[0] experiarSoC_core0/csb1[0] experiarSoC_core0/web0 experiarSoC_core0/clk0
+ experiarSoC_core0/clk1 experiarSoC_core0/wmask0[0] experiarSoC_core0/wmask0[1] experiarSoC_core0/wmask0[2]
+ experiarSoC_core0/wmask0[3] experiarSoC_core0/dout0[0] experiarSoC_core0/dout0[1]
+ experiarSoC_core0/dout0[2] experiarSoC_core0/dout0[3] experiarSoC_core0/dout0[4]
+ experiarSoC_core0/dout0[5] experiarSoC_core0/dout0[6] experiarSoC_core0/dout0[7]
+ experiarSoC_core0/dout0[8] experiarSoC_core0/dout0[9] experiarSoC_core0/dout0[10]
+ experiarSoC_core0/dout0[11] experiarSoC_core0/dout0[12] experiarSoC_core0/dout0[13]
+ experiarSoC_core0/dout0[14] experiarSoC_core0/dout0[15] experiarSoC_core0/dout0[16]
+ experiarSoC_core0/dout0[17] experiarSoC_core0/dout0[18] experiarSoC_core0/dout0[19]
+ experiarSoC_core0/dout0[20] experiarSoC_core0/dout0[21] experiarSoC_core0/dout0[22]
+ experiarSoC_core0/dout0[23] experiarSoC_core0/dout0[24] experiarSoC_core0/dout0[25]
+ experiarSoC_core0/dout0[26] experiarSoC_core0/dout0[27] experiarSoC_core0/dout0[28]
+ experiarSoC_core0/dout0[29] experiarSoC_core0/dout0[30] experiarSoC_core0/dout0[31]
+ experiarSoC_core0/dout1[0] experiarSoC_core0/dout1[1] experiarSoC_core0/dout1[2]
+ experiarSoC_core0/dout1[3] experiarSoC_core0/dout1[4] experiarSoC_core0/dout1[5]
+ experiarSoC_core0/dout1[6] experiarSoC_core0/dout1[7] experiarSoC_core0/dout1[8]
+ experiarSoC_core0/dout1[9] experiarSoC_core0/dout1[10] experiarSoC_core0/dout1[11]
+ experiarSoC_core0/dout1[12] experiarSoC_core0/dout1[13] experiarSoC_core0/dout1[14]
+ experiarSoC_core0/dout1[15] experiarSoC_core0/dout1[16] experiarSoC_core0/dout1[17]
+ experiarSoC_core0/dout1[18] experiarSoC_core0/dout1[19] experiarSoC_core0/dout1[20]
+ experiarSoC_core0/dout1[21] experiarSoC_core0/dout1[22] experiarSoC_core0/dout1[23]
+ experiarSoC_core0/dout1[24] experiarSoC_core0/dout1[25] experiarSoC_core0/dout1[26]
+ experiarSoC_core0/dout1[27] experiarSoC_core0/dout1[28] experiarSoC_core0/dout1[29]
+ experiarSoC_core0/dout1[30] experiarSoC_core0/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_core0SRAM1 experiarSoC_core0/din0[0] experiarSoC_core0/din0[1] experiarSoC_core0/din0[2]
+ experiarSoC_core0/din0[3] experiarSoC_core0/din0[4] experiarSoC_core0/din0[5] experiarSoC_core0/din0[6]
+ experiarSoC_core0/din0[7] experiarSoC_core0/din0[8] experiarSoC_core0/din0[9] experiarSoC_core0/din0[10]
+ experiarSoC_core0/din0[11] experiarSoC_core0/din0[12] experiarSoC_core0/din0[13]
+ experiarSoC_core0/din0[14] experiarSoC_core0/din0[15] experiarSoC_core0/din0[16]
+ experiarSoC_core0/din0[17] experiarSoC_core0/din0[18] experiarSoC_core0/din0[19]
+ experiarSoC_core0/din0[20] experiarSoC_core0/din0[21] experiarSoC_core0/din0[22]
+ experiarSoC_core0/din0[23] experiarSoC_core0/din0[24] experiarSoC_core0/din0[25]
+ experiarSoC_core0/din0[26] experiarSoC_core0/din0[27] experiarSoC_core0/din0[28]
+ experiarSoC_core0/din0[29] experiarSoC_core0/din0[30] experiarSoC_core0/din0[31]
+ experiarSoC_core0/addr0[0] experiarSoC_core0/addr0[1] experiarSoC_core0/addr0[2]
+ experiarSoC_core0/addr0[3] experiarSoC_core0/addr0[4] experiarSoC_core0/addr0[5]
+ experiarSoC_core0/addr0[6] experiarSoC_core0/addr0[7] experiarSoC_core0/addr0[8]
+ experiarSoC_core0/addr1[0] experiarSoC_core0/addr1[1] experiarSoC_core0/addr1[2]
+ experiarSoC_core0/addr1[3] experiarSoC_core0/addr1[4] experiarSoC_core0/addr1[5]
+ experiarSoC_core0/addr1[6] experiarSoC_core0/addr1[7] experiarSoC_core0/addr1[8]
+ experiarSoC_core0/csb0[1] experiarSoC_core0/csb1[1] experiarSoC_core0/web0 experiarSoC_core0/clk0
+ experiarSoC_core0/clk1 experiarSoC_core0/wmask0[0] experiarSoC_core0/wmask0[1] experiarSoC_core0/wmask0[2]
+ experiarSoC_core0/wmask0[3] experiarSoC_core0/dout0[32] experiarSoC_core0/dout0[33]
+ experiarSoC_core0/dout0[34] experiarSoC_core0/dout0[35] experiarSoC_core0/dout0[36]
+ experiarSoC_core0/dout0[37] experiarSoC_core0/dout0[38] experiarSoC_core0/dout0[39]
+ experiarSoC_core0/dout0[40] experiarSoC_core0/dout0[41] experiarSoC_core0/dout0[42]
+ experiarSoC_core0/dout0[43] experiarSoC_core0/dout0[44] experiarSoC_core0/dout0[45]
+ experiarSoC_core0/dout0[46] experiarSoC_core0/dout0[47] experiarSoC_core0/dout0[48]
+ experiarSoC_core0/dout0[49] experiarSoC_core0/dout0[50] experiarSoC_core0/dout0[51]
+ experiarSoC_core0/dout0[52] experiarSoC_core0/dout0[53] experiarSoC_core0/dout0[54]
+ experiarSoC_core0/dout0[55] experiarSoC_core0/dout0[56] experiarSoC_core0/dout0[57]
+ experiarSoC_core0/dout0[58] experiarSoC_core0/dout0[59] experiarSoC_core0/dout0[60]
+ experiarSoC_core0/dout0[61] experiarSoC_core0/dout0[62] experiarSoC_core0/dout0[63]
+ experiarSoC_core0/dout1[32] experiarSoC_core0/dout1[33] experiarSoC_core0/dout1[34]
+ experiarSoC_core0/dout1[35] experiarSoC_core0/dout1[36] experiarSoC_core0/dout1[37]
+ experiarSoC_core0/dout1[38] experiarSoC_core0/dout1[39] experiarSoC_core0/dout1[40]
+ experiarSoC_core0/dout1[41] experiarSoC_core0/dout1[42] experiarSoC_core0/dout1[43]
+ experiarSoC_core0/dout1[44] experiarSoC_core0/dout1[45] experiarSoC_core0/dout1[46]
+ experiarSoC_core0/dout1[47] experiarSoC_core0/dout1[48] experiarSoC_core0/dout1[49]
+ experiarSoC_core0/dout1[50] experiarSoC_core0/dout1[51] experiarSoC_core0/dout1[52]
+ experiarSoC_core0/dout1[53] experiarSoC_core0/dout1[54] experiarSoC_core0/dout1[55]
+ experiarSoC_core0/dout1[56] experiarSoC_core0/dout1[57] experiarSoC_core0/dout1[58]
+ experiarSoC_core0/dout1[59] experiarSoC_core0/dout1[60] experiarSoC_core0/dout1[61]
+ experiarSoC_core0/dout1[62] experiarSoC_core0/dout1[63] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_flashSRAM experiarSoC_flashSRAM/din0[0] experiarSoC_flashSRAM/din0[1]
+ experiarSoC_flashSRAM/din0[2] experiarSoC_flashSRAM/din0[3] experiarSoC_flashSRAM/din0[4]
+ experiarSoC_flashSRAM/din0[5] experiarSoC_flashSRAM/din0[6] experiarSoC_flashSRAM/din0[7]
+ experiarSoC_flashSRAM/din0[8] experiarSoC_flashSRAM/din0[9] experiarSoC_flashSRAM/din0[10]
+ experiarSoC_flashSRAM/din0[11] experiarSoC_flashSRAM/din0[12] experiarSoC_flashSRAM/din0[13]
+ experiarSoC_flashSRAM/din0[14] experiarSoC_flashSRAM/din0[15] experiarSoC_flashSRAM/din0[16]
+ experiarSoC_flashSRAM/din0[17] experiarSoC_flashSRAM/din0[18] experiarSoC_flashSRAM/din0[19]
+ experiarSoC_flashSRAM/din0[20] experiarSoC_flashSRAM/din0[21] experiarSoC_flashSRAM/din0[22]
+ experiarSoC_flashSRAM/din0[23] experiarSoC_flashSRAM/din0[24] experiarSoC_flashSRAM/din0[25]
+ experiarSoC_flashSRAM/din0[26] experiarSoC_flashSRAM/din0[27] experiarSoC_flashSRAM/din0[28]
+ experiarSoC_flashSRAM/din0[29] experiarSoC_flashSRAM/din0[30] experiarSoC_flashSRAM/din0[31]
+ experiarSoC_flashSRAM/addr0[0] experiarSoC_flashSRAM/addr0[1] experiarSoC_flashSRAM/addr0[2]
+ experiarSoC_flashSRAM/addr0[3] experiarSoC_flashSRAM/addr0[4] experiarSoC_flashSRAM/addr0[5]
+ experiarSoC_flashSRAM/addr0[6] experiarSoC_flashSRAM/addr0[7] experiarSoC_flashSRAM/addr0[8]
+ experiarSoC_flashSRAM/addr1[0] experiarSoC_flashSRAM/addr1[1] experiarSoC_flashSRAM/addr1[2]
+ experiarSoC_flashSRAM/addr1[3] experiarSoC_flashSRAM/addr1[4] experiarSoC_flashSRAM/addr1[5]
+ experiarSoC_flashSRAM/addr1[6] experiarSoC_flashSRAM/addr1[7] experiarSoC_flashSRAM/addr1[8]
+ experiarSoC_flashSRAM/csb0 experiarSoC_flashSRAM/csb1 experiarSoC_flashSRAM/web0
+ experiarSoC_flashSRAM/clk0 experiarSoC_flashSRAM/clk1 experiarSoC_flashSRAM/wmask0[0]
+ experiarSoC_flashSRAM/wmask0[1] experiarSoC_flashSRAM/wmask0[2] experiarSoC_flashSRAM/wmask0[3]
+ experiarSoC_flashSRAM/dout0[0] experiarSoC_flashSRAM/dout0[1] experiarSoC_flashSRAM/dout0[2]
+ experiarSoC_flashSRAM/dout0[3] experiarSoC_flashSRAM/dout0[4] experiarSoC_flashSRAM/dout0[5]
+ experiarSoC_flashSRAM/dout0[6] experiarSoC_flashSRAM/dout0[7] experiarSoC_flashSRAM/dout0[8]
+ experiarSoC_flashSRAM/dout0[9] experiarSoC_flashSRAM/dout0[10] experiarSoC_flashSRAM/dout0[11]
+ experiarSoC_flashSRAM/dout0[12] experiarSoC_flashSRAM/dout0[13] experiarSoC_flashSRAM/dout0[14]
+ experiarSoC_flashSRAM/dout0[15] experiarSoC_flashSRAM/dout0[16] experiarSoC_flashSRAM/dout0[17]
+ experiarSoC_flashSRAM/dout0[18] experiarSoC_flashSRAM/dout0[19] experiarSoC_flashSRAM/dout0[20]
+ experiarSoC_flashSRAM/dout0[21] experiarSoC_flashSRAM/dout0[22] experiarSoC_flashSRAM/dout0[23]
+ experiarSoC_flashSRAM/dout0[24] experiarSoC_flashSRAM/dout0[25] experiarSoC_flashSRAM/dout0[26]
+ experiarSoC_flashSRAM/dout0[27] experiarSoC_flashSRAM/dout0[28] experiarSoC_flashSRAM/dout0[29]
+ experiarSoC_flashSRAM/dout0[30] experiarSoC_flashSRAM/dout0[31] experiarSoC_flashSRAM/dout1[0]
+ experiarSoC_flashSRAM/dout1[1] experiarSoC_flashSRAM/dout1[2] experiarSoC_flashSRAM/dout1[3]
+ experiarSoC_flashSRAM/dout1[4] experiarSoC_flashSRAM/dout1[5] experiarSoC_flashSRAM/dout1[6]
+ experiarSoC_flashSRAM/dout1[7] experiarSoC_flashSRAM/dout1[8] experiarSoC_flashSRAM/dout1[9]
+ experiarSoC_flashSRAM/dout1[10] experiarSoC_flashSRAM/dout1[11] experiarSoC_flashSRAM/dout1[12]
+ experiarSoC_flashSRAM/dout1[13] experiarSoC_flashSRAM/dout1[14] experiarSoC_flashSRAM/dout1[15]
+ experiarSoC_flashSRAM/dout1[16] experiarSoC_flashSRAM/dout1[17] experiarSoC_flashSRAM/dout1[18]
+ experiarSoC_flashSRAM/dout1[19] experiarSoC_flashSRAM/dout1[20] experiarSoC_flashSRAM/dout1[21]
+ experiarSoC_flashSRAM/dout1[22] experiarSoC_flashSRAM/dout1[23] experiarSoC_flashSRAM/dout1[24]
+ experiarSoC_flashSRAM/dout1[25] experiarSoC_flashSRAM/dout1[26] experiarSoC_flashSRAM/dout1[27]
+ experiarSoC_flashSRAM/dout1[28] experiarSoC_flashSRAM/dout1[29] experiarSoC_flashSRAM/dout1[30]
+ experiarSoC_flashSRAM/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xart vccd1 vssd1 Art
XexperiarSoC_core0 experiarSoC_core0/addr0[0] experiarSoC_core0/addr0[1] experiarSoC_core0/addr0[2]
+ experiarSoC_core0/addr0[3] experiarSoC_core0/addr0[4] experiarSoC_core0/addr0[5]
+ experiarSoC_core0/addr0[6] experiarSoC_core0/addr0[7] experiarSoC_core0/addr0[8]
+ experiarSoC_core0/addr1[0] experiarSoC_core0/addr1[1] experiarSoC_core0/addr1[2]
+ experiarSoC_core0/addr1[3] experiarSoC_core0/addr1[4] experiarSoC_core0/addr1[5]
+ experiarSoC_core0/addr1[6] experiarSoC_core0/addr1[7] experiarSoC_core0/addr1[8]
+ experiarSoC_core0/clk0 experiarSoC_core0/clk1 caravelHost/core0Index[0] caravelHost/core0Index[1]
+ caravelHost/core0Index[2] caravelHost/core0Index[3] caravelHost/core0Index[4] caravelHost/core0Index[5]
+ caravelHost/core0Index[6] caravelHost/core0Index[7] experiarSoC_core0/core_wb_ack_i
+ experiarSoC_core0/core_wb_adr_o[0] experiarSoC_core0/core_wb_adr_o[10] experiarSoC_core0/core_wb_adr_o[11]
+ experiarSoC_core0/core_wb_adr_o[12] experiarSoC_core0/core_wb_adr_o[13] experiarSoC_core0/core_wb_adr_o[14]
+ experiarSoC_core0/core_wb_adr_o[15] experiarSoC_core0/core_wb_adr_o[16] experiarSoC_core0/core_wb_adr_o[17]
+ experiarSoC_core0/core_wb_adr_o[18] experiarSoC_core0/core_wb_adr_o[19] experiarSoC_core0/core_wb_adr_o[1]
+ experiarSoC_core0/core_wb_adr_o[20] experiarSoC_core0/core_wb_adr_o[21] experiarSoC_core0/core_wb_adr_o[22]
+ experiarSoC_core0/core_wb_adr_o[23] experiarSoC_core0/core_wb_adr_o[24] experiarSoC_core0/core_wb_adr_o[25]
+ experiarSoC_core0/core_wb_adr_o[26] experiarSoC_core0/core_wb_adr_o[27] experiarSoC_core0/core_wb_adr_o[2]
+ experiarSoC_core0/core_wb_adr_o[3] experiarSoC_core0/core_wb_adr_o[4] experiarSoC_core0/core_wb_adr_o[5]
+ experiarSoC_core0/core_wb_adr_o[6] experiarSoC_core0/core_wb_adr_o[7] experiarSoC_core0/core_wb_adr_o[8]
+ experiarSoC_core0/core_wb_adr_o[9] experiarSoC_core0/core_wb_cyc_o experiarSoC_core0/core_wb_data_i[0]
+ experiarSoC_core0/core_wb_data_i[10] experiarSoC_core0/core_wb_data_i[11] experiarSoC_core0/core_wb_data_i[12]
+ experiarSoC_core0/core_wb_data_i[13] experiarSoC_core0/core_wb_data_i[14] experiarSoC_core0/core_wb_data_i[15]
+ experiarSoC_core0/core_wb_data_i[16] experiarSoC_core0/core_wb_data_i[17] experiarSoC_core0/core_wb_data_i[18]
+ experiarSoC_core0/core_wb_data_i[19] experiarSoC_core0/core_wb_data_i[1] experiarSoC_core0/core_wb_data_i[20]
+ experiarSoC_core0/core_wb_data_i[21] experiarSoC_core0/core_wb_data_i[22] experiarSoC_core0/core_wb_data_i[23]
+ experiarSoC_core0/core_wb_data_i[24] experiarSoC_core0/core_wb_data_i[25] experiarSoC_core0/core_wb_data_i[26]
+ experiarSoC_core0/core_wb_data_i[27] experiarSoC_core0/core_wb_data_i[28] experiarSoC_core0/core_wb_data_i[29]
+ experiarSoC_core0/core_wb_data_i[2] experiarSoC_core0/core_wb_data_i[30] experiarSoC_core0/core_wb_data_i[31]
+ experiarSoC_core0/core_wb_data_i[3] experiarSoC_core0/core_wb_data_i[4] experiarSoC_core0/core_wb_data_i[5]
+ experiarSoC_core0/core_wb_data_i[6] experiarSoC_core0/core_wb_data_i[7] experiarSoC_core0/core_wb_data_i[8]
+ experiarSoC_core0/core_wb_data_i[9] experiarSoC_core0/core_wb_data_o[0] experiarSoC_core0/core_wb_data_o[10]
+ experiarSoC_core0/core_wb_data_o[11] experiarSoC_core0/core_wb_data_o[12] experiarSoC_core0/core_wb_data_o[13]
+ experiarSoC_core0/core_wb_data_o[14] experiarSoC_core0/core_wb_data_o[15] experiarSoC_core0/core_wb_data_o[16]
+ experiarSoC_core0/core_wb_data_o[17] experiarSoC_core0/core_wb_data_o[18] experiarSoC_core0/core_wb_data_o[19]
+ experiarSoC_core0/core_wb_data_o[1] experiarSoC_core0/core_wb_data_o[20] experiarSoC_core0/core_wb_data_o[21]
+ experiarSoC_core0/core_wb_data_o[22] experiarSoC_core0/core_wb_data_o[23] experiarSoC_core0/core_wb_data_o[24]
+ experiarSoC_core0/core_wb_data_o[25] experiarSoC_core0/core_wb_data_o[26] experiarSoC_core0/core_wb_data_o[27]
+ experiarSoC_core0/core_wb_data_o[28] experiarSoC_core0/core_wb_data_o[29] experiarSoC_core0/core_wb_data_o[2]
+ experiarSoC_core0/core_wb_data_o[30] experiarSoC_core0/core_wb_data_o[31] experiarSoC_core0/core_wb_data_o[3]
+ experiarSoC_core0/core_wb_data_o[4] experiarSoC_core0/core_wb_data_o[5] experiarSoC_core0/core_wb_data_o[6]
+ experiarSoC_core0/core_wb_data_o[7] experiarSoC_core0/core_wb_data_o[8] experiarSoC_core0/core_wb_data_o[9]
+ experiarSoC_core0/core_wb_error_i experiarSoC_core0/core_wb_sel_o[0] experiarSoC_core0/core_wb_sel_o[1]
+ experiarSoC_core0/core_wb_sel_o[2] experiarSoC_core0/core_wb_sel_o[3] experiarSoC_core0/core_wb_stall_i
+ experiarSoC_core0/core_wb_stb_o experiarSoC_core0/core_wb_we_o experiarSoC_core0/csb0[0]
+ experiarSoC_core0/csb0[1] experiarSoC_core0/csb1[0] experiarSoC_core0/csb1[1] experiarSoC_core0/din0[0]
+ experiarSoC_core0/din0[10] experiarSoC_core0/din0[11] experiarSoC_core0/din0[12]
+ experiarSoC_core0/din0[13] experiarSoC_core0/din0[14] experiarSoC_core0/din0[15]
+ experiarSoC_core0/din0[16] experiarSoC_core0/din0[17] experiarSoC_core0/din0[18]
+ experiarSoC_core0/din0[19] experiarSoC_core0/din0[1] experiarSoC_core0/din0[20]
+ experiarSoC_core0/din0[21] experiarSoC_core0/din0[22] experiarSoC_core0/din0[23]
+ experiarSoC_core0/din0[24] experiarSoC_core0/din0[25] experiarSoC_core0/din0[26]
+ experiarSoC_core0/din0[27] experiarSoC_core0/din0[28] experiarSoC_core0/din0[29]
+ experiarSoC_core0/din0[2] experiarSoC_core0/din0[30] experiarSoC_core0/din0[31]
+ experiarSoC_core0/din0[3] experiarSoC_core0/din0[4] experiarSoC_core0/din0[5] experiarSoC_core0/din0[6]
+ experiarSoC_core0/din0[7] experiarSoC_core0/din0[8] experiarSoC_core0/din0[9] experiarSoC_core0/dout0[0]
+ experiarSoC_core0/dout0[10] experiarSoC_core0/dout0[11] experiarSoC_core0/dout0[12]
+ experiarSoC_core0/dout0[13] experiarSoC_core0/dout0[14] experiarSoC_core0/dout0[15]
+ experiarSoC_core0/dout0[16] experiarSoC_core0/dout0[17] experiarSoC_core0/dout0[18]
+ experiarSoC_core0/dout0[19] experiarSoC_core0/dout0[1] experiarSoC_core0/dout0[20]
+ experiarSoC_core0/dout0[21] experiarSoC_core0/dout0[22] experiarSoC_core0/dout0[23]
+ experiarSoC_core0/dout0[24] experiarSoC_core0/dout0[25] experiarSoC_core0/dout0[26]
+ experiarSoC_core0/dout0[27] experiarSoC_core0/dout0[28] experiarSoC_core0/dout0[29]
+ experiarSoC_core0/dout0[2] experiarSoC_core0/dout0[30] experiarSoC_core0/dout0[31]
+ experiarSoC_core0/dout0[32] experiarSoC_core0/dout0[33] experiarSoC_core0/dout0[34]
+ experiarSoC_core0/dout0[35] experiarSoC_core0/dout0[36] experiarSoC_core0/dout0[37]
+ experiarSoC_core0/dout0[38] experiarSoC_core0/dout0[39] experiarSoC_core0/dout0[3]
+ experiarSoC_core0/dout0[40] experiarSoC_core0/dout0[41] experiarSoC_core0/dout0[42]
+ experiarSoC_core0/dout0[43] experiarSoC_core0/dout0[44] experiarSoC_core0/dout0[45]
+ experiarSoC_core0/dout0[46] experiarSoC_core0/dout0[47] experiarSoC_core0/dout0[48]
+ experiarSoC_core0/dout0[49] experiarSoC_core0/dout0[4] experiarSoC_core0/dout0[50]
+ experiarSoC_core0/dout0[51] experiarSoC_core0/dout0[52] experiarSoC_core0/dout0[53]
+ experiarSoC_core0/dout0[54] experiarSoC_core0/dout0[55] experiarSoC_core0/dout0[56]
+ experiarSoC_core0/dout0[57] experiarSoC_core0/dout0[58] experiarSoC_core0/dout0[59]
+ experiarSoC_core0/dout0[5] experiarSoC_core0/dout0[60] experiarSoC_core0/dout0[61]
+ experiarSoC_core0/dout0[62] experiarSoC_core0/dout0[63] experiarSoC_core0/dout0[6]
+ experiarSoC_core0/dout0[7] experiarSoC_core0/dout0[8] experiarSoC_core0/dout0[9]
+ experiarSoC_core0/dout1[0] experiarSoC_core0/dout1[10] experiarSoC_core0/dout1[11]
+ experiarSoC_core0/dout1[12] experiarSoC_core0/dout1[13] experiarSoC_core0/dout1[14]
+ experiarSoC_core0/dout1[15] experiarSoC_core0/dout1[16] experiarSoC_core0/dout1[17]
+ experiarSoC_core0/dout1[18] experiarSoC_core0/dout1[19] experiarSoC_core0/dout1[1]
+ experiarSoC_core0/dout1[20] experiarSoC_core0/dout1[21] experiarSoC_core0/dout1[22]
+ experiarSoC_core0/dout1[23] experiarSoC_core0/dout1[24] experiarSoC_core0/dout1[25]
+ experiarSoC_core0/dout1[26] experiarSoC_core0/dout1[27] experiarSoC_core0/dout1[28]
+ experiarSoC_core0/dout1[29] experiarSoC_core0/dout1[2] experiarSoC_core0/dout1[30]
+ experiarSoC_core0/dout1[31] experiarSoC_core0/dout1[32] experiarSoC_core0/dout1[33]
+ experiarSoC_core0/dout1[34] experiarSoC_core0/dout1[35] experiarSoC_core0/dout1[36]
+ experiarSoC_core0/dout1[37] experiarSoC_core0/dout1[38] experiarSoC_core0/dout1[39]
+ experiarSoC_core0/dout1[3] experiarSoC_core0/dout1[40] experiarSoC_core0/dout1[41]
+ experiarSoC_core0/dout1[42] experiarSoC_core0/dout1[43] experiarSoC_core0/dout1[44]
+ experiarSoC_core0/dout1[45] experiarSoC_core0/dout1[46] experiarSoC_core0/dout1[47]
+ experiarSoC_core0/dout1[48] experiarSoC_core0/dout1[49] experiarSoC_core0/dout1[4]
+ experiarSoC_core0/dout1[50] experiarSoC_core0/dout1[51] experiarSoC_core0/dout1[52]
+ experiarSoC_core0/dout1[53] experiarSoC_core0/dout1[54] experiarSoC_core0/dout1[55]
+ experiarSoC_core0/dout1[56] experiarSoC_core0/dout1[57] experiarSoC_core0/dout1[58]
+ experiarSoC_core0/dout1[59] experiarSoC_core0/dout1[5] experiarSoC_core0/dout1[60]
+ experiarSoC_core0/dout1[61] experiarSoC_core0/dout1[62] experiarSoC_core0/dout1[63]
+ experiarSoC_core0/dout1[6] experiarSoC_core0/dout1[7] experiarSoC_core0/dout1[8]
+ experiarSoC_core0/dout1[9] experiarSoC_core1/irq[0] experiarSoC_core1/irq[10] experiarSoC_core1/irq[11]
+ experiarSoC_core1/irq[12] experiarSoC_core1/irq[13] experiarSoC_core1/irq[14] experiarSoC_core1/irq[15]
+ experiarSoC_core1/irq[1] experiarSoC_core1/irq[2] experiarSoC_core1/irq[3] experiarSoC_core1/irq[4]
+ experiarSoC_core1/irq[5] experiarSoC_core1/irq[6] experiarSoC_core1/irq[7] experiarSoC_core1/irq[8]
+ experiarSoC_core1/irq[9] experiarSoC_core1/jtag_tck experiarSoC_core0/jtag_tdi experiarSoC_core1/jtag_tdi
+ experiarSoC_core1/jtag_tms experiarSoC_core0/localMemory_wb_ack_o experiarSoC_core0/localMemory_wb_adr_i[0]
+ experiarSoC_core0/localMemory_wb_adr_i[10] experiarSoC_core0/localMemory_wb_adr_i[11]
+ experiarSoC_core0/localMemory_wb_adr_i[12] experiarSoC_core0/localMemory_wb_adr_i[13]
+ experiarSoC_core0/localMemory_wb_adr_i[14] experiarSoC_core0/localMemory_wb_adr_i[15]
+ experiarSoC_core0/localMemory_wb_adr_i[16] experiarSoC_core0/localMemory_wb_adr_i[17]
+ experiarSoC_core0/localMemory_wb_adr_i[18] experiarSoC_core0/localMemory_wb_adr_i[19]
+ experiarSoC_core0/localMemory_wb_adr_i[1] experiarSoC_core0/localMemory_wb_adr_i[20]
+ experiarSoC_core0/localMemory_wb_adr_i[21] experiarSoC_core0/localMemory_wb_adr_i[22]
+ experiarSoC_core0/localMemory_wb_adr_i[23] experiarSoC_core0/localMemory_wb_adr_i[2]
+ experiarSoC_core0/localMemory_wb_adr_i[3] experiarSoC_core0/localMemory_wb_adr_i[4]
+ experiarSoC_core0/localMemory_wb_adr_i[5] experiarSoC_core0/localMemory_wb_adr_i[6]
+ experiarSoC_core0/localMemory_wb_adr_i[7] experiarSoC_core0/localMemory_wb_adr_i[8]
+ experiarSoC_core0/localMemory_wb_adr_i[9] experiarSoC_core0/localMemory_wb_cyc_i
+ experiarSoC_core0/localMemory_wb_data_i[0] experiarSoC_core0/localMemory_wb_data_i[10]
+ experiarSoC_core0/localMemory_wb_data_i[11] experiarSoC_core0/localMemory_wb_data_i[12]
+ experiarSoC_core0/localMemory_wb_data_i[13] experiarSoC_core0/localMemory_wb_data_i[14]
+ experiarSoC_core0/localMemory_wb_data_i[15] experiarSoC_core0/localMemory_wb_data_i[16]
+ experiarSoC_core0/localMemory_wb_data_i[17] experiarSoC_core0/localMemory_wb_data_i[18]
+ experiarSoC_core0/localMemory_wb_data_i[19] experiarSoC_core0/localMemory_wb_data_i[1]
+ experiarSoC_core0/localMemory_wb_data_i[20] experiarSoC_core0/localMemory_wb_data_i[21]
+ experiarSoC_core0/localMemory_wb_data_i[22] experiarSoC_core0/localMemory_wb_data_i[23]
+ experiarSoC_core0/localMemory_wb_data_i[24] experiarSoC_core0/localMemory_wb_data_i[25]
+ experiarSoC_core0/localMemory_wb_data_i[26] experiarSoC_core0/localMemory_wb_data_i[27]
+ experiarSoC_core0/localMemory_wb_data_i[28] experiarSoC_core0/localMemory_wb_data_i[29]
+ experiarSoC_core0/localMemory_wb_data_i[2] experiarSoC_core0/localMemory_wb_data_i[30]
+ experiarSoC_core0/localMemory_wb_data_i[31] experiarSoC_core0/localMemory_wb_data_i[3]
+ experiarSoC_core0/localMemory_wb_data_i[4] experiarSoC_core0/localMemory_wb_data_i[5]
+ experiarSoC_core0/localMemory_wb_data_i[6] experiarSoC_core0/localMemory_wb_data_i[7]
+ experiarSoC_core0/localMemory_wb_data_i[8] experiarSoC_core0/localMemory_wb_data_i[9]
+ experiarSoC_core0/localMemory_wb_data_o[0] experiarSoC_core0/localMemory_wb_data_o[10]
+ experiarSoC_core0/localMemory_wb_data_o[11] experiarSoC_core0/localMemory_wb_data_o[12]
+ experiarSoC_core0/localMemory_wb_data_o[13] experiarSoC_core0/localMemory_wb_data_o[14]
+ experiarSoC_core0/localMemory_wb_data_o[15] experiarSoC_core0/localMemory_wb_data_o[16]
+ experiarSoC_core0/localMemory_wb_data_o[17] experiarSoC_core0/localMemory_wb_data_o[18]
+ experiarSoC_core0/localMemory_wb_data_o[19] experiarSoC_core0/localMemory_wb_data_o[1]
+ experiarSoC_core0/localMemory_wb_data_o[20] experiarSoC_core0/localMemory_wb_data_o[21]
+ experiarSoC_core0/localMemory_wb_data_o[22] experiarSoC_core0/localMemory_wb_data_o[23]
+ experiarSoC_core0/localMemory_wb_data_o[24] experiarSoC_core0/localMemory_wb_data_o[25]
+ experiarSoC_core0/localMemory_wb_data_o[26] experiarSoC_core0/localMemory_wb_data_o[27]
+ experiarSoC_core0/localMemory_wb_data_o[28] experiarSoC_core0/localMemory_wb_data_o[29]
+ experiarSoC_core0/localMemory_wb_data_o[2] experiarSoC_core0/localMemory_wb_data_o[30]
+ experiarSoC_core0/localMemory_wb_data_o[31] experiarSoC_core0/localMemory_wb_data_o[3]
+ experiarSoC_core0/localMemory_wb_data_o[4] experiarSoC_core0/localMemory_wb_data_o[5]
+ experiarSoC_core0/localMemory_wb_data_o[6] experiarSoC_core0/localMemory_wb_data_o[7]
+ experiarSoC_core0/localMemory_wb_data_o[8] experiarSoC_core0/localMemory_wb_data_o[9]
+ experiarSoC_core0/localMemory_wb_error_o experiarSoC_core0/localMemory_wb_sel_i[0]
+ experiarSoC_core0/localMemory_wb_sel_i[1] experiarSoC_core0/localMemory_wb_sel_i[2]
+ experiarSoC_core0/localMemory_wb_sel_i[3] experiarSoC_core0/localMemory_wb_stall_o
+ experiarSoC_core0/localMemory_wb_stb_i experiarSoC_core0/localMemory_wb_we_i caravelHost/manufacturerID[0]
+ caravelHost/manufacturerID[10] caravelHost/manufacturerID[1] caravelHost/manufacturerID[2]
+ caravelHost/manufacturerID[3] caravelHost/manufacturerID[4] caravelHost/manufacturerID[5]
+ caravelHost/manufacturerID[6] caravelHost/manufacturerID[7] caravelHost/manufacturerID[8]
+ caravelHost/manufacturerID[9] caravelHost/partID[0] caravelHost/partID[10] caravelHost/partID[11]
+ caravelHost/partID[12] caravelHost/partID[13] caravelHost/partID[14] caravelHost/partID[15]
+ caravelHost/partID[1] caravelHost/partID[2] caravelHost/partID[3] caravelHost/partID[4]
+ caravelHost/partID[5] caravelHost/partID[6] caravelHost/partID[7] caravelHost/partID[8]
+ caravelHost/partID[9] la_data_out[69] la_data_out[70] la_data_out[28] la_data_out[29]
+ la_data_out[27] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[18]
+ la_data_out[19] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[38] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[39] la_data_out[67]
+ la_data_out[68] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[71] la_data_out[72]
+ la_data_out[26] vccd1 caravelHost/versionID[0] caravelHost/versionID[1] caravelHost/versionID[2]
+ caravelHost/versionID[3] vssd1 wb_clk_i wb_rst_i experiarSoC_core0/web0 experiarSoC_core0/wmask0[0]
+ experiarSoC_core0/wmask0[1] experiarSoC_core0/wmask0[2] experiarSoC_core0/wmask0[3]
+ ExperiarCore
XexperiarSoC_core1 experiarSoC_core1/addr0[0] experiarSoC_core1/addr0[1] experiarSoC_core1/addr0[2]
+ experiarSoC_core1/addr0[3] experiarSoC_core1/addr0[4] experiarSoC_core1/addr0[5]
+ experiarSoC_core1/addr0[6] experiarSoC_core1/addr0[7] experiarSoC_core1/addr0[8]
+ experiarSoC_core1/addr1[0] experiarSoC_core1/addr1[1] experiarSoC_core1/addr1[2]
+ experiarSoC_core1/addr1[3] experiarSoC_core1/addr1[4] experiarSoC_core1/addr1[5]
+ experiarSoC_core1/addr1[6] experiarSoC_core1/addr1[7] experiarSoC_core1/addr1[8]
+ experiarSoC_core1/clk0 experiarSoC_core1/clk1 caravelHost/core1Index[0] caravelHost/core1Index[1]
+ caravelHost/core1Index[2] caravelHost/core1Index[3] caravelHost/core1Index[4] caravelHost/core1Index[5]
+ caravelHost/core1Index[6] caravelHost/core1Index[7] experiarSoC_core1/core_wb_ack_i
+ experiarSoC_core1/core_wb_adr_o[0] experiarSoC_core1/core_wb_adr_o[10] experiarSoC_core1/core_wb_adr_o[11]
+ experiarSoC_core1/core_wb_adr_o[12] experiarSoC_core1/core_wb_adr_o[13] experiarSoC_core1/core_wb_adr_o[14]
+ experiarSoC_core1/core_wb_adr_o[15] experiarSoC_core1/core_wb_adr_o[16] experiarSoC_core1/core_wb_adr_o[17]
+ experiarSoC_core1/core_wb_adr_o[18] experiarSoC_core1/core_wb_adr_o[19] experiarSoC_core1/core_wb_adr_o[1]
+ experiarSoC_core1/core_wb_adr_o[20] experiarSoC_core1/core_wb_adr_o[21] experiarSoC_core1/core_wb_adr_o[22]
+ experiarSoC_core1/core_wb_adr_o[23] experiarSoC_core1/core_wb_adr_o[24] experiarSoC_core1/core_wb_adr_o[25]
+ experiarSoC_core1/core_wb_adr_o[26] experiarSoC_core1/core_wb_adr_o[27] experiarSoC_core1/core_wb_adr_o[2]
+ experiarSoC_core1/core_wb_adr_o[3] experiarSoC_core1/core_wb_adr_o[4] experiarSoC_core1/core_wb_adr_o[5]
+ experiarSoC_core1/core_wb_adr_o[6] experiarSoC_core1/core_wb_adr_o[7] experiarSoC_core1/core_wb_adr_o[8]
+ experiarSoC_core1/core_wb_adr_o[9] experiarSoC_core1/core_wb_cyc_o experiarSoC_core1/core_wb_data_i[0]
+ experiarSoC_core1/core_wb_data_i[10] experiarSoC_core1/core_wb_data_i[11] experiarSoC_core1/core_wb_data_i[12]
+ experiarSoC_core1/core_wb_data_i[13] experiarSoC_core1/core_wb_data_i[14] experiarSoC_core1/core_wb_data_i[15]
+ experiarSoC_core1/core_wb_data_i[16] experiarSoC_core1/core_wb_data_i[17] experiarSoC_core1/core_wb_data_i[18]
+ experiarSoC_core1/core_wb_data_i[19] experiarSoC_core1/core_wb_data_i[1] experiarSoC_core1/core_wb_data_i[20]
+ experiarSoC_core1/core_wb_data_i[21] experiarSoC_core1/core_wb_data_i[22] experiarSoC_core1/core_wb_data_i[23]
+ experiarSoC_core1/core_wb_data_i[24] experiarSoC_core1/core_wb_data_i[25] experiarSoC_core1/core_wb_data_i[26]
+ experiarSoC_core1/core_wb_data_i[27] experiarSoC_core1/core_wb_data_i[28] experiarSoC_core1/core_wb_data_i[29]
+ experiarSoC_core1/core_wb_data_i[2] experiarSoC_core1/core_wb_data_i[30] experiarSoC_core1/core_wb_data_i[31]
+ experiarSoC_core1/core_wb_data_i[3] experiarSoC_core1/core_wb_data_i[4] experiarSoC_core1/core_wb_data_i[5]
+ experiarSoC_core1/core_wb_data_i[6] experiarSoC_core1/core_wb_data_i[7] experiarSoC_core1/core_wb_data_i[8]
+ experiarSoC_core1/core_wb_data_i[9] experiarSoC_core1/core_wb_data_o[0] experiarSoC_core1/core_wb_data_o[10]
+ experiarSoC_core1/core_wb_data_o[11] experiarSoC_core1/core_wb_data_o[12] experiarSoC_core1/core_wb_data_o[13]
+ experiarSoC_core1/core_wb_data_o[14] experiarSoC_core1/core_wb_data_o[15] experiarSoC_core1/core_wb_data_o[16]
+ experiarSoC_core1/core_wb_data_o[17] experiarSoC_core1/core_wb_data_o[18] experiarSoC_core1/core_wb_data_o[19]
+ experiarSoC_core1/core_wb_data_o[1] experiarSoC_core1/core_wb_data_o[20] experiarSoC_core1/core_wb_data_o[21]
+ experiarSoC_core1/core_wb_data_o[22] experiarSoC_core1/core_wb_data_o[23] experiarSoC_core1/core_wb_data_o[24]
+ experiarSoC_core1/core_wb_data_o[25] experiarSoC_core1/core_wb_data_o[26] experiarSoC_core1/core_wb_data_o[27]
+ experiarSoC_core1/core_wb_data_o[28] experiarSoC_core1/core_wb_data_o[29] experiarSoC_core1/core_wb_data_o[2]
+ experiarSoC_core1/core_wb_data_o[30] experiarSoC_core1/core_wb_data_o[31] experiarSoC_core1/core_wb_data_o[3]
+ experiarSoC_core1/core_wb_data_o[4] experiarSoC_core1/core_wb_data_o[5] experiarSoC_core1/core_wb_data_o[6]
+ experiarSoC_core1/core_wb_data_o[7] experiarSoC_core1/core_wb_data_o[8] experiarSoC_core1/core_wb_data_o[9]
+ experiarSoC_core1/core_wb_error_i experiarSoC_core1/core_wb_sel_o[0] experiarSoC_core1/core_wb_sel_o[1]
+ experiarSoC_core1/core_wb_sel_o[2] experiarSoC_core1/core_wb_sel_o[3] experiarSoC_core1/core_wb_stall_i
+ experiarSoC_core1/core_wb_stb_o experiarSoC_core1/core_wb_we_o experiarSoC_core1/csb0[0]
+ experiarSoC_core1/csb0[1] experiarSoC_core1/csb1[0] experiarSoC_core1/csb1[1] experiarSoC_core1/din0[0]
+ experiarSoC_core1/din0[10] experiarSoC_core1/din0[11] experiarSoC_core1/din0[12]
+ experiarSoC_core1/din0[13] experiarSoC_core1/din0[14] experiarSoC_core1/din0[15]
+ experiarSoC_core1/din0[16] experiarSoC_core1/din0[17] experiarSoC_core1/din0[18]
+ experiarSoC_core1/din0[19] experiarSoC_core1/din0[1] experiarSoC_core1/din0[20]
+ experiarSoC_core1/din0[21] experiarSoC_core1/din0[22] experiarSoC_core1/din0[23]
+ experiarSoC_core1/din0[24] experiarSoC_core1/din0[25] experiarSoC_core1/din0[26]
+ experiarSoC_core1/din0[27] experiarSoC_core1/din0[28] experiarSoC_core1/din0[29]
+ experiarSoC_core1/din0[2] experiarSoC_core1/din0[30] experiarSoC_core1/din0[31]
+ experiarSoC_core1/din0[3] experiarSoC_core1/din0[4] experiarSoC_core1/din0[5] experiarSoC_core1/din0[6]
+ experiarSoC_core1/din0[7] experiarSoC_core1/din0[8] experiarSoC_core1/din0[9] experiarSoC_core1/dout0[0]
+ experiarSoC_core1/dout0[10] experiarSoC_core1/dout0[11] experiarSoC_core1/dout0[12]
+ experiarSoC_core1/dout0[13] experiarSoC_core1/dout0[14] experiarSoC_core1/dout0[15]
+ experiarSoC_core1/dout0[16] experiarSoC_core1/dout0[17] experiarSoC_core1/dout0[18]
+ experiarSoC_core1/dout0[19] experiarSoC_core1/dout0[1] experiarSoC_core1/dout0[20]
+ experiarSoC_core1/dout0[21] experiarSoC_core1/dout0[22] experiarSoC_core1/dout0[23]
+ experiarSoC_core1/dout0[24] experiarSoC_core1/dout0[25] experiarSoC_core1/dout0[26]
+ experiarSoC_core1/dout0[27] experiarSoC_core1/dout0[28] experiarSoC_core1/dout0[29]
+ experiarSoC_core1/dout0[2] experiarSoC_core1/dout0[30] experiarSoC_core1/dout0[31]
+ experiarSoC_core1/dout0[32] experiarSoC_core1/dout0[33] experiarSoC_core1/dout0[34]
+ experiarSoC_core1/dout0[35] experiarSoC_core1/dout0[36] experiarSoC_core1/dout0[37]
+ experiarSoC_core1/dout0[38] experiarSoC_core1/dout0[39] experiarSoC_core1/dout0[3]
+ experiarSoC_core1/dout0[40] experiarSoC_core1/dout0[41] experiarSoC_core1/dout0[42]
+ experiarSoC_core1/dout0[43] experiarSoC_core1/dout0[44] experiarSoC_core1/dout0[45]
+ experiarSoC_core1/dout0[46] experiarSoC_core1/dout0[47] experiarSoC_core1/dout0[48]
+ experiarSoC_core1/dout0[49] experiarSoC_core1/dout0[4] experiarSoC_core1/dout0[50]
+ experiarSoC_core1/dout0[51] experiarSoC_core1/dout0[52] experiarSoC_core1/dout0[53]
+ experiarSoC_core1/dout0[54] experiarSoC_core1/dout0[55] experiarSoC_core1/dout0[56]
+ experiarSoC_core1/dout0[57] experiarSoC_core1/dout0[58] experiarSoC_core1/dout0[59]
+ experiarSoC_core1/dout0[5] experiarSoC_core1/dout0[60] experiarSoC_core1/dout0[61]
+ experiarSoC_core1/dout0[62] experiarSoC_core1/dout0[63] experiarSoC_core1/dout0[6]
+ experiarSoC_core1/dout0[7] experiarSoC_core1/dout0[8] experiarSoC_core1/dout0[9]
+ experiarSoC_core1/dout1[0] experiarSoC_core1/dout1[10] experiarSoC_core1/dout1[11]
+ experiarSoC_core1/dout1[12] experiarSoC_core1/dout1[13] experiarSoC_core1/dout1[14]
+ experiarSoC_core1/dout1[15] experiarSoC_core1/dout1[16] experiarSoC_core1/dout1[17]
+ experiarSoC_core1/dout1[18] experiarSoC_core1/dout1[19] experiarSoC_core1/dout1[1]
+ experiarSoC_core1/dout1[20] experiarSoC_core1/dout1[21] experiarSoC_core1/dout1[22]
+ experiarSoC_core1/dout1[23] experiarSoC_core1/dout1[24] experiarSoC_core1/dout1[25]
+ experiarSoC_core1/dout1[26] experiarSoC_core1/dout1[27] experiarSoC_core1/dout1[28]
+ experiarSoC_core1/dout1[29] experiarSoC_core1/dout1[2] experiarSoC_core1/dout1[30]
+ experiarSoC_core1/dout1[31] experiarSoC_core1/dout1[32] experiarSoC_core1/dout1[33]
+ experiarSoC_core1/dout1[34] experiarSoC_core1/dout1[35] experiarSoC_core1/dout1[36]
+ experiarSoC_core1/dout1[37] experiarSoC_core1/dout1[38] experiarSoC_core1/dout1[39]
+ experiarSoC_core1/dout1[3] experiarSoC_core1/dout1[40] experiarSoC_core1/dout1[41]
+ experiarSoC_core1/dout1[42] experiarSoC_core1/dout1[43] experiarSoC_core1/dout1[44]
+ experiarSoC_core1/dout1[45] experiarSoC_core1/dout1[46] experiarSoC_core1/dout1[47]
+ experiarSoC_core1/dout1[48] experiarSoC_core1/dout1[49] experiarSoC_core1/dout1[4]
+ experiarSoC_core1/dout1[50] experiarSoC_core1/dout1[51] experiarSoC_core1/dout1[52]
+ experiarSoC_core1/dout1[53] experiarSoC_core1/dout1[54] experiarSoC_core1/dout1[55]
+ experiarSoC_core1/dout1[56] experiarSoC_core1/dout1[57] experiarSoC_core1/dout1[58]
+ experiarSoC_core1/dout1[59] experiarSoC_core1/dout1[5] experiarSoC_core1/dout1[60]
+ experiarSoC_core1/dout1[61] experiarSoC_core1/dout1[62] experiarSoC_core1/dout1[63]
+ experiarSoC_core1/dout1[6] experiarSoC_core1/dout1[7] experiarSoC_core1/dout1[8]
+ experiarSoC_core1/dout1[9] experiarSoC_core1/irq[0] experiarSoC_core1/irq[10] experiarSoC_core1/irq[11]
+ experiarSoC_core1/irq[12] experiarSoC_core1/irq[13] experiarSoC_core1/irq[14] experiarSoC_core1/irq[15]
+ experiarSoC_core1/irq[1] experiarSoC_core1/irq[2] experiarSoC_core1/irq[3] experiarSoC_core1/irq[4]
+ experiarSoC_core1/irq[5] experiarSoC_core1/irq[6] experiarSoC_core1/irq[7] experiarSoC_core1/irq[8]
+ experiarSoC_core1/irq[9] experiarSoC_core1/jtag_tck experiarSoC_core1/jtag_tdi experiarSoC_core1/jtag_tdo
+ experiarSoC_core1/jtag_tms experiarSoC_core1/localMemory_wb_ack_o experiarSoC_core1/localMemory_wb_adr_i[0]
+ experiarSoC_core1/localMemory_wb_adr_i[10] experiarSoC_core1/localMemory_wb_adr_i[11]
+ experiarSoC_core1/localMemory_wb_adr_i[12] experiarSoC_core1/localMemory_wb_adr_i[13]
+ experiarSoC_core1/localMemory_wb_adr_i[14] experiarSoC_core1/localMemory_wb_adr_i[15]
+ experiarSoC_core1/localMemory_wb_adr_i[16] experiarSoC_core1/localMemory_wb_adr_i[17]
+ experiarSoC_core1/localMemory_wb_adr_i[18] experiarSoC_core1/localMemory_wb_adr_i[19]
+ experiarSoC_core1/localMemory_wb_adr_i[1] experiarSoC_core1/localMemory_wb_adr_i[20]
+ experiarSoC_core1/localMemory_wb_adr_i[21] experiarSoC_core1/localMemory_wb_adr_i[22]
+ experiarSoC_core1/localMemory_wb_adr_i[23] experiarSoC_core1/localMemory_wb_adr_i[2]
+ experiarSoC_core1/localMemory_wb_adr_i[3] experiarSoC_core1/localMemory_wb_adr_i[4]
+ experiarSoC_core1/localMemory_wb_adr_i[5] experiarSoC_core1/localMemory_wb_adr_i[6]
+ experiarSoC_core1/localMemory_wb_adr_i[7] experiarSoC_core1/localMemory_wb_adr_i[8]
+ experiarSoC_core1/localMemory_wb_adr_i[9] experiarSoC_core1/localMemory_wb_cyc_i
+ experiarSoC_core1/localMemory_wb_data_i[0] experiarSoC_core1/localMemory_wb_data_i[10]
+ experiarSoC_core1/localMemory_wb_data_i[11] experiarSoC_core1/localMemory_wb_data_i[12]
+ experiarSoC_core1/localMemory_wb_data_i[13] experiarSoC_core1/localMemory_wb_data_i[14]
+ experiarSoC_core1/localMemory_wb_data_i[15] experiarSoC_core1/localMemory_wb_data_i[16]
+ experiarSoC_core1/localMemory_wb_data_i[17] experiarSoC_core1/localMemory_wb_data_i[18]
+ experiarSoC_core1/localMemory_wb_data_i[19] experiarSoC_core1/localMemory_wb_data_i[1]
+ experiarSoC_core1/localMemory_wb_data_i[20] experiarSoC_core1/localMemory_wb_data_i[21]
+ experiarSoC_core1/localMemory_wb_data_i[22] experiarSoC_core1/localMemory_wb_data_i[23]
+ experiarSoC_core1/localMemory_wb_data_i[24] experiarSoC_core1/localMemory_wb_data_i[25]
+ experiarSoC_core1/localMemory_wb_data_i[26] experiarSoC_core1/localMemory_wb_data_i[27]
+ experiarSoC_core1/localMemory_wb_data_i[28] experiarSoC_core1/localMemory_wb_data_i[29]
+ experiarSoC_core1/localMemory_wb_data_i[2] experiarSoC_core1/localMemory_wb_data_i[30]
+ experiarSoC_core1/localMemory_wb_data_i[31] experiarSoC_core1/localMemory_wb_data_i[3]
+ experiarSoC_core1/localMemory_wb_data_i[4] experiarSoC_core1/localMemory_wb_data_i[5]
+ experiarSoC_core1/localMemory_wb_data_i[6] experiarSoC_core1/localMemory_wb_data_i[7]
+ experiarSoC_core1/localMemory_wb_data_i[8] experiarSoC_core1/localMemory_wb_data_i[9]
+ experiarSoC_core1/localMemory_wb_data_o[0] experiarSoC_core1/localMemory_wb_data_o[10]
+ experiarSoC_core1/localMemory_wb_data_o[11] experiarSoC_core1/localMemory_wb_data_o[12]
+ experiarSoC_core1/localMemory_wb_data_o[13] experiarSoC_core1/localMemory_wb_data_o[14]
+ experiarSoC_core1/localMemory_wb_data_o[15] experiarSoC_core1/localMemory_wb_data_o[16]
+ experiarSoC_core1/localMemory_wb_data_o[17] experiarSoC_core1/localMemory_wb_data_o[18]
+ experiarSoC_core1/localMemory_wb_data_o[19] experiarSoC_core1/localMemory_wb_data_o[1]
+ experiarSoC_core1/localMemory_wb_data_o[20] experiarSoC_core1/localMemory_wb_data_o[21]
+ experiarSoC_core1/localMemory_wb_data_o[22] experiarSoC_core1/localMemory_wb_data_o[23]
+ experiarSoC_core1/localMemory_wb_data_o[24] experiarSoC_core1/localMemory_wb_data_o[25]
+ experiarSoC_core1/localMemory_wb_data_o[26] experiarSoC_core1/localMemory_wb_data_o[27]
+ experiarSoC_core1/localMemory_wb_data_o[28] experiarSoC_core1/localMemory_wb_data_o[29]
+ experiarSoC_core1/localMemory_wb_data_o[2] experiarSoC_core1/localMemory_wb_data_o[30]
+ experiarSoC_core1/localMemory_wb_data_o[31] experiarSoC_core1/localMemory_wb_data_o[3]
+ experiarSoC_core1/localMemory_wb_data_o[4] experiarSoC_core1/localMemory_wb_data_o[5]
+ experiarSoC_core1/localMemory_wb_data_o[6] experiarSoC_core1/localMemory_wb_data_o[7]
+ experiarSoC_core1/localMemory_wb_data_o[8] experiarSoC_core1/localMemory_wb_data_o[9]
+ experiarSoC_core1/localMemory_wb_error_o experiarSoC_core1/localMemory_wb_sel_i[0]
+ experiarSoC_core1/localMemory_wb_sel_i[1] experiarSoC_core1/localMemory_wb_sel_i[2]
+ experiarSoC_core1/localMemory_wb_sel_i[3] experiarSoC_core1/localMemory_wb_stall_o
+ experiarSoC_core1/localMemory_wb_stb_i experiarSoC_core1/localMemory_wb_we_i caravelHost/manufacturerID[0]
+ caravelHost/manufacturerID[10] caravelHost/manufacturerID[1] caravelHost/manufacturerID[2]
+ caravelHost/manufacturerID[3] caravelHost/manufacturerID[4] caravelHost/manufacturerID[5]
+ caravelHost/manufacturerID[6] caravelHost/manufacturerID[7] caravelHost/manufacturerID[8]
+ caravelHost/manufacturerID[9] caravelHost/partID[0] caravelHost/partID[10] caravelHost/partID[11]
+ caravelHost/partID[12] caravelHost/partID[13] caravelHost/partID[14] caravelHost/partID[15]
+ caravelHost/partID[1] caravelHost/partID[2] caravelHost/partID[3] caravelHost/partID[4]
+ caravelHost/partID[5] caravelHost/partID[6] caravelHost/partID[7] caravelHost/partID[8]
+ caravelHost/partID[9] la_data_out[124] la_data_out[125] la_data_out[83] la_data_out[84]
+ la_data_out[82] la_data_out[78] la_data_out[79] la_data_out[80] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[85]
+ la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[90]
+ la_data_out[91] la_data_out[92] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[110] la_data_out[111] la_data_out[93] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[120] la_data_out[121] la_data_out[94] la_data_out[122]
+ la_data_out[123] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[100] la_data_out[101] la_data_out[126] la_data_out[127]
+ la_data_out[81] vccd1 caravelHost/versionID[0] caravelHost/versionID[1] caravelHost/versionID[2]
+ caravelHost/versionID[3] vssd1 wb_clk_i wb_rst_i experiarSoC_core1/web0 experiarSoC_core1/wmask0[0]
+ experiarSoC_core1/wmask0[1] experiarSoC_core1/wmask0[2] experiarSoC_core1/wmask0[3]
+ ExperiarCore
XexperiarSoC_peripherals experiarSoC_flash/flash_csb experiarSoC_flash/flash_io0_read
+ experiarSoC_flash/flash_io0_we experiarSoC_flash/flash_io0_write experiarSoC_flash/flash_io1_read
+ experiarSoC_flash/flash_io1_we experiarSoC_flash/flash_io1_write experiarSoC_flash/flash_sck
+ caravelHost/caravel_uart_tx caravelHost/caravel_uart_rx io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9]
+ io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16]
+ io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23]
+ io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30]
+ io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] experiarSoC_core1/jtag_tck experiarSoC_core0/jtag_tdi
+ experiarSoC_core1/jtag_tdo experiarSoC_core1/jtag_tms experiarSoC_core1/irq[0] experiarSoC_core1/irq[1]
+ experiarSoC_core1/irq[2] experiarSoC_core1/irq[3] experiarSoC_core1/irq[4] experiarSoC_core1/irq[5]
+ experiarSoC_core1/irq[6] experiarSoC_core1/irq[7] experiarSoC_core1/irq[8] experiarSoC_core1/irq[9]
+ la_data_out[0] la_data_out[1] vccd1 experiarSoC_video/vga_b[0] experiarSoC_video/vga_b[1]
+ experiarSoC_video/vga_g[0] experiarSoC_video/vga_g[1] experiarSoC_video/vga_hsync
+ experiarSoC_video/vga_r[0] experiarSoC_video/vga_r[1] experiarSoC_video/vga_vsync
+ vssd1 experiarSoC_peripherals/wb_ack_o experiarSoC_peripherals/wb_adr_i[0] experiarSoC_peripherals/wb_adr_i[10]
+ experiarSoC_peripherals/wb_adr_i[11] experiarSoC_peripherals/wb_adr_i[12] experiarSoC_peripherals/wb_adr_i[13]
+ experiarSoC_peripherals/wb_adr_i[14] experiarSoC_peripherals/wb_adr_i[15] experiarSoC_peripherals/wb_adr_i[16]
+ experiarSoC_peripherals/wb_adr_i[17] experiarSoC_peripherals/wb_adr_i[18] experiarSoC_peripherals/wb_adr_i[19]
+ experiarSoC_peripherals/wb_adr_i[1] experiarSoC_peripherals/wb_adr_i[20] experiarSoC_peripherals/wb_adr_i[21]
+ experiarSoC_peripherals/wb_adr_i[22] experiarSoC_peripherals/wb_adr_i[23] experiarSoC_peripherals/wb_adr_i[2]
+ experiarSoC_peripherals/wb_adr_i[3] experiarSoC_peripherals/wb_adr_i[4] experiarSoC_peripherals/wb_adr_i[5]
+ experiarSoC_peripherals/wb_adr_i[6] experiarSoC_peripherals/wb_adr_i[7] experiarSoC_peripherals/wb_adr_i[8]
+ experiarSoC_peripherals/wb_adr_i[9] wb_clk_i experiarSoC_peripherals/wb_cyc_i experiarSoC_peripherals/wb_data_i[0]
+ experiarSoC_peripherals/wb_data_i[10] experiarSoC_peripherals/wb_data_i[11] experiarSoC_peripherals/wb_data_i[12]
+ experiarSoC_peripherals/wb_data_i[13] experiarSoC_peripherals/wb_data_i[14] experiarSoC_peripherals/wb_data_i[15]
+ experiarSoC_peripherals/wb_data_i[16] experiarSoC_peripherals/wb_data_i[17] experiarSoC_peripherals/wb_data_i[18]
+ experiarSoC_peripherals/wb_data_i[19] experiarSoC_peripherals/wb_data_i[1] experiarSoC_peripherals/wb_data_i[20]
+ experiarSoC_peripherals/wb_data_i[21] experiarSoC_peripherals/wb_data_i[22] experiarSoC_peripherals/wb_data_i[23]
+ experiarSoC_peripherals/wb_data_i[24] experiarSoC_peripherals/wb_data_i[25] experiarSoC_peripherals/wb_data_i[26]
+ experiarSoC_peripherals/wb_data_i[27] experiarSoC_peripherals/wb_data_i[28] experiarSoC_peripherals/wb_data_i[29]
+ experiarSoC_peripherals/wb_data_i[2] experiarSoC_peripherals/wb_data_i[30] experiarSoC_peripherals/wb_data_i[31]
+ experiarSoC_peripherals/wb_data_i[3] experiarSoC_peripherals/wb_data_i[4] experiarSoC_peripherals/wb_data_i[5]
+ experiarSoC_peripherals/wb_data_i[6] experiarSoC_peripherals/wb_data_i[7] experiarSoC_peripherals/wb_data_i[8]
+ experiarSoC_peripherals/wb_data_i[9] experiarSoC_peripherals/wb_data_o[0] experiarSoC_peripherals/wb_data_o[10]
+ experiarSoC_peripherals/wb_data_o[11] experiarSoC_peripherals/wb_data_o[12] experiarSoC_peripherals/wb_data_o[13]
+ experiarSoC_peripherals/wb_data_o[14] experiarSoC_peripherals/wb_data_o[15] experiarSoC_peripherals/wb_data_o[16]
+ experiarSoC_peripherals/wb_data_o[17] experiarSoC_peripherals/wb_data_o[18] experiarSoC_peripherals/wb_data_o[19]
+ experiarSoC_peripherals/wb_data_o[1] experiarSoC_peripherals/wb_data_o[20] experiarSoC_peripherals/wb_data_o[21]
+ experiarSoC_peripherals/wb_data_o[22] experiarSoC_peripherals/wb_data_o[23] experiarSoC_peripherals/wb_data_o[24]
+ experiarSoC_peripherals/wb_data_o[25] experiarSoC_peripherals/wb_data_o[26] experiarSoC_peripherals/wb_data_o[27]
+ experiarSoC_peripherals/wb_data_o[28] experiarSoC_peripherals/wb_data_o[29] experiarSoC_peripherals/wb_data_o[2]
+ experiarSoC_peripherals/wb_data_o[30] experiarSoC_peripherals/wb_data_o[31] experiarSoC_peripherals/wb_data_o[3]
+ experiarSoC_peripherals/wb_data_o[4] experiarSoC_peripherals/wb_data_o[5] experiarSoC_peripherals/wb_data_o[6]
+ experiarSoC_peripherals/wb_data_o[7] experiarSoC_peripherals/wb_data_o[8] experiarSoC_peripherals/wb_data_o[9]
+ experiarSoC_peripherals/wb_error_o wb_rst_i experiarSoC_peripherals/wb_sel_i[0]
+ experiarSoC_peripherals/wb_sel_i[1] experiarSoC_peripherals/wb_sel_i[2] experiarSoC_peripherals/wb_sel_i[3]
+ experiarSoC_peripherals/wb_stall_o experiarSoC_peripherals/wb_stb_i experiarSoC_peripherals/wb_we_i
+ Peripherals
XexperiarSoC_wishboneInterconnect caravelHost/caravel_wb_ack_i caravelHost/caravel_wb_adr_o[0]
+ caravelHost/caravel_wb_adr_o[10] caravelHost/caravel_wb_adr_o[11] caravelHost/caravel_wb_adr_o[12]
+ caravelHost/caravel_wb_adr_o[13] caravelHost/caravel_wb_adr_o[14] caravelHost/caravel_wb_adr_o[15]
+ caravelHost/caravel_wb_adr_o[16] caravelHost/caravel_wb_adr_o[17] caravelHost/caravel_wb_adr_o[18]
+ caravelHost/caravel_wb_adr_o[19] caravelHost/caravel_wb_adr_o[1] caravelHost/caravel_wb_adr_o[20]
+ caravelHost/caravel_wb_adr_o[21] caravelHost/caravel_wb_adr_o[22] caravelHost/caravel_wb_adr_o[23]
+ caravelHost/caravel_wb_adr_o[24] caravelHost/caravel_wb_adr_o[25] caravelHost/caravel_wb_adr_o[26]
+ caravelHost/caravel_wb_adr_o[27] caravelHost/caravel_wb_adr_o[2] caravelHost/caravel_wb_adr_o[3]
+ caravelHost/caravel_wb_adr_o[4] caravelHost/caravel_wb_adr_o[5] caravelHost/caravel_wb_adr_o[6]
+ caravelHost/caravel_wb_adr_o[7] caravelHost/caravel_wb_adr_o[8] caravelHost/caravel_wb_adr_o[9]
+ caravelHost/caravel_wb_cyc_o caravelHost/caravel_wb_data_i[0] caravelHost/caravel_wb_data_i[10]
+ caravelHost/caravel_wb_data_i[11] caravelHost/caravel_wb_data_i[12] caravelHost/caravel_wb_data_i[13]
+ caravelHost/caravel_wb_data_i[14] caravelHost/caravel_wb_data_i[15] caravelHost/caravel_wb_data_i[16]
+ caravelHost/caravel_wb_data_i[17] caravelHost/caravel_wb_data_i[18] caravelHost/caravel_wb_data_i[19]
+ caravelHost/caravel_wb_data_i[1] caravelHost/caravel_wb_data_i[20] caravelHost/caravel_wb_data_i[21]
+ caravelHost/caravel_wb_data_i[22] caravelHost/caravel_wb_data_i[23] caravelHost/caravel_wb_data_i[24]
+ caravelHost/caravel_wb_data_i[25] caravelHost/caravel_wb_data_i[26] caravelHost/caravel_wb_data_i[27]
+ caravelHost/caravel_wb_data_i[28] caravelHost/caravel_wb_data_i[29] caravelHost/caravel_wb_data_i[2]
+ caravelHost/caravel_wb_data_i[30] caravelHost/caravel_wb_data_i[31] caravelHost/caravel_wb_data_i[3]
+ caravelHost/caravel_wb_data_i[4] caravelHost/caravel_wb_data_i[5] caravelHost/caravel_wb_data_i[6]
+ caravelHost/caravel_wb_data_i[7] caravelHost/caravel_wb_data_i[8] caravelHost/caravel_wb_data_i[9]
+ caravelHost/caravel_wb_data_o[0] caravelHost/caravel_wb_data_o[10] caravelHost/caravel_wb_data_o[11]
+ caravelHost/caravel_wb_data_o[12] caravelHost/caravel_wb_data_o[13] caravelHost/caravel_wb_data_o[14]
+ caravelHost/caravel_wb_data_o[15] caravelHost/caravel_wb_data_o[16] caravelHost/caravel_wb_data_o[17]
+ caravelHost/caravel_wb_data_o[18] caravelHost/caravel_wb_data_o[19] caravelHost/caravel_wb_data_o[1]
+ caravelHost/caravel_wb_data_o[20] caravelHost/caravel_wb_data_o[21] caravelHost/caravel_wb_data_o[22]
+ caravelHost/caravel_wb_data_o[23] caravelHost/caravel_wb_data_o[24] caravelHost/caravel_wb_data_o[25]
+ caravelHost/caravel_wb_data_o[26] caravelHost/caravel_wb_data_o[27] caravelHost/caravel_wb_data_o[28]
+ caravelHost/caravel_wb_data_o[29] caravelHost/caravel_wb_data_o[2] caravelHost/caravel_wb_data_o[30]
+ caravelHost/caravel_wb_data_o[31] caravelHost/caravel_wb_data_o[3] caravelHost/caravel_wb_data_o[4]
+ caravelHost/caravel_wb_data_o[5] caravelHost/caravel_wb_data_o[6] caravelHost/caravel_wb_data_o[7]
+ caravelHost/caravel_wb_data_o[8] caravelHost/caravel_wb_data_o[9] caravelHost/caravel_wb_error_i
+ caravelHost/caravel_wb_sel_o[0] caravelHost/caravel_wb_sel_o[1] caravelHost/caravel_wb_sel_o[2]
+ caravelHost/caravel_wb_sel_o[3] caravelHost/caravel_wb_stall_i caravelHost/caravel_wb_stb_o
+ caravelHost/caravel_wb_we_o experiarSoC_core0/core_wb_ack_i experiarSoC_core0/core_wb_adr_o[0]
+ experiarSoC_core0/core_wb_adr_o[10] experiarSoC_core0/core_wb_adr_o[11] experiarSoC_core0/core_wb_adr_o[12]
+ experiarSoC_core0/core_wb_adr_o[13] experiarSoC_core0/core_wb_adr_o[14] experiarSoC_core0/core_wb_adr_o[15]
+ experiarSoC_core0/core_wb_adr_o[16] experiarSoC_core0/core_wb_adr_o[17] experiarSoC_core0/core_wb_adr_o[18]
+ experiarSoC_core0/core_wb_adr_o[19] experiarSoC_core0/core_wb_adr_o[1] experiarSoC_core0/core_wb_adr_o[20]
+ experiarSoC_core0/core_wb_adr_o[21] experiarSoC_core0/core_wb_adr_o[22] experiarSoC_core0/core_wb_adr_o[23]
+ experiarSoC_core0/core_wb_adr_o[24] experiarSoC_core0/core_wb_adr_o[25] experiarSoC_core0/core_wb_adr_o[26]
+ experiarSoC_core0/core_wb_adr_o[27] experiarSoC_core0/core_wb_adr_o[2] experiarSoC_core0/core_wb_adr_o[3]
+ experiarSoC_core0/core_wb_adr_o[4] experiarSoC_core0/core_wb_adr_o[5] experiarSoC_core0/core_wb_adr_o[6]
+ experiarSoC_core0/core_wb_adr_o[7] experiarSoC_core0/core_wb_adr_o[8] experiarSoC_core0/core_wb_adr_o[9]
+ experiarSoC_core0/core_wb_cyc_o experiarSoC_core0/core_wb_data_i[0] experiarSoC_core0/core_wb_data_i[10]
+ experiarSoC_core0/core_wb_data_i[11] experiarSoC_core0/core_wb_data_i[12] experiarSoC_core0/core_wb_data_i[13]
+ experiarSoC_core0/core_wb_data_i[14] experiarSoC_core0/core_wb_data_i[15] experiarSoC_core0/core_wb_data_i[16]
+ experiarSoC_core0/core_wb_data_i[17] experiarSoC_core0/core_wb_data_i[18] experiarSoC_core0/core_wb_data_i[19]
+ experiarSoC_core0/core_wb_data_i[1] experiarSoC_core0/core_wb_data_i[20] experiarSoC_core0/core_wb_data_i[21]
+ experiarSoC_core0/core_wb_data_i[22] experiarSoC_core0/core_wb_data_i[23] experiarSoC_core0/core_wb_data_i[24]
+ experiarSoC_core0/core_wb_data_i[25] experiarSoC_core0/core_wb_data_i[26] experiarSoC_core0/core_wb_data_i[27]
+ experiarSoC_core0/core_wb_data_i[28] experiarSoC_core0/core_wb_data_i[29] experiarSoC_core0/core_wb_data_i[2]
+ experiarSoC_core0/core_wb_data_i[30] experiarSoC_core0/core_wb_data_i[31] experiarSoC_core0/core_wb_data_i[3]
+ experiarSoC_core0/core_wb_data_i[4] experiarSoC_core0/core_wb_data_i[5] experiarSoC_core0/core_wb_data_i[6]
+ experiarSoC_core0/core_wb_data_i[7] experiarSoC_core0/core_wb_data_i[8] experiarSoC_core0/core_wb_data_i[9]
+ experiarSoC_core0/core_wb_data_o[0] experiarSoC_core0/core_wb_data_o[10] experiarSoC_core0/core_wb_data_o[11]
+ experiarSoC_core0/core_wb_data_o[12] experiarSoC_core0/core_wb_data_o[13] experiarSoC_core0/core_wb_data_o[14]
+ experiarSoC_core0/core_wb_data_o[15] experiarSoC_core0/core_wb_data_o[16] experiarSoC_core0/core_wb_data_o[17]
+ experiarSoC_core0/core_wb_data_o[18] experiarSoC_core0/core_wb_data_o[19] experiarSoC_core0/core_wb_data_o[1]
+ experiarSoC_core0/core_wb_data_o[20] experiarSoC_core0/core_wb_data_o[21] experiarSoC_core0/core_wb_data_o[22]
+ experiarSoC_core0/core_wb_data_o[23] experiarSoC_core0/core_wb_data_o[24] experiarSoC_core0/core_wb_data_o[25]
+ experiarSoC_core0/core_wb_data_o[26] experiarSoC_core0/core_wb_data_o[27] experiarSoC_core0/core_wb_data_o[28]
+ experiarSoC_core0/core_wb_data_o[29] experiarSoC_core0/core_wb_data_o[2] experiarSoC_core0/core_wb_data_o[30]
+ experiarSoC_core0/core_wb_data_o[31] experiarSoC_core0/core_wb_data_o[3] experiarSoC_core0/core_wb_data_o[4]
+ experiarSoC_core0/core_wb_data_o[5] experiarSoC_core0/core_wb_data_o[6] experiarSoC_core0/core_wb_data_o[7]
+ experiarSoC_core0/core_wb_data_o[8] experiarSoC_core0/core_wb_data_o[9] experiarSoC_core0/core_wb_error_i
+ experiarSoC_core0/core_wb_sel_o[0] experiarSoC_core0/core_wb_sel_o[1] experiarSoC_core0/core_wb_sel_o[2]
+ experiarSoC_core0/core_wb_sel_o[3] experiarSoC_core0/core_wb_stall_i experiarSoC_core0/core_wb_stb_o
+ experiarSoC_core0/core_wb_we_o experiarSoC_core1/core_wb_ack_i experiarSoC_core1/core_wb_adr_o[0]
+ experiarSoC_core1/core_wb_adr_o[10] experiarSoC_core1/core_wb_adr_o[11] experiarSoC_core1/core_wb_adr_o[12]
+ experiarSoC_core1/core_wb_adr_o[13] experiarSoC_core1/core_wb_adr_o[14] experiarSoC_core1/core_wb_adr_o[15]
+ experiarSoC_core1/core_wb_adr_o[16] experiarSoC_core1/core_wb_adr_o[17] experiarSoC_core1/core_wb_adr_o[18]
+ experiarSoC_core1/core_wb_adr_o[19] experiarSoC_core1/core_wb_adr_o[1] experiarSoC_core1/core_wb_adr_o[20]
+ experiarSoC_core1/core_wb_adr_o[21] experiarSoC_core1/core_wb_adr_o[22] experiarSoC_core1/core_wb_adr_o[23]
+ experiarSoC_core1/core_wb_adr_o[24] experiarSoC_core1/core_wb_adr_o[25] experiarSoC_core1/core_wb_adr_o[26]
+ experiarSoC_core1/core_wb_adr_o[27] experiarSoC_core1/core_wb_adr_o[2] experiarSoC_core1/core_wb_adr_o[3]
+ experiarSoC_core1/core_wb_adr_o[4] experiarSoC_core1/core_wb_adr_o[5] experiarSoC_core1/core_wb_adr_o[6]
+ experiarSoC_core1/core_wb_adr_o[7] experiarSoC_core1/core_wb_adr_o[8] experiarSoC_core1/core_wb_adr_o[9]
+ experiarSoC_core1/core_wb_cyc_o experiarSoC_core1/core_wb_data_i[0] experiarSoC_core1/core_wb_data_i[10]
+ experiarSoC_core1/core_wb_data_i[11] experiarSoC_core1/core_wb_data_i[12] experiarSoC_core1/core_wb_data_i[13]
+ experiarSoC_core1/core_wb_data_i[14] experiarSoC_core1/core_wb_data_i[15] experiarSoC_core1/core_wb_data_i[16]
+ experiarSoC_core1/core_wb_data_i[17] experiarSoC_core1/core_wb_data_i[18] experiarSoC_core1/core_wb_data_i[19]
+ experiarSoC_core1/core_wb_data_i[1] experiarSoC_core1/core_wb_data_i[20] experiarSoC_core1/core_wb_data_i[21]
+ experiarSoC_core1/core_wb_data_i[22] experiarSoC_core1/core_wb_data_i[23] experiarSoC_core1/core_wb_data_i[24]
+ experiarSoC_core1/core_wb_data_i[25] experiarSoC_core1/core_wb_data_i[26] experiarSoC_core1/core_wb_data_i[27]
+ experiarSoC_core1/core_wb_data_i[28] experiarSoC_core1/core_wb_data_i[29] experiarSoC_core1/core_wb_data_i[2]
+ experiarSoC_core1/core_wb_data_i[30] experiarSoC_core1/core_wb_data_i[31] experiarSoC_core1/core_wb_data_i[3]
+ experiarSoC_core1/core_wb_data_i[4] experiarSoC_core1/core_wb_data_i[5] experiarSoC_core1/core_wb_data_i[6]
+ experiarSoC_core1/core_wb_data_i[7] experiarSoC_core1/core_wb_data_i[8] experiarSoC_core1/core_wb_data_i[9]
+ experiarSoC_core1/core_wb_data_o[0] experiarSoC_core1/core_wb_data_o[10] experiarSoC_core1/core_wb_data_o[11]
+ experiarSoC_core1/core_wb_data_o[12] experiarSoC_core1/core_wb_data_o[13] experiarSoC_core1/core_wb_data_o[14]
+ experiarSoC_core1/core_wb_data_o[15] experiarSoC_core1/core_wb_data_o[16] experiarSoC_core1/core_wb_data_o[17]
+ experiarSoC_core1/core_wb_data_o[18] experiarSoC_core1/core_wb_data_o[19] experiarSoC_core1/core_wb_data_o[1]
+ experiarSoC_core1/core_wb_data_o[20] experiarSoC_core1/core_wb_data_o[21] experiarSoC_core1/core_wb_data_o[22]
+ experiarSoC_core1/core_wb_data_o[23] experiarSoC_core1/core_wb_data_o[24] experiarSoC_core1/core_wb_data_o[25]
+ experiarSoC_core1/core_wb_data_o[26] experiarSoC_core1/core_wb_data_o[27] experiarSoC_core1/core_wb_data_o[28]
+ experiarSoC_core1/core_wb_data_o[29] experiarSoC_core1/core_wb_data_o[2] experiarSoC_core1/core_wb_data_o[30]
+ experiarSoC_core1/core_wb_data_o[31] experiarSoC_core1/core_wb_data_o[3] experiarSoC_core1/core_wb_data_o[4]
+ experiarSoC_core1/core_wb_data_o[5] experiarSoC_core1/core_wb_data_o[6] experiarSoC_core1/core_wb_data_o[7]
+ experiarSoC_core1/core_wb_data_o[8] experiarSoC_core1/core_wb_data_o[9] experiarSoC_core1/core_wb_error_i
+ experiarSoC_core1/core_wb_sel_o[0] experiarSoC_core1/core_wb_sel_o[1] experiarSoC_core1/core_wb_sel_o[2]
+ experiarSoC_core1/core_wb_sel_o[3] experiarSoC_core1/core_wb_stall_i experiarSoC_core1/core_wb_stb_o
+ experiarSoC_core1/core_wb_we_o la_data_out[2] la_data_out[3] la_data_out[4] la_data_out[5]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] experiarSoC_core0/localMemory_wb_ack_o experiarSoC_core0/localMemory_wb_adr_i[0]
+ experiarSoC_core0/localMemory_wb_adr_i[10] experiarSoC_core0/localMemory_wb_adr_i[11]
+ experiarSoC_core0/localMemory_wb_adr_i[12] experiarSoC_core0/localMemory_wb_adr_i[13]
+ experiarSoC_core0/localMemory_wb_adr_i[14] experiarSoC_core0/localMemory_wb_adr_i[15]
+ experiarSoC_core0/localMemory_wb_adr_i[16] experiarSoC_core0/localMemory_wb_adr_i[17]
+ experiarSoC_core0/localMemory_wb_adr_i[18] experiarSoC_core0/localMemory_wb_adr_i[19]
+ experiarSoC_core0/localMemory_wb_adr_i[1] experiarSoC_core0/localMemory_wb_adr_i[20]
+ experiarSoC_core0/localMemory_wb_adr_i[21] experiarSoC_core0/localMemory_wb_adr_i[22]
+ experiarSoC_core0/localMemory_wb_adr_i[23] experiarSoC_core0/localMemory_wb_adr_i[2]
+ experiarSoC_core0/localMemory_wb_adr_i[3] experiarSoC_core0/localMemory_wb_adr_i[4]
+ experiarSoC_core0/localMemory_wb_adr_i[5] experiarSoC_core0/localMemory_wb_adr_i[6]
+ experiarSoC_core0/localMemory_wb_adr_i[7] experiarSoC_core0/localMemory_wb_adr_i[8]
+ experiarSoC_core0/localMemory_wb_adr_i[9] experiarSoC_core0/localMemory_wb_cyc_i
+ experiarSoC_core0/localMemory_wb_data_i[0] experiarSoC_core0/localMemory_wb_data_i[10]
+ experiarSoC_core0/localMemory_wb_data_i[11] experiarSoC_core0/localMemory_wb_data_i[12]
+ experiarSoC_core0/localMemory_wb_data_i[13] experiarSoC_core0/localMemory_wb_data_i[14]
+ experiarSoC_core0/localMemory_wb_data_i[15] experiarSoC_core0/localMemory_wb_data_i[16]
+ experiarSoC_core0/localMemory_wb_data_i[17] experiarSoC_core0/localMemory_wb_data_i[18]
+ experiarSoC_core0/localMemory_wb_data_i[19] experiarSoC_core0/localMemory_wb_data_i[1]
+ experiarSoC_core0/localMemory_wb_data_i[20] experiarSoC_core0/localMemory_wb_data_i[21]
+ experiarSoC_core0/localMemory_wb_data_i[22] experiarSoC_core0/localMemory_wb_data_i[23]
+ experiarSoC_core0/localMemory_wb_data_i[24] experiarSoC_core0/localMemory_wb_data_i[25]
+ experiarSoC_core0/localMemory_wb_data_i[26] experiarSoC_core0/localMemory_wb_data_i[27]
+ experiarSoC_core0/localMemory_wb_data_i[28] experiarSoC_core0/localMemory_wb_data_i[29]
+ experiarSoC_core0/localMemory_wb_data_i[2] experiarSoC_core0/localMemory_wb_data_i[30]
+ experiarSoC_core0/localMemory_wb_data_i[31] experiarSoC_core0/localMemory_wb_data_i[3]
+ experiarSoC_core0/localMemory_wb_data_i[4] experiarSoC_core0/localMemory_wb_data_i[5]
+ experiarSoC_core0/localMemory_wb_data_i[6] experiarSoC_core0/localMemory_wb_data_i[7]
+ experiarSoC_core0/localMemory_wb_data_i[8] experiarSoC_core0/localMemory_wb_data_i[9]
+ experiarSoC_core0/localMemory_wb_data_o[0] experiarSoC_core0/localMemory_wb_data_o[10]
+ experiarSoC_core0/localMemory_wb_data_o[11] experiarSoC_core0/localMemory_wb_data_o[12]
+ experiarSoC_core0/localMemory_wb_data_o[13] experiarSoC_core0/localMemory_wb_data_o[14]
+ experiarSoC_core0/localMemory_wb_data_o[15] experiarSoC_core0/localMemory_wb_data_o[16]
+ experiarSoC_core0/localMemory_wb_data_o[17] experiarSoC_core0/localMemory_wb_data_o[18]
+ experiarSoC_core0/localMemory_wb_data_o[19] experiarSoC_core0/localMemory_wb_data_o[1]
+ experiarSoC_core0/localMemory_wb_data_o[20] experiarSoC_core0/localMemory_wb_data_o[21]
+ experiarSoC_core0/localMemory_wb_data_o[22] experiarSoC_core0/localMemory_wb_data_o[23]
+ experiarSoC_core0/localMemory_wb_data_o[24] experiarSoC_core0/localMemory_wb_data_o[25]
+ experiarSoC_core0/localMemory_wb_data_o[26] experiarSoC_core0/localMemory_wb_data_o[27]
+ experiarSoC_core0/localMemory_wb_data_o[28] experiarSoC_core0/localMemory_wb_data_o[29]
+ experiarSoC_core0/localMemory_wb_data_o[2] experiarSoC_core0/localMemory_wb_data_o[30]
+ experiarSoC_core0/localMemory_wb_data_o[31] experiarSoC_core0/localMemory_wb_data_o[3]
+ experiarSoC_core0/localMemory_wb_data_o[4] experiarSoC_core0/localMemory_wb_data_o[5]
+ experiarSoC_core0/localMemory_wb_data_o[6] experiarSoC_core0/localMemory_wb_data_o[7]
+ experiarSoC_core0/localMemory_wb_data_o[8] experiarSoC_core0/localMemory_wb_data_o[9]
+ experiarSoC_core0/localMemory_wb_error_o experiarSoC_core0/localMemory_wb_sel_i[0]
+ experiarSoC_core0/localMemory_wb_sel_i[1] experiarSoC_core0/localMemory_wb_sel_i[2]
+ experiarSoC_core0/localMemory_wb_sel_i[3] experiarSoC_core0/localMemory_wb_stall_o
+ experiarSoC_core0/localMemory_wb_stb_i experiarSoC_core0/localMemory_wb_we_i experiarSoC_core1/localMemory_wb_ack_o
+ experiarSoC_core1/localMemory_wb_adr_i[0] experiarSoC_core1/localMemory_wb_adr_i[10]
+ experiarSoC_core1/localMemory_wb_adr_i[11] experiarSoC_core1/localMemory_wb_adr_i[12]
+ experiarSoC_core1/localMemory_wb_adr_i[13] experiarSoC_core1/localMemory_wb_adr_i[14]
+ experiarSoC_core1/localMemory_wb_adr_i[15] experiarSoC_core1/localMemory_wb_adr_i[16]
+ experiarSoC_core1/localMemory_wb_adr_i[17] experiarSoC_core1/localMemory_wb_adr_i[18]
+ experiarSoC_core1/localMemory_wb_adr_i[19] experiarSoC_core1/localMemory_wb_adr_i[1]
+ experiarSoC_core1/localMemory_wb_adr_i[20] experiarSoC_core1/localMemory_wb_adr_i[21]
+ experiarSoC_core1/localMemory_wb_adr_i[22] experiarSoC_core1/localMemory_wb_adr_i[23]
+ experiarSoC_core1/localMemory_wb_adr_i[2] experiarSoC_core1/localMemory_wb_adr_i[3]
+ experiarSoC_core1/localMemory_wb_adr_i[4] experiarSoC_core1/localMemory_wb_adr_i[5]
+ experiarSoC_core1/localMemory_wb_adr_i[6] experiarSoC_core1/localMemory_wb_adr_i[7]
+ experiarSoC_core1/localMemory_wb_adr_i[8] experiarSoC_core1/localMemory_wb_adr_i[9]
+ experiarSoC_core1/localMemory_wb_cyc_i experiarSoC_core1/localMemory_wb_data_i[0]
+ experiarSoC_core1/localMemory_wb_data_i[10] experiarSoC_core1/localMemory_wb_data_i[11]
+ experiarSoC_core1/localMemory_wb_data_i[12] experiarSoC_core1/localMemory_wb_data_i[13]
+ experiarSoC_core1/localMemory_wb_data_i[14] experiarSoC_core1/localMemory_wb_data_i[15]
+ experiarSoC_core1/localMemory_wb_data_i[16] experiarSoC_core1/localMemory_wb_data_i[17]
+ experiarSoC_core1/localMemory_wb_data_i[18] experiarSoC_core1/localMemory_wb_data_i[19]
+ experiarSoC_core1/localMemory_wb_data_i[1] experiarSoC_core1/localMemory_wb_data_i[20]
+ experiarSoC_core1/localMemory_wb_data_i[21] experiarSoC_core1/localMemory_wb_data_i[22]
+ experiarSoC_core1/localMemory_wb_data_i[23] experiarSoC_core1/localMemory_wb_data_i[24]
+ experiarSoC_core1/localMemory_wb_data_i[25] experiarSoC_core1/localMemory_wb_data_i[26]
+ experiarSoC_core1/localMemory_wb_data_i[27] experiarSoC_core1/localMemory_wb_data_i[28]
+ experiarSoC_core1/localMemory_wb_data_i[29] experiarSoC_core1/localMemory_wb_data_i[2]
+ experiarSoC_core1/localMemory_wb_data_i[30] experiarSoC_core1/localMemory_wb_data_i[31]
+ experiarSoC_core1/localMemory_wb_data_i[3] experiarSoC_core1/localMemory_wb_data_i[4]
+ experiarSoC_core1/localMemory_wb_data_i[5] experiarSoC_core1/localMemory_wb_data_i[6]
+ experiarSoC_core1/localMemory_wb_data_i[7] experiarSoC_core1/localMemory_wb_data_i[8]
+ experiarSoC_core1/localMemory_wb_data_i[9] experiarSoC_core1/localMemory_wb_data_o[0]
+ experiarSoC_core1/localMemory_wb_data_o[10] experiarSoC_core1/localMemory_wb_data_o[11]
+ experiarSoC_core1/localMemory_wb_data_o[12] experiarSoC_core1/localMemory_wb_data_o[13]
+ experiarSoC_core1/localMemory_wb_data_o[14] experiarSoC_core1/localMemory_wb_data_o[15]
+ experiarSoC_core1/localMemory_wb_data_o[16] experiarSoC_core1/localMemory_wb_data_o[17]
+ experiarSoC_core1/localMemory_wb_data_o[18] experiarSoC_core1/localMemory_wb_data_o[19]
+ experiarSoC_core1/localMemory_wb_data_o[1] experiarSoC_core1/localMemory_wb_data_o[20]
+ experiarSoC_core1/localMemory_wb_data_o[21] experiarSoC_core1/localMemory_wb_data_o[22]
+ experiarSoC_core1/localMemory_wb_data_o[23] experiarSoC_core1/localMemory_wb_data_o[24]
+ experiarSoC_core1/localMemory_wb_data_o[25] experiarSoC_core1/localMemory_wb_data_o[26]
+ experiarSoC_core1/localMemory_wb_data_o[27] experiarSoC_core1/localMemory_wb_data_o[28]
+ experiarSoC_core1/localMemory_wb_data_o[29] experiarSoC_core1/localMemory_wb_data_o[2]
+ experiarSoC_core1/localMemory_wb_data_o[30] experiarSoC_core1/localMemory_wb_data_o[31]
+ experiarSoC_core1/localMemory_wb_data_o[3] experiarSoC_core1/localMemory_wb_data_o[4]
+ experiarSoC_core1/localMemory_wb_data_o[5] experiarSoC_core1/localMemory_wb_data_o[6]
+ experiarSoC_core1/localMemory_wb_data_o[7] experiarSoC_core1/localMemory_wb_data_o[8]
+ experiarSoC_core1/localMemory_wb_data_o[9] experiarSoC_core1/localMemory_wb_error_o
+ experiarSoC_core1/localMemory_wb_sel_i[0] experiarSoC_core1/localMemory_wb_sel_i[1]
+ experiarSoC_core1/localMemory_wb_sel_i[2] experiarSoC_core1/localMemory_wb_sel_i[3]
+ experiarSoC_core1/localMemory_wb_stall_o experiarSoC_core1/localMemory_wb_stb_i
+ experiarSoC_core1/localMemory_wb_we_i experiarSoC_video/wb_ack_o experiarSoC_video/wb_adr_i[0]
+ experiarSoC_video/wb_adr_i[10] experiarSoC_video/wb_adr_i[11] experiarSoC_video/wb_adr_i[12]
+ experiarSoC_video/wb_adr_i[13] experiarSoC_video/wb_adr_i[14] experiarSoC_video/wb_adr_i[15]
+ experiarSoC_video/wb_adr_i[16] experiarSoC_video/wb_adr_i[17] experiarSoC_video/wb_adr_i[18]
+ experiarSoC_video/wb_adr_i[19] experiarSoC_video/wb_adr_i[1] experiarSoC_video/wb_adr_i[20]
+ experiarSoC_video/wb_adr_i[21] experiarSoC_video/wb_adr_i[22] experiarSoC_video/wb_adr_i[23]
+ experiarSoC_video/wb_adr_i[2] experiarSoC_video/wb_adr_i[3] experiarSoC_video/wb_adr_i[4]
+ experiarSoC_video/wb_adr_i[5] experiarSoC_video/wb_adr_i[6] experiarSoC_video/wb_adr_i[7]
+ experiarSoC_video/wb_adr_i[8] experiarSoC_video/wb_adr_i[9] experiarSoC_video/wb_cyc_i
+ experiarSoC_video/wb_data_i[0] experiarSoC_video/wb_data_i[10] experiarSoC_video/wb_data_i[11]
+ experiarSoC_video/wb_data_i[12] experiarSoC_video/wb_data_i[13] experiarSoC_video/wb_data_i[14]
+ experiarSoC_video/wb_data_i[15] experiarSoC_video/wb_data_i[16] experiarSoC_video/wb_data_i[17]
+ experiarSoC_video/wb_data_i[18] experiarSoC_video/wb_data_i[19] experiarSoC_video/wb_data_i[1]
+ experiarSoC_video/wb_data_i[20] experiarSoC_video/wb_data_i[21] experiarSoC_video/wb_data_i[22]
+ experiarSoC_video/wb_data_i[23] experiarSoC_video/wb_data_i[24] experiarSoC_video/wb_data_i[25]
+ experiarSoC_video/wb_data_i[26] experiarSoC_video/wb_data_i[27] experiarSoC_video/wb_data_i[28]
+ experiarSoC_video/wb_data_i[29] experiarSoC_video/wb_data_i[2] experiarSoC_video/wb_data_i[30]
+ experiarSoC_video/wb_data_i[31] experiarSoC_video/wb_data_i[3] experiarSoC_video/wb_data_i[4]
+ experiarSoC_video/wb_data_i[5] experiarSoC_video/wb_data_i[6] experiarSoC_video/wb_data_i[7]
+ experiarSoC_video/wb_data_i[8] experiarSoC_video/wb_data_i[9] experiarSoC_video/wb_data_o[0]
+ experiarSoC_video/wb_data_o[10] experiarSoC_video/wb_data_o[11] experiarSoC_video/wb_data_o[12]
+ experiarSoC_video/wb_data_o[13] experiarSoC_video/wb_data_o[14] experiarSoC_video/wb_data_o[15]
+ experiarSoC_video/wb_data_o[16] experiarSoC_video/wb_data_o[17] experiarSoC_video/wb_data_o[18]
+ experiarSoC_video/wb_data_o[19] experiarSoC_video/wb_data_o[1] experiarSoC_video/wb_data_o[20]
+ experiarSoC_video/wb_data_o[21] experiarSoC_video/wb_data_o[22] experiarSoC_video/wb_data_o[23]
+ experiarSoC_video/wb_data_o[24] experiarSoC_video/wb_data_o[25] experiarSoC_video/wb_data_o[26]
+ experiarSoC_video/wb_data_o[27] experiarSoC_video/wb_data_o[28] experiarSoC_video/wb_data_o[29]
+ experiarSoC_video/wb_data_o[2] experiarSoC_video/wb_data_o[30] experiarSoC_video/wb_data_o[31]
+ experiarSoC_video/wb_data_o[3] experiarSoC_video/wb_data_o[4] experiarSoC_video/wb_data_o[5]
+ experiarSoC_video/wb_data_o[6] experiarSoC_video/wb_data_o[7] experiarSoC_video/wb_data_o[8]
+ experiarSoC_video/wb_data_o[9] experiarSoC_video/wb_error_o experiarSoC_video/wb_sel_i[0]
+ experiarSoC_video/wb_sel_i[1] experiarSoC_video/wb_sel_i[2] experiarSoC_video/wb_sel_i[3]
+ experiarSoC_video/wb_stall_o experiarSoC_video/wb_stb_i experiarSoC_video/wb_we_i
+ experiarSoC_peripherals/wb_ack_o experiarSoC_peripherals/wb_adr_i[0] experiarSoC_peripherals/wb_adr_i[10]
+ experiarSoC_peripherals/wb_adr_i[11] experiarSoC_peripherals/wb_adr_i[12] experiarSoC_peripherals/wb_adr_i[13]
+ experiarSoC_peripherals/wb_adr_i[14] experiarSoC_peripherals/wb_adr_i[15] experiarSoC_peripherals/wb_adr_i[16]
+ experiarSoC_peripherals/wb_adr_i[17] experiarSoC_peripherals/wb_adr_i[18] experiarSoC_peripherals/wb_adr_i[19]
+ experiarSoC_peripherals/wb_adr_i[1] experiarSoC_peripherals/wb_adr_i[20] experiarSoC_peripherals/wb_adr_i[21]
+ experiarSoC_peripherals/wb_adr_i[22] experiarSoC_peripherals/wb_adr_i[23] experiarSoC_peripherals/wb_adr_i[2]
+ experiarSoC_peripherals/wb_adr_i[3] experiarSoC_peripherals/wb_adr_i[4] experiarSoC_peripherals/wb_adr_i[5]
+ experiarSoC_peripherals/wb_adr_i[6] experiarSoC_peripherals/wb_adr_i[7] experiarSoC_peripherals/wb_adr_i[8]
+ experiarSoC_peripherals/wb_adr_i[9] experiarSoC_peripherals/wb_cyc_i experiarSoC_peripherals/wb_data_i[0]
+ experiarSoC_peripherals/wb_data_i[10] experiarSoC_peripherals/wb_data_i[11] experiarSoC_peripherals/wb_data_i[12]
+ experiarSoC_peripherals/wb_data_i[13] experiarSoC_peripherals/wb_data_i[14] experiarSoC_peripherals/wb_data_i[15]
+ experiarSoC_peripherals/wb_data_i[16] experiarSoC_peripherals/wb_data_i[17] experiarSoC_peripherals/wb_data_i[18]
+ experiarSoC_peripherals/wb_data_i[19] experiarSoC_peripherals/wb_data_i[1] experiarSoC_peripherals/wb_data_i[20]
+ experiarSoC_peripherals/wb_data_i[21] experiarSoC_peripherals/wb_data_i[22] experiarSoC_peripherals/wb_data_i[23]
+ experiarSoC_peripherals/wb_data_i[24] experiarSoC_peripherals/wb_data_i[25] experiarSoC_peripherals/wb_data_i[26]
+ experiarSoC_peripherals/wb_data_i[27] experiarSoC_peripherals/wb_data_i[28] experiarSoC_peripherals/wb_data_i[29]
+ experiarSoC_peripherals/wb_data_i[2] experiarSoC_peripherals/wb_data_i[30] experiarSoC_peripherals/wb_data_i[31]
+ experiarSoC_peripherals/wb_data_i[3] experiarSoC_peripherals/wb_data_i[4] experiarSoC_peripherals/wb_data_i[5]
+ experiarSoC_peripherals/wb_data_i[6] experiarSoC_peripherals/wb_data_i[7] experiarSoC_peripherals/wb_data_i[8]
+ experiarSoC_peripherals/wb_data_i[9] experiarSoC_peripherals/wb_data_o[0] experiarSoC_peripherals/wb_data_o[10]
+ experiarSoC_peripherals/wb_data_o[11] experiarSoC_peripherals/wb_data_o[12] experiarSoC_peripherals/wb_data_o[13]
+ experiarSoC_peripherals/wb_data_o[14] experiarSoC_peripherals/wb_data_o[15] experiarSoC_peripherals/wb_data_o[16]
+ experiarSoC_peripherals/wb_data_o[17] experiarSoC_peripherals/wb_data_o[18] experiarSoC_peripherals/wb_data_o[19]
+ experiarSoC_peripherals/wb_data_o[1] experiarSoC_peripherals/wb_data_o[20] experiarSoC_peripherals/wb_data_o[21]
+ experiarSoC_peripherals/wb_data_o[22] experiarSoC_peripherals/wb_data_o[23] experiarSoC_peripherals/wb_data_o[24]
+ experiarSoC_peripherals/wb_data_o[25] experiarSoC_peripherals/wb_data_o[26] experiarSoC_peripherals/wb_data_o[27]
+ experiarSoC_peripherals/wb_data_o[28] experiarSoC_peripherals/wb_data_o[29] experiarSoC_peripherals/wb_data_o[2]
+ experiarSoC_peripherals/wb_data_o[30] experiarSoC_peripherals/wb_data_o[31] experiarSoC_peripherals/wb_data_o[3]
+ experiarSoC_peripherals/wb_data_o[4] experiarSoC_peripherals/wb_data_o[5] experiarSoC_peripherals/wb_data_o[6]
+ experiarSoC_peripherals/wb_data_o[7] experiarSoC_peripherals/wb_data_o[8] experiarSoC_peripherals/wb_data_o[9]
+ experiarSoC_peripherals/wb_error_o experiarSoC_peripherals/wb_sel_i[0] experiarSoC_peripherals/wb_sel_i[1]
+ experiarSoC_peripherals/wb_sel_i[2] experiarSoC_peripherals/wb_sel_i[3] experiarSoC_peripherals/wb_stall_o
+ experiarSoC_peripherals/wb_stb_i experiarSoC_peripherals/wb_we_i experiarSoC_flash/wb_ack_o
+ experiarSoC_flash/wb_adr_i[0] experiarSoC_flash/wb_adr_i[10] experiarSoC_flash/wb_adr_i[11]
+ experiarSoC_flash/wb_adr_i[12] experiarSoC_flash/wb_adr_i[13] experiarSoC_flash/wb_adr_i[14]
+ experiarSoC_flash/wb_adr_i[15] experiarSoC_flash/wb_adr_i[16] experiarSoC_flash/wb_adr_i[17]
+ experiarSoC_flash/wb_adr_i[18] experiarSoC_flash/wb_adr_i[19] experiarSoC_flash/wb_adr_i[1]
+ experiarSoC_flash/wb_adr_i[20] experiarSoC_flash/wb_adr_i[21] experiarSoC_flash/wb_adr_i[22]
+ experiarSoC_flash/wb_adr_i[23] experiarSoC_flash/wb_adr_i[2] experiarSoC_flash/wb_adr_i[3]
+ experiarSoC_flash/wb_adr_i[4] experiarSoC_flash/wb_adr_i[5] experiarSoC_flash/wb_adr_i[6]
+ experiarSoC_flash/wb_adr_i[7] experiarSoC_flash/wb_adr_i[8] experiarSoC_flash/wb_adr_i[9]
+ experiarSoC_flash/wb_cyc_i experiarSoC_flash/wb_data_i[0] experiarSoC_flash/wb_data_i[10]
+ experiarSoC_flash/wb_data_i[11] experiarSoC_flash/wb_data_i[12] experiarSoC_flash/wb_data_i[13]
+ experiarSoC_flash/wb_data_i[14] experiarSoC_flash/wb_data_i[15] experiarSoC_flash/wb_data_i[16]
+ experiarSoC_flash/wb_data_i[17] experiarSoC_flash/wb_data_i[18] experiarSoC_flash/wb_data_i[19]
+ experiarSoC_flash/wb_data_i[1] experiarSoC_flash/wb_data_i[20] experiarSoC_flash/wb_data_i[21]
+ experiarSoC_flash/wb_data_i[22] experiarSoC_flash/wb_data_i[23] experiarSoC_flash/wb_data_i[24]
+ experiarSoC_flash/wb_data_i[25] experiarSoC_flash/wb_data_i[26] experiarSoC_flash/wb_data_i[27]
+ experiarSoC_flash/wb_data_i[28] experiarSoC_flash/wb_data_i[29] experiarSoC_flash/wb_data_i[2]
+ experiarSoC_flash/wb_data_i[30] experiarSoC_flash/wb_data_i[31] experiarSoC_flash/wb_data_i[3]
+ experiarSoC_flash/wb_data_i[4] experiarSoC_flash/wb_data_i[5] experiarSoC_flash/wb_data_i[6]
+ experiarSoC_flash/wb_data_i[7] experiarSoC_flash/wb_data_i[8] experiarSoC_flash/wb_data_i[9]
+ experiarSoC_flash/wb_data_o[0] experiarSoC_flash/wb_data_o[10] experiarSoC_flash/wb_data_o[11]
+ experiarSoC_flash/wb_data_o[12] experiarSoC_flash/wb_data_o[13] experiarSoC_flash/wb_data_o[14]
+ experiarSoC_flash/wb_data_o[15] experiarSoC_flash/wb_data_o[16] experiarSoC_flash/wb_data_o[17]
+ experiarSoC_flash/wb_data_o[18] experiarSoC_flash/wb_data_o[19] experiarSoC_flash/wb_data_o[1]
+ experiarSoC_flash/wb_data_o[20] experiarSoC_flash/wb_data_o[21] experiarSoC_flash/wb_data_o[22]
+ experiarSoC_flash/wb_data_o[23] experiarSoC_flash/wb_data_o[24] experiarSoC_flash/wb_data_o[25]
+ experiarSoC_flash/wb_data_o[26] experiarSoC_flash/wb_data_o[27] experiarSoC_flash/wb_data_o[28]
+ experiarSoC_flash/wb_data_o[29] experiarSoC_flash/wb_data_o[2] experiarSoC_flash/wb_data_o[30]
+ experiarSoC_flash/wb_data_o[31] experiarSoC_flash/wb_data_o[3] experiarSoC_flash/wb_data_o[4]
+ experiarSoC_flash/wb_data_o[5] experiarSoC_flash/wb_data_o[6] experiarSoC_flash/wb_data_o[7]
+ experiarSoC_flash/wb_data_o[8] experiarSoC_flash/wb_data_o[9] experiarSoC_flash/wb_error_o
+ experiarSoC_flash/wb_sel_i[0] experiarSoC_flash/wb_sel_i[1] experiarSoC_flash/wb_sel_i[2]
+ experiarSoC_flash/wb_sel_i[3] experiarSoC_flash/wb_stall_o experiarSoC_flash/wb_stb_i
+ experiarSoC_flash/wb_we_i vccd1 vssd1 wb_clk_i wb_rst_i WishboneInterconnect
XcaravelHost caravelHost/caravel_irq[0] caravelHost/caravel_irq[1] caravelHost/caravel_irq[2]
+ caravelHost/caravel_irq[3] caravelHost/caravel_uart_rx caravelHost/caravel_uart_tx
+ caravelHost/caravel_wb_ack_i caravelHost/caravel_wb_adr_o[0] caravelHost/caravel_wb_adr_o[10]
+ caravelHost/caravel_wb_adr_o[11] caravelHost/caravel_wb_adr_o[12] caravelHost/caravel_wb_adr_o[13]
+ caravelHost/caravel_wb_adr_o[14] caravelHost/caravel_wb_adr_o[15] caravelHost/caravel_wb_adr_o[16]
+ caravelHost/caravel_wb_adr_o[17] caravelHost/caravel_wb_adr_o[18] caravelHost/caravel_wb_adr_o[19]
+ caravelHost/caravel_wb_adr_o[1] caravelHost/caravel_wb_adr_o[20] caravelHost/caravel_wb_adr_o[21]
+ caravelHost/caravel_wb_adr_o[22] caravelHost/caravel_wb_adr_o[23] caravelHost/caravel_wb_adr_o[24]
+ caravelHost/caravel_wb_adr_o[25] caravelHost/caravel_wb_adr_o[26] caravelHost/caravel_wb_adr_o[27]
+ caravelHost/caravel_wb_adr_o[2] caravelHost/caravel_wb_adr_o[3] caravelHost/caravel_wb_adr_o[4]
+ caravelHost/caravel_wb_adr_o[5] caravelHost/caravel_wb_adr_o[6] caravelHost/caravel_wb_adr_o[7]
+ caravelHost/caravel_wb_adr_o[8] caravelHost/caravel_wb_adr_o[9] caravelHost/caravel_wb_cyc_o
+ caravelHost/caravel_wb_data_i[0] caravelHost/caravel_wb_data_i[10] caravelHost/caravel_wb_data_i[11]
+ caravelHost/caravel_wb_data_i[12] caravelHost/caravel_wb_data_i[13] caravelHost/caravel_wb_data_i[14]
+ caravelHost/caravel_wb_data_i[15] caravelHost/caravel_wb_data_i[16] caravelHost/caravel_wb_data_i[17]
+ caravelHost/caravel_wb_data_i[18] caravelHost/caravel_wb_data_i[19] caravelHost/caravel_wb_data_i[1]
+ caravelHost/caravel_wb_data_i[20] caravelHost/caravel_wb_data_i[21] caravelHost/caravel_wb_data_i[22]
+ caravelHost/caravel_wb_data_i[23] caravelHost/caravel_wb_data_i[24] caravelHost/caravel_wb_data_i[25]
+ caravelHost/caravel_wb_data_i[26] caravelHost/caravel_wb_data_i[27] caravelHost/caravel_wb_data_i[28]
+ caravelHost/caravel_wb_data_i[29] caravelHost/caravel_wb_data_i[2] caravelHost/caravel_wb_data_i[30]
+ caravelHost/caravel_wb_data_i[31] caravelHost/caravel_wb_data_i[3] caravelHost/caravel_wb_data_i[4]
+ caravelHost/caravel_wb_data_i[5] caravelHost/caravel_wb_data_i[6] caravelHost/caravel_wb_data_i[7]
+ caravelHost/caravel_wb_data_i[8] caravelHost/caravel_wb_data_i[9] caravelHost/caravel_wb_data_o[0]
+ caravelHost/caravel_wb_data_o[10] caravelHost/caravel_wb_data_o[11] caravelHost/caravel_wb_data_o[12]
+ caravelHost/caravel_wb_data_o[13] caravelHost/caravel_wb_data_o[14] caravelHost/caravel_wb_data_o[15]
+ caravelHost/caravel_wb_data_o[16] caravelHost/caravel_wb_data_o[17] caravelHost/caravel_wb_data_o[18]
+ caravelHost/caravel_wb_data_o[19] caravelHost/caravel_wb_data_o[1] caravelHost/caravel_wb_data_o[20]
+ caravelHost/caravel_wb_data_o[21] caravelHost/caravel_wb_data_o[22] caravelHost/caravel_wb_data_o[23]
+ caravelHost/caravel_wb_data_o[24] caravelHost/caravel_wb_data_o[25] caravelHost/caravel_wb_data_o[26]
+ caravelHost/caravel_wb_data_o[27] caravelHost/caravel_wb_data_o[28] caravelHost/caravel_wb_data_o[29]
+ caravelHost/caravel_wb_data_o[2] caravelHost/caravel_wb_data_o[30] caravelHost/caravel_wb_data_o[31]
+ caravelHost/caravel_wb_data_o[3] caravelHost/caravel_wb_data_o[4] caravelHost/caravel_wb_data_o[5]
+ caravelHost/caravel_wb_data_o[6] caravelHost/caravel_wb_data_o[7] caravelHost/caravel_wb_data_o[8]
+ caravelHost/caravel_wb_data_o[9] caravelHost/caravel_wb_error_i caravelHost/caravel_wb_sel_o[0]
+ caravelHost/caravel_wb_sel_o[1] caravelHost/caravel_wb_sel_o[2] caravelHost/caravel_wb_sel_o[3]
+ caravelHost/caravel_wb_stall_i caravelHost/caravel_wb_stb_o caravelHost/caravel_wb_we_o
+ caravelHost/core0Index[0] caravelHost/core0Index[1] caravelHost/core0Index[2] caravelHost/core0Index[3]
+ caravelHost/core0Index[4] caravelHost/core0Index[5] caravelHost/core0Index[6] caravelHost/core0Index[7]
+ caravelHost/core1Index[0] caravelHost/core1Index[1] caravelHost/core1Index[2] caravelHost/core1Index[3]
+ caravelHost/core1Index[4] caravelHost/core1Index[5] caravelHost/core1Index[6] caravelHost/core1Index[7]
+ caravelHost/manufacturerID[0] caravelHost/manufacturerID[10] caravelHost/manufacturerID[1]
+ caravelHost/manufacturerID[2] caravelHost/manufacturerID[3] caravelHost/manufacturerID[4]
+ caravelHost/manufacturerID[5] caravelHost/manufacturerID[6] caravelHost/manufacturerID[7]
+ caravelHost/manufacturerID[8] caravelHost/manufacturerID[9] caravelHost/partID[0]
+ caravelHost/partID[10] caravelHost/partID[11] caravelHost/partID[12] caravelHost/partID[13]
+ caravelHost/partID[14] caravelHost/partID[15] caravelHost/partID[1] caravelHost/partID[2]
+ caravelHost/partID[3] caravelHost/partID[4] caravelHost/partID[5] caravelHost/partID[6]
+ caravelHost/partID[7] caravelHost/partID[8] caravelHost/partID[9] vccd1 caravelHost/versionID[0]
+ caravelHost/versionID[1] caravelHost/versionID[2] caravelHost/versionID[3] vssd1
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i CaravelHost
XexperiarSoC_core1SRAM0 experiarSoC_core1/din0[0] experiarSoC_core1/din0[1] experiarSoC_core1/din0[2]
+ experiarSoC_core1/din0[3] experiarSoC_core1/din0[4] experiarSoC_core1/din0[5] experiarSoC_core1/din0[6]
+ experiarSoC_core1/din0[7] experiarSoC_core1/din0[8] experiarSoC_core1/din0[9] experiarSoC_core1/din0[10]
+ experiarSoC_core1/din0[11] experiarSoC_core1/din0[12] experiarSoC_core1/din0[13]
+ experiarSoC_core1/din0[14] experiarSoC_core1/din0[15] experiarSoC_core1/din0[16]
+ experiarSoC_core1/din0[17] experiarSoC_core1/din0[18] experiarSoC_core1/din0[19]
+ experiarSoC_core1/din0[20] experiarSoC_core1/din0[21] experiarSoC_core1/din0[22]
+ experiarSoC_core1/din0[23] experiarSoC_core1/din0[24] experiarSoC_core1/din0[25]
+ experiarSoC_core1/din0[26] experiarSoC_core1/din0[27] experiarSoC_core1/din0[28]
+ experiarSoC_core1/din0[29] experiarSoC_core1/din0[30] experiarSoC_core1/din0[31]
+ experiarSoC_core1/addr0[0] experiarSoC_core1/addr0[1] experiarSoC_core1/addr0[2]
+ experiarSoC_core1/addr0[3] experiarSoC_core1/addr0[4] experiarSoC_core1/addr0[5]
+ experiarSoC_core1/addr0[6] experiarSoC_core1/addr0[7] experiarSoC_core1/addr0[8]
+ experiarSoC_core1/addr1[0] experiarSoC_core1/addr1[1] experiarSoC_core1/addr1[2]
+ experiarSoC_core1/addr1[3] experiarSoC_core1/addr1[4] experiarSoC_core1/addr1[5]
+ experiarSoC_core1/addr1[6] experiarSoC_core1/addr1[7] experiarSoC_core1/addr1[8]
+ experiarSoC_core1/csb0[0] experiarSoC_core1/csb1[0] experiarSoC_core1/web0 experiarSoC_core1/clk0
+ experiarSoC_core1/clk1 experiarSoC_core1/wmask0[0] experiarSoC_core1/wmask0[1] experiarSoC_core1/wmask0[2]
+ experiarSoC_core1/wmask0[3] experiarSoC_core1/dout0[0] experiarSoC_core1/dout0[1]
+ experiarSoC_core1/dout0[2] experiarSoC_core1/dout0[3] experiarSoC_core1/dout0[4]
+ experiarSoC_core1/dout0[5] experiarSoC_core1/dout0[6] experiarSoC_core1/dout0[7]
+ experiarSoC_core1/dout0[8] experiarSoC_core1/dout0[9] experiarSoC_core1/dout0[10]
+ experiarSoC_core1/dout0[11] experiarSoC_core1/dout0[12] experiarSoC_core1/dout0[13]
+ experiarSoC_core1/dout0[14] experiarSoC_core1/dout0[15] experiarSoC_core1/dout0[16]
+ experiarSoC_core1/dout0[17] experiarSoC_core1/dout0[18] experiarSoC_core1/dout0[19]
+ experiarSoC_core1/dout0[20] experiarSoC_core1/dout0[21] experiarSoC_core1/dout0[22]
+ experiarSoC_core1/dout0[23] experiarSoC_core1/dout0[24] experiarSoC_core1/dout0[25]
+ experiarSoC_core1/dout0[26] experiarSoC_core1/dout0[27] experiarSoC_core1/dout0[28]
+ experiarSoC_core1/dout0[29] experiarSoC_core1/dout0[30] experiarSoC_core1/dout0[31]
+ experiarSoC_core1/dout1[0] experiarSoC_core1/dout1[1] experiarSoC_core1/dout1[2]
+ experiarSoC_core1/dout1[3] experiarSoC_core1/dout1[4] experiarSoC_core1/dout1[5]
+ experiarSoC_core1/dout1[6] experiarSoC_core1/dout1[7] experiarSoC_core1/dout1[8]
+ experiarSoC_core1/dout1[9] experiarSoC_core1/dout1[10] experiarSoC_core1/dout1[11]
+ experiarSoC_core1/dout1[12] experiarSoC_core1/dout1[13] experiarSoC_core1/dout1[14]
+ experiarSoC_core1/dout1[15] experiarSoC_core1/dout1[16] experiarSoC_core1/dout1[17]
+ experiarSoC_core1/dout1[18] experiarSoC_core1/dout1[19] experiarSoC_core1/dout1[20]
+ experiarSoC_core1/dout1[21] experiarSoC_core1/dout1[22] experiarSoC_core1/dout1[23]
+ experiarSoC_core1/dout1[24] experiarSoC_core1/dout1[25] experiarSoC_core1/dout1[26]
+ experiarSoC_core1/dout1[27] experiarSoC_core1/dout1[28] experiarSoC_core1/dout1[29]
+ experiarSoC_core1/dout1[30] experiarSoC_core1/dout1[31] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_core1SRAM1 experiarSoC_core1/din0[0] experiarSoC_core1/din0[1] experiarSoC_core1/din0[2]
+ experiarSoC_core1/din0[3] experiarSoC_core1/din0[4] experiarSoC_core1/din0[5] experiarSoC_core1/din0[6]
+ experiarSoC_core1/din0[7] experiarSoC_core1/din0[8] experiarSoC_core1/din0[9] experiarSoC_core1/din0[10]
+ experiarSoC_core1/din0[11] experiarSoC_core1/din0[12] experiarSoC_core1/din0[13]
+ experiarSoC_core1/din0[14] experiarSoC_core1/din0[15] experiarSoC_core1/din0[16]
+ experiarSoC_core1/din0[17] experiarSoC_core1/din0[18] experiarSoC_core1/din0[19]
+ experiarSoC_core1/din0[20] experiarSoC_core1/din0[21] experiarSoC_core1/din0[22]
+ experiarSoC_core1/din0[23] experiarSoC_core1/din0[24] experiarSoC_core1/din0[25]
+ experiarSoC_core1/din0[26] experiarSoC_core1/din0[27] experiarSoC_core1/din0[28]
+ experiarSoC_core1/din0[29] experiarSoC_core1/din0[30] experiarSoC_core1/din0[31]
+ experiarSoC_core1/addr0[0] experiarSoC_core1/addr0[1] experiarSoC_core1/addr0[2]
+ experiarSoC_core1/addr0[3] experiarSoC_core1/addr0[4] experiarSoC_core1/addr0[5]
+ experiarSoC_core1/addr0[6] experiarSoC_core1/addr0[7] experiarSoC_core1/addr0[8]
+ experiarSoC_core1/addr1[0] experiarSoC_core1/addr1[1] experiarSoC_core1/addr1[2]
+ experiarSoC_core1/addr1[3] experiarSoC_core1/addr1[4] experiarSoC_core1/addr1[5]
+ experiarSoC_core1/addr1[6] experiarSoC_core1/addr1[7] experiarSoC_core1/addr1[8]
+ experiarSoC_core1/csb0[1] experiarSoC_core1/csb1[1] experiarSoC_core1/web0 experiarSoC_core1/clk0
+ experiarSoC_core1/clk1 experiarSoC_core1/wmask0[0] experiarSoC_core1/wmask0[1] experiarSoC_core1/wmask0[2]
+ experiarSoC_core1/wmask0[3] experiarSoC_core1/dout0[32] experiarSoC_core1/dout0[33]
+ experiarSoC_core1/dout0[34] experiarSoC_core1/dout0[35] experiarSoC_core1/dout0[36]
+ experiarSoC_core1/dout0[37] experiarSoC_core1/dout0[38] experiarSoC_core1/dout0[39]
+ experiarSoC_core1/dout0[40] experiarSoC_core1/dout0[41] experiarSoC_core1/dout0[42]
+ experiarSoC_core1/dout0[43] experiarSoC_core1/dout0[44] experiarSoC_core1/dout0[45]
+ experiarSoC_core1/dout0[46] experiarSoC_core1/dout0[47] experiarSoC_core1/dout0[48]
+ experiarSoC_core1/dout0[49] experiarSoC_core1/dout0[50] experiarSoC_core1/dout0[51]
+ experiarSoC_core1/dout0[52] experiarSoC_core1/dout0[53] experiarSoC_core1/dout0[54]
+ experiarSoC_core1/dout0[55] experiarSoC_core1/dout0[56] experiarSoC_core1/dout0[57]
+ experiarSoC_core1/dout0[58] experiarSoC_core1/dout0[59] experiarSoC_core1/dout0[60]
+ experiarSoC_core1/dout0[61] experiarSoC_core1/dout0[62] experiarSoC_core1/dout0[63]
+ experiarSoC_core1/dout1[32] experiarSoC_core1/dout1[33] experiarSoC_core1/dout1[34]
+ experiarSoC_core1/dout1[35] experiarSoC_core1/dout1[36] experiarSoC_core1/dout1[37]
+ experiarSoC_core1/dout1[38] experiarSoC_core1/dout1[39] experiarSoC_core1/dout1[40]
+ experiarSoC_core1/dout1[41] experiarSoC_core1/dout1[42] experiarSoC_core1/dout1[43]
+ experiarSoC_core1/dout1[44] experiarSoC_core1/dout1[45] experiarSoC_core1/dout1[46]
+ experiarSoC_core1/dout1[47] experiarSoC_core1/dout1[48] experiarSoC_core1/dout1[49]
+ experiarSoC_core1/dout1[50] experiarSoC_core1/dout1[51] experiarSoC_core1/dout1[52]
+ experiarSoC_core1/dout1[53] experiarSoC_core1/dout1[54] experiarSoC_core1/dout1[55]
+ experiarSoC_core1/dout1[56] experiarSoC_core1/dout1[57] experiarSoC_core1/dout1[58]
+ experiarSoC_core1/dout1[59] experiarSoC_core1/dout1[60] experiarSoC_core1/dout1[61]
+ experiarSoC_core1/dout1[62] experiarSoC_core1/dout1[63] vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
XexperiarSoC_video experiarSoC_videoSRAM1/addr0[0] experiarSoC_videoSRAM1/addr0[1]
+ experiarSoC_videoSRAM1/addr0[2] experiarSoC_videoSRAM1/addr0[3] experiarSoC_videoSRAM1/addr0[4]
+ experiarSoC_videoSRAM1/addr0[5] experiarSoC_videoSRAM1/addr0[6] experiarSoC_videoSRAM1/addr0[7]
+ experiarSoC_videoSRAM1/addr0[8] experiarSoC_videoSRAM1/addr1[0] experiarSoC_videoSRAM1/addr1[1]
+ experiarSoC_videoSRAM1/addr1[2] experiarSoC_videoSRAM1/addr1[3] experiarSoC_videoSRAM1/addr1[4]
+ experiarSoC_videoSRAM1/addr1[5] experiarSoC_videoSRAM1/addr1[6] experiarSoC_videoSRAM1/addr1[7]
+ experiarSoC_videoSRAM1/addr1[8] experiarSoC_videoSRAM1/clk0 experiarSoC_videoSRAM1/clk1
+ experiarSoC_videoSRAM0/csb0 experiarSoC_videoSRAM1/csb0 experiarSoC_videoSRAM0/csb1
+ experiarSoC_videoSRAM1/csb1 experiarSoC_videoSRAM1/din0[0] experiarSoC_videoSRAM1/din0[10]
+ experiarSoC_videoSRAM1/din0[11] experiarSoC_videoSRAM1/din0[12] experiarSoC_videoSRAM1/din0[13]
+ experiarSoC_videoSRAM1/din0[14] experiarSoC_videoSRAM1/din0[15] experiarSoC_videoSRAM1/din0[16]
+ experiarSoC_videoSRAM1/din0[17] experiarSoC_videoSRAM1/din0[18] experiarSoC_videoSRAM1/din0[19]
+ experiarSoC_videoSRAM1/din0[1] experiarSoC_videoSRAM1/din0[20] experiarSoC_videoSRAM1/din0[21]
+ experiarSoC_videoSRAM1/din0[22] experiarSoC_videoSRAM1/din0[23] experiarSoC_videoSRAM1/din0[24]
+ experiarSoC_videoSRAM1/din0[25] experiarSoC_videoSRAM1/din0[26] experiarSoC_videoSRAM1/din0[27]
+ experiarSoC_videoSRAM1/din0[28] experiarSoC_videoSRAM1/din0[29] experiarSoC_videoSRAM1/din0[2]
+ experiarSoC_videoSRAM1/din0[30] experiarSoC_videoSRAM1/din0[31] experiarSoC_videoSRAM1/din0[3]
+ experiarSoC_videoSRAM1/din0[4] experiarSoC_videoSRAM1/din0[5] experiarSoC_videoSRAM1/din0[6]
+ experiarSoC_videoSRAM1/din0[7] experiarSoC_videoSRAM1/din0[8] experiarSoC_videoSRAM1/din0[9]
+ experiarSoC_videoSRAM0/dout0[0] experiarSoC_videoSRAM0/dout0[10] experiarSoC_videoSRAM0/dout0[11]
+ experiarSoC_videoSRAM0/dout0[12] experiarSoC_videoSRAM0/dout0[13] experiarSoC_videoSRAM0/dout0[14]
+ experiarSoC_videoSRAM0/dout0[15] experiarSoC_videoSRAM0/dout0[16] experiarSoC_videoSRAM0/dout0[17]
+ experiarSoC_videoSRAM0/dout0[18] experiarSoC_videoSRAM0/dout0[19] experiarSoC_videoSRAM0/dout0[1]
+ experiarSoC_videoSRAM0/dout0[20] experiarSoC_videoSRAM0/dout0[21] experiarSoC_videoSRAM0/dout0[22]
+ experiarSoC_videoSRAM0/dout0[23] experiarSoC_videoSRAM0/dout0[24] experiarSoC_videoSRAM0/dout0[25]
+ experiarSoC_videoSRAM0/dout0[26] experiarSoC_videoSRAM0/dout0[27] experiarSoC_videoSRAM0/dout0[28]
+ experiarSoC_videoSRAM0/dout0[29] experiarSoC_videoSRAM0/dout0[2] experiarSoC_videoSRAM0/dout0[30]
+ experiarSoC_videoSRAM0/dout0[31] experiarSoC_videoSRAM1/dout0[0] experiarSoC_videoSRAM1/dout0[1]
+ experiarSoC_videoSRAM1/dout0[2] experiarSoC_videoSRAM1/dout0[3] experiarSoC_videoSRAM1/dout0[4]
+ experiarSoC_videoSRAM1/dout0[5] experiarSoC_videoSRAM1/dout0[6] experiarSoC_videoSRAM1/dout0[7]
+ experiarSoC_videoSRAM0/dout0[3] experiarSoC_videoSRAM1/dout0[8] experiarSoC_videoSRAM1/dout0[9]
+ experiarSoC_videoSRAM1/dout0[10] experiarSoC_videoSRAM1/dout0[11] experiarSoC_videoSRAM1/dout0[12]
+ experiarSoC_videoSRAM1/dout0[13] experiarSoC_videoSRAM1/dout0[14] experiarSoC_videoSRAM1/dout0[15]
+ experiarSoC_videoSRAM1/dout0[16] experiarSoC_videoSRAM1/dout0[17] experiarSoC_videoSRAM0/dout0[4]
+ experiarSoC_videoSRAM1/dout0[18] experiarSoC_videoSRAM1/dout0[19] experiarSoC_videoSRAM1/dout0[20]
+ experiarSoC_videoSRAM1/dout0[21] experiarSoC_videoSRAM1/dout0[22] experiarSoC_videoSRAM1/dout0[23]
+ experiarSoC_videoSRAM1/dout0[24] experiarSoC_videoSRAM1/dout0[25] experiarSoC_videoSRAM1/dout0[26]
+ experiarSoC_videoSRAM1/dout0[27] experiarSoC_videoSRAM0/dout0[5] experiarSoC_videoSRAM1/dout0[28]
+ experiarSoC_videoSRAM1/dout0[29] experiarSoC_videoSRAM1/dout0[30] experiarSoC_videoSRAM1/dout0[31]
+ experiarSoC_videoSRAM0/dout0[6] experiarSoC_videoSRAM0/dout0[7] experiarSoC_videoSRAM0/dout0[8]
+ experiarSoC_videoSRAM0/dout0[9] experiarSoC_videoSRAM0/dout1[0] experiarSoC_videoSRAM0/dout1[10]
+ experiarSoC_videoSRAM0/dout1[11] experiarSoC_videoSRAM0/dout1[12] experiarSoC_videoSRAM0/dout1[13]
+ experiarSoC_videoSRAM0/dout1[14] experiarSoC_videoSRAM0/dout1[15] experiarSoC_videoSRAM0/dout1[16]
+ experiarSoC_videoSRAM0/dout1[17] experiarSoC_videoSRAM0/dout1[18] experiarSoC_videoSRAM0/dout1[19]
+ experiarSoC_videoSRAM0/dout1[1] experiarSoC_videoSRAM0/dout1[20] experiarSoC_videoSRAM0/dout1[21]
+ experiarSoC_videoSRAM0/dout1[22] experiarSoC_videoSRAM0/dout1[23] experiarSoC_videoSRAM0/dout1[24]
+ experiarSoC_videoSRAM0/dout1[25] experiarSoC_videoSRAM0/dout1[26] experiarSoC_videoSRAM0/dout1[27]
+ experiarSoC_videoSRAM0/dout1[28] experiarSoC_videoSRAM0/dout1[29] experiarSoC_videoSRAM0/dout1[2]
+ experiarSoC_videoSRAM0/dout1[30] experiarSoC_videoSRAM0/dout1[31] experiarSoC_videoSRAM1/dout1[0]
+ experiarSoC_videoSRAM1/dout1[1] experiarSoC_videoSRAM1/dout1[2] experiarSoC_videoSRAM1/dout1[3]
+ experiarSoC_videoSRAM1/dout1[4] experiarSoC_videoSRAM1/dout1[5] experiarSoC_videoSRAM1/dout1[6]
+ experiarSoC_videoSRAM1/dout1[7] experiarSoC_videoSRAM0/dout1[3] experiarSoC_videoSRAM1/dout1[8]
+ experiarSoC_videoSRAM1/dout1[9] experiarSoC_videoSRAM1/dout1[10] experiarSoC_videoSRAM1/dout1[11]
+ experiarSoC_videoSRAM1/dout1[12] experiarSoC_videoSRAM1/dout1[13] experiarSoC_videoSRAM1/dout1[14]
+ experiarSoC_videoSRAM1/dout1[15] experiarSoC_videoSRAM1/dout1[16] experiarSoC_videoSRAM1/dout1[17]
+ experiarSoC_videoSRAM0/dout1[4] experiarSoC_videoSRAM1/dout1[18] experiarSoC_videoSRAM1/dout1[19]
+ experiarSoC_videoSRAM1/dout1[20] experiarSoC_videoSRAM1/dout1[21] experiarSoC_videoSRAM1/dout1[22]
+ experiarSoC_videoSRAM1/dout1[23] experiarSoC_videoSRAM1/dout1[24] experiarSoC_videoSRAM1/dout1[25]
+ experiarSoC_videoSRAM1/dout1[26] experiarSoC_videoSRAM1/dout1[27] experiarSoC_videoSRAM0/dout1[5]
+ experiarSoC_videoSRAM1/dout1[28] experiarSoC_videoSRAM1/dout1[29] experiarSoC_videoSRAM1/dout1[30]
+ experiarSoC_videoSRAM1/dout1[31] experiarSoC_videoSRAM0/dout1[6] experiarSoC_videoSRAM0/dout1[7]
+ experiarSoC_videoSRAM0/dout1[8] experiarSoC_videoSRAM0/dout1[9] experiarSoC_videoSRAM1/web0
+ experiarSoC_videoSRAM1/wmask0[0] experiarSoC_videoSRAM1/wmask0[1] experiarSoC_videoSRAM1/wmask0[2]
+ experiarSoC_videoSRAM1/wmask0[3] experiarSoC_videoSRAM3/addr0[0] experiarSoC_videoSRAM3/addr0[1]
+ experiarSoC_videoSRAM3/addr0[2] experiarSoC_videoSRAM3/addr0[3] experiarSoC_videoSRAM3/addr0[4]
+ experiarSoC_videoSRAM3/addr0[5] experiarSoC_videoSRAM3/addr0[6] experiarSoC_videoSRAM3/addr0[7]
+ experiarSoC_videoSRAM3/addr0[8] experiarSoC_videoSRAM3/addr1[0] experiarSoC_videoSRAM3/addr1[1]
+ experiarSoC_videoSRAM3/addr1[2] experiarSoC_videoSRAM3/addr1[3] experiarSoC_videoSRAM3/addr1[4]
+ experiarSoC_videoSRAM3/addr1[5] experiarSoC_videoSRAM3/addr1[6] experiarSoC_videoSRAM3/addr1[7]
+ experiarSoC_videoSRAM3/addr1[8] experiarSoC_videoSRAM3/clk0 experiarSoC_videoSRAM3/clk1
+ experiarSoC_videoSRAM2/csb0 experiarSoC_videoSRAM3/csb0 experiarSoC_videoSRAM2/csb1
+ experiarSoC_videoSRAM3/csb1 experiarSoC_videoSRAM3/din0[0] experiarSoC_videoSRAM3/din0[10]
+ experiarSoC_videoSRAM3/din0[11] experiarSoC_videoSRAM3/din0[12] experiarSoC_videoSRAM3/din0[13]
+ experiarSoC_videoSRAM3/din0[14] experiarSoC_videoSRAM3/din0[15] experiarSoC_videoSRAM3/din0[16]
+ experiarSoC_videoSRAM3/din0[17] experiarSoC_videoSRAM3/din0[18] experiarSoC_videoSRAM3/din0[19]
+ experiarSoC_videoSRAM3/din0[1] experiarSoC_videoSRAM3/din0[20] experiarSoC_videoSRAM3/din0[21]
+ experiarSoC_videoSRAM3/din0[22] experiarSoC_videoSRAM3/din0[23] experiarSoC_videoSRAM3/din0[24]
+ experiarSoC_videoSRAM3/din0[25] experiarSoC_videoSRAM3/din0[26] experiarSoC_videoSRAM3/din0[27]
+ experiarSoC_videoSRAM3/din0[28] experiarSoC_videoSRAM3/din0[29] experiarSoC_videoSRAM3/din0[2]
+ experiarSoC_videoSRAM3/din0[30] experiarSoC_videoSRAM3/din0[31] experiarSoC_videoSRAM3/din0[3]
+ experiarSoC_videoSRAM3/din0[4] experiarSoC_videoSRAM3/din0[5] experiarSoC_videoSRAM3/din0[6]
+ experiarSoC_videoSRAM3/din0[7] experiarSoC_videoSRAM3/din0[8] experiarSoC_videoSRAM3/din0[9]
+ experiarSoC_videoSRAM2/dout0[0] experiarSoC_videoSRAM2/dout0[10] experiarSoC_videoSRAM2/dout0[11]
+ experiarSoC_videoSRAM2/dout0[12] experiarSoC_videoSRAM2/dout0[13] experiarSoC_videoSRAM2/dout0[14]
+ experiarSoC_videoSRAM2/dout0[15] experiarSoC_videoSRAM2/dout0[16] experiarSoC_videoSRAM2/dout0[17]
+ experiarSoC_videoSRAM2/dout0[18] experiarSoC_videoSRAM2/dout0[19] experiarSoC_videoSRAM2/dout0[1]
+ experiarSoC_videoSRAM2/dout0[20] experiarSoC_videoSRAM2/dout0[21] experiarSoC_videoSRAM2/dout0[22]
+ experiarSoC_videoSRAM2/dout0[23] experiarSoC_videoSRAM2/dout0[24] experiarSoC_videoSRAM2/dout0[25]
+ experiarSoC_videoSRAM2/dout0[26] experiarSoC_videoSRAM2/dout0[27] experiarSoC_videoSRAM2/dout0[28]
+ experiarSoC_videoSRAM2/dout0[29] experiarSoC_videoSRAM2/dout0[2] experiarSoC_videoSRAM2/dout0[30]
+ experiarSoC_videoSRAM2/dout0[31] experiarSoC_videoSRAM3/dout0[0] experiarSoC_videoSRAM3/dout0[1]
+ experiarSoC_videoSRAM3/dout0[2] experiarSoC_videoSRAM3/dout0[3] experiarSoC_videoSRAM3/dout0[4]
+ experiarSoC_videoSRAM3/dout0[5] experiarSoC_videoSRAM3/dout0[6] experiarSoC_videoSRAM3/dout0[7]
+ experiarSoC_videoSRAM2/dout0[3] experiarSoC_videoSRAM3/dout0[8] experiarSoC_videoSRAM3/dout0[9]
+ experiarSoC_videoSRAM3/dout0[10] experiarSoC_videoSRAM3/dout0[11] experiarSoC_videoSRAM3/dout0[12]
+ experiarSoC_videoSRAM3/dout0[13] experiarSoC_videoSRAM3/dout0[14] experiarSoC_videoSRAM3/dout0[15]
+ experiarSoC_videoSRAM3/dout0[16] experiarSoC_videoSRAM3/dout0[17] experiarSoC_videoSRAM2/dout0[4]
+ experiarSoC_videoSRAM3/dout0[18] experiarSoC_videoSRAM3/dout0[19] experiarSoC_videoSRAM3/dout0[20]
+ experiarSoC_videoSRAM3/dout0[21] experiarSoC_videoSRAM3/dout0[22] experiarSoC_videoSRAM3/dout0[23]
+ experiarSoC_videoSRAM3/dout0[24] experiarSoC_videoSRAM3/dout0[25] experiarSoC_videoSRAM3/dout0[26]
+ experiarSoC_videoSRAM3/dout0[27] experiarSoC_videoSRAM2/dout0[5] experiarSoC_videoSRAM3/dout0[28]
+ experiarSoC_videoSRAM3/dout0[29] experiarSoC_videoSRAM3/dout0[30] experiarSoC_videoSRAM3/dout0[31]
+ experiarSoC_videoSRAM2/dout0[6] experiarSoC_videoSRAM2/dout0[7] experiarSoC_videoSRAM2/dout0[8]
+ experiarSoC_videoSRAM2/dout0[9] experiarSoC_videoSRAM2/dout1[0] experiarSoC_videoSRAM2/dout1[10]
+ experiarSoC_videoSRAM2/dout1[11] experiarSoC_videoSRAM2/dout1[12] experiarSoC_videoSRAM2/dout1[13]
+ experiarSoC_videoSRAM2/dout1[14] experiarSoC_videoSRAM2/dout1[15] experiarSoC_videoSRAM2/dout1[16]
+ experiarSoC_videoSRAM2/dout1[17] experiarSoC_videoSRAM2/dout1[18] experiarSoC_videoSRAM2/dout1[19]
+ experiarSoC_videoSRAM2/dout1[1] experiarSoC_videoSRAM2/dout1[20] experiarSoC_videoSRAM2/dout1[21]
+ experiarSoC_videoSRAM2/dout1[22] experiarSoC_videoSRAM2/dout1[23] experiarSoC_videoSRAM2/dout1[24]
+ experiarSoC_videoSRAM2/dout1[25] experiarSoC_videoSRAM2/dout1[26] experiarSoC_videoSRAM2/dout1[27]
+ experiarSoC_videoSRAM2/dout1[28] experiarSoC_videoSRAM2/dout1[29] experiarSoC_videoSRAM2/dout1[2]
+ experiarSoC_videoSRAM2/dout1[30] experiarSoC_videoSRAM2/dout1[31] experiarSoC_videoSRAM3/dout1[0]
+ experiarSoC_videoSRAM3/dout1[1] experiarSoC_videoSRAM3/dout1[2] experiarSoC_videoSRAM3/dout1[3]
+ experiarSoC_videoSRAM3/dout1[4] experiarSoC_videoSRAM3/dout1[5] experiarSoC_videoSRAM3/dout1[6]
+ experiarSoC_videoSRAM3/dout1[7] experiarSoC_videoSRAM2/dout1[3] experiarSoC_videoSRAM3/dout1[8]
+ experiarSoC_videoSRAM3/dout1[9] experiarSoC_videoSRAM3/dout1[10] experiarSoC_videoSRAM3/dout1[11]
+ experiarSoC_videoSRAM3/dout1[12] experiarSoC_videoSRAM3/dout1[13] experiarSoC_videoSRAM3/dout1[14]
+ experiarSoC_videoSRAM3/dout1[15] experiarSoC_videoSRAM3/dout1[16] experiarSoC_videoSRAM3/dout1[17]
+ experiarSoC_videoSRAM2/dout1[4] experiarSoC_videoSRAM3/dout1[18] experiarSoC_videoSRAM3/dout1[19]
+ experiarSoC_videoSRAM3/dout1[20] experiarSoC_videoSRAM3/dout1[21] experiarSoC_videoSRAM3/dout1[22]
+ experiarSoC_videoSRAM3/dout1[23] experiarSoC_videoSRAM3/dout1[24] experiarSoC_videoSRAM3/dout1[25]
+ experiarSoC_videoSRAM3/dout1[26] experiarSoC_videoSRAM3/dout1[27] experiarSoC_videoSRAM2/dout1[5]
+ experiarSoC_videoSRAM3/dout1[28] experiarSoC_videoSRAM3/dout1[29] experiarSoC_videoSRAM3/dout1[30]
+ experiarSoC_videoSRAM3/dout1[31] experiarSoC_videoSRAM2/dout1[6] experiarSoC_videoSRAM2/dout1[7]
+ experiarSoC_videoSRAM2/dout1[8] experiarSoC_videoSRAM2/dout1[9] experiarSoC_videoSRAM3/web0
+ experiarSoC_videoSRAM3/wmask0[0] experiarSoC_videoSRAM3/wmask0[1] experiarSoC_videoSRAM3/wmask0[2]
+ experiarSoC_videoSRAM3/wmask0[3] vccd1 experiarSoC_video/vga_b[0] experiarSoC_video/vga_b[1]
+ experiarSoC_video/vga_g[0] experiarSoC_video/vga_g[1] experiarSoC_video/vga_hsync
+ experiarSoC_video/vga_r[0] experiarSoC_video/vga_r[1] experiarSoC_video/vga_vsync
+ experiarSoC_core1/irq[10] experiarSoC_core1/irq[11] vssd1 experiarSoC_video/wb_ack_o
+ experiarSoC_video/wb_adr_i[0] experiarSoC_video/wb_adr_i[10] experiarSoC_video/wb_adr_i[11]
+ experiarSoC_video/wb_adr_i[12] experiarSoC_video/wb_adr_i[13] experiarSoC_video/wb_adr_i[14]
+ experiarSoC_video/wb_adr_i[15] experiarSoC_video/wb_adr_i[16] experiarSoC_video/wb_adr_i[17]
+ experiarSoC_video/wb_adr_i[18] experiarSoC_video/wb_adr_i[19] experiarSoC_video/wb_adr_i[1]
+ experiarSoC_video/wb_adr_i[20] experiarSoC_video/wb_adr_i[21] experiarSoC_video/wb_adr_i[22]
+ experiarSoC_video/wb_adr_i[23] experiarSoC_video/wb_adr_i[2] experiarSoC_video/wb_adr_i[3]
+ experiarSoC_video/wb_adr_i[4] experiarSoC_video/wb_adr_i[5] experiarSoC_video/wb_adr_i[6]
+ experiarSoC_video/wb_adr_i[7] experiarSoC_video/wb_adr_i[8] experiarSoC_video/wb_adr_i[9]
+ wb_clk_i experiarSoC_video/wb_cyc_i experiarSoC_video/wb_data_i[0] experiarSoC_video/wb_data_i[10]
+ experiarSoC_video/wb_data_i[11] experiarSoC_video/wb_data_i[12] experiarSoC_video/wb_data_i[13]
+ experiarSoC_video/wb_data_i[14] experiarSoC_video/wb_data_i[15] experiarSoC_video/wb_data_i[16]
+ experiarSoC_video/wb_data_i[17] experiarSoC_video/wb_data_i[18] experiarSoC_video/wb_data_i[19]
+ experiarSoC_video/wb_data_i[1] experiarSoC_video/wb_data_i[20] experiarSoC_video/wb_data_i[21]
+ experiarSoC_video/wb_data_i[22] experiarSoC_video/wb_data_i[23] experiarSoC_video/wb_data_i[24]
+ experiarSoC_video/wb_data_i[25] experiarSoC_video/wb_data_i[26] experiarSoC_video/wb_data_i[27]
+ experiarSoC_video/wb_data_i[28] experiarSoC_video/wb_data_i[29] experiarSoC_video/wb_data_i[2]
+ experiarSoC_video/wb_data_i[30] experiarSoC_video/wb_data_i[31] experiarSoC_video/wb_data_i[3]
+ experiarSoC_video/wb_data_i[4] experiarSoC_video/wb_data_i[5] experiarSoC_video/wb_data_i[6]
+ experiarSoC_video/wb_data_i[7] experiarSoC_video/wb_data_i[8] experiarSoC_video/wb_data_i[9]
+ experiarSoC_video/wb_data_o[0] experiarSoC_video/wb_data_o[10] experiarSoC_video/wb_data_o[11]
+ experiarSoC_video/wb_data_o[12] experiarSoC_video/wb_data_o[13] experiarSoC_video/wb_data_o[14]
+ experiarSoC_video/wb_data_o[15] experiarSoC_video/wb_data_o[16] experiarSoC_video/wb_data_o[17]
+ experiarSoC_video/wb_data_o[18] experiarSoC_video/wb_data_o[19] experiarSoC_video/wb_data_o[1]
+ experiarSoC_video/wb_data_o[20] experiarSoC_video/wb_data_o[21] experiarSoC_video/wb_data_o[22]
+ experiarSoC_video/wb_data_o[23] experiarSoC_video/wb_data_o[24] experiarSoC_video/wb_data_o[25]
+ experiarSoC_video/wb_data_o[26] experiarSoC_video/wb_data_o[27] experiarSoC_video/wb_data_o[28]
+ experiarSoC_video/wb_data_o[29] experiarSoC_video/wb_data_o[2] experiarSoC_video/wb_data_o[30]
+ experiarSoC_video/wb_data_o[31] experiarSoC_video/wb_data_o[3] experiarSoC_video/wb_data_o[4]
+ experiarSoC_video/wb_data_o[5] experiarSoC_video/wb_data_o[6] experiarSoC_video/wb_data_o[7]
+ experiarSoC_video/wb_data_o[8] experiarSoC_video/wb_data_o[9] experiarSoC_video/wb_error_o
+ wb_rst_i experiarSoC_video/wb_sel_i[0] experiarSoC_video/wb_sel_i[1] experiarSoC_video/wb_sel_i[2]
+ experiarSoC_video/wb_sel_i[3] experiarSoC_video/wb_stall_o experiarSoC_video/wb_stb_i
+ experiarSoC_video/wb_we_i Video
XexperiarSoC_flash experiarSoC_flash/flash_csb experiarSoC_flash/flash_io0_read experiarSoC_flash/flash_io0_we
+ experiarSoC_flash/flash_io0_write experiarSoC_flash/flash_io1_read experiarSoC_flash/flash_io1_we
+ experiarSoC_flash/flash_io1_write experiarSoC_flash/flash_sck experiarSoC_flashSRAM/addr0[0]
+ experiarSoC_flashSRAM/addr0[1] experiarSoC_flashSRAM/addr0[2] experiarSoC_flashSRAM/addr0[3]
+ experiarSoC_flashSRAM/addr0[4] experiarSoC_flashSRAM/addr0[5] experiarSoC_flashSRAM/addr0[6]
+ experiarSoC_flashSRAM/addr0[7] experiarSoC_flashSRAM/addr0[8] experiarSoC_flashSRAM/addr1[0]
+ experiarSoC_flashSRAM/addr1[1] experiarSoC_flashSRAM/addr1[2] experiarSoC_flashSRAM/addr1[3]
+ experiarSoC_flashSRAM/addr1[4] experiarSoC_flashSRAM/addr1[5] experiarSoC_flashSRAM/addr1[6]
+ experiarSoC_flashSRAM/addr1[7] experiarSoC_flashSRAM/addr1[8] experiarSoC_flashSRAM/clk0
+ experiarSoC_flashSRAM/clk1 experiarSoC_flashSRAM/csb0 experiarSoC_flashSRAM/csb1
+ experiarSoC_flashSRAM/din0[0] experiarSoC_flashSRAM/din0[10] experiarSoC_flashSRAM/din0[11]
+ experiarSoC_flashSRAM/din0[12] experiarSoC_flashSRAM/din0[13] experiarSoC_flashSRAM/din0[14]
+ experiarSoC_flashSRAM/din0[15] experiarSoC_flashSRAM/din0[16] experiarSoC_flashSRAM/din0[17]
+ experiarSoC_flashSRAM/din0[18] experiarSoC_flashSRAM/din0[19] experiarSoC_flashSRAM/din0[1]
+ experiarSoC_flashSRAM/din0[20] experiarSoC_flashSRAM/din0[21] experiarSoC_flashSRAM/din0[22]
+ experiarSoC_flashSRAM/din0[23] experiarSoC_flashSRAM/din0[24] experiarSoC_flashSRAM/din0[25]
+ experiarSoC_flashSRAM/din0[26] experiarSoC_flashSRAM/din0[27] experiarSoC_flashSRAM/din0[28]
+ experiarSoC_flashSRAM/din0[29] experiarSoC_flashSRAM/din0[2] experiarSoC_flashSRAM/din0[30]
+ experiarSoC_flashSRAM/din0[31] experiarSoC_flashSRAM/din0[3] experiarSoC_flashSRAM/din0[4]
+ experiarSoC_flashSRAM/din0[5] experiarSoC_flashSRAM/din0[6] experiarSoC_flashSRAM/din0[7]
+ experiarSoC_flashSRAM/din0[8] experiarSoC_flashSRAM/din0[9] experiarSoC_flashSRAM/dout0[0]
+ experiarSoC_flashSRAM/dout0[10] experiarSoC_flashSRAM/dout0[11] experiarSoC_flashSRAM/dout0[12]
+ experiarSoC_flashSRAM/dout0[13] experiarSoC_flashSRAM/dout0[14] experiarSoC_flashSRAM/dout0[15]
+ experiarSoC_flashSRAM/dout0[16] experiarSoC_flashSRAM/dout0[17] experiarSoC_flashSRAM/dout0[18]
+ experiarSoC_flashSRAM/dout0[19] experiarSoC_flashSRAM/dout0[1] experiarSoC_flashSRAM/dout0[20]
+ experiarSoC_flashSRAM/dout0[21] experiarSoC_flashSRAM/dout0[22] experiarSoC_flashSRAM/dout0[23]
+ experiarSoC_flashSRAM/dout0[24] experiarSoC_flashSRAM/dout0[25] experiarSoC_flashSRAM/dout0[26]
+ experiarSoC_flashSRAM/dout0[27] experiarSoC_flashSRAM/dout0[28] experiarSoC_flashSRAM/dout0[29]
+ experiarSoC_flashSRAM/dout0[2] experiarSoC_flashSRAM/dout0[30] experiarSoC_flashSRAM/dout0[31]
+ experiarSoC_flashSRAM/dout0[3] experiarSoC_flashSRAM/dout0[4] experiarSoC_flashSRAM/dout0[5]
+ experiarSoC_flashSRAM/dout0[6] experiarSoC_flashSRAM/dout0[7] experiarSoC_flashSRAM/dout0[8]
+ experiarSoC_flashSRAM/dout0[9] experiarSoC_flashSRAM/dout1[0] experiarSoC_flashSRAM/dout1[10]
+ experiarSoC_flashSRAM/dout1[11] experiarSoC_flashSRAM/dout1[12] experiarSoC_flashSRAM/dout1[13]
+ experiarSoC_flashSRAM/dout1[14] experiarSoC_flashSRAM/dout1[15] experiarSoC_flashSRAM/dout1[16]
+ experiarSoC_flashSRAM/dout1[17] experiarSoC_flashSRAM/dout1[18] experiarSoC_flashSRAM/dout1[19]
+ experiarSoC_flashSRAM/dout1[1] experiarSoC_flashSRAM/dout1[20] experiarSoC_flashSRAM/dout1[21]
+ experiarSoC_flashSRAM/dout1[22] experiarSoC_flashSRAM/dout1[23] experiarSoC_flashSRAM/dout1[24]
+ experiarSoC_flashSRAM/dout1[25] experiarSoC_flashSRAM/dout1[26] experiarSoC_flashSRAM/dout1[27]
+ experiarSoC_flashSRAM/dout1[28] experiarSoC_flashSRAM/dout1[29] experiarSoC_flashSRAM/dout1[2]
+ experiarSoC_flashSRAM/dout1[30] experiarSoC_flashSRAM/dout1[31] experiarSoC_flashSRAM/dout1[3]
+ experiarSoC_flashSRAM/dout1[4] experiarSoC_flashSRAM/dout1[5] experiarSoC_flashSRAM/dout1[6]
+ experiarSoC_flashSRAM/dout1[7] experiarSoC_flashSRAM/dout1[8] experiarSoC_flashSRAM/dout1[9]
+ experiarSoC_flashSRAM/web0 experiarSoC_flashSRAM/wmask0[0] experiarSoC_flashSRAM/wmask0[1]
+ experiarSoC_flashSRAM/wmask0[2] experiarSoC_flashSRAM/wmask0[3] vccd1 vssd1 experiarSoC_flash/wb_ack_o
+ experiarSoC_flash/wb_adr_i[0] experiarSoC_flash/wb_adr_i[10] experiarSoC_flash/wb_adr_i[11]
+ experiarSoC_flash/wb_adr_i[12] experiarSoC_flash/wb_adr_i[13] experiarSoC_flash/wb_adr_i[14]
+ experiarSoC_flash/wb_adr_i[15] experiarSoC_flash/wb_adr_i[16] experiarSoC_flash/wb_adr_i[17]
+ experiarSoC_flash/wb_adr_i[18] experiarSoC_flash/wb_adr_i[19] experiarSoC_flash/wb_adr_i[1]
+ experiarSoC_flash/wb_adr_i[20] experiarSoC_flash/wb_adr_i[21] experiarSoC_flash/wb_adr_i[22]
+ experiarSoC_flash/wb_adr_i[23] experiarSoC_flash/wb_adr_i[2] experiarSoC_flash/wb_adr_i[3]
+ experiarSoC_flash/wb_adr_i[4] experiarSoC_flash/wb_adr_i[5] experiarSoC_flash/wb_adr_i[6]
+ experiarSoC_flash/wb_adr_i[7] experiarSoC_flash/wb_adr_i[8] experiarSoC_flash/wb_adr_i[9]
+ wb_clk_i experiarSoC_flash/wb_cyc_i experiarSoC_flash/wb_data_i[0] experiarSoC_flash/wb_data_i[10]
+ experiarSoC_flash/wb_data_i[11] experiarSoC_flash/wb_data_i[12] experiarSoC_flash/wb_data_i[13]
+ experiarSoC_flash/wb_data_i[14] experiarSoC_flash/wb_data_i[15] experiarSoC_flash/wb_data_i[16]
+ experiarSoC_flash/wb_data_i[17] experiarSoC_flash/wb_data_i[18] experiarSoC_flash/wb_data_i[19]
+ experiarSoC_flash/wb_data_i[1] experiarSoC_flash/wb_data_i[20] experiarSoC_flash/wb_data_i[21]
+ experiarSoC_flash/wb_data_i[22] experiarSoC_flash/wb_data_i[23] experiarSoC_flash/wb_data_i[24]
+ experiarSoC_flash/wb_data_i[25] experiarSoC_flash/wb_data_i[26] experiarSoC_flash/wb_data_i[27]
+ experiarSoC_flash/wb_data_i[28] experiarSoC_flash/wb_data_i[29] experiarSoC_flash/wb_data_i[2]
+ experiarSoC_flash/wb_data_i[30] experiarSoC_flash/wb_data_i[31] experiarSoC_flash/wb_data_i[3]
+ experiarSoC_flash/wb_data_i[4] experiarSoC_flash/wb_data_i[5] experiarSoC_flash/wb_data_i[6]
+ experiarSoC_flash/wb_data_i[7] experiarSoC_flash/wb_data_i[8] experiarSoC_flash/wb_data_i[9]
+ experiarSoC_flash/wb_data_o[0] experiarSoC_flash/wb_data_o[10] experiarSoC_flash/wb_data_o[11]
+ experiarSoC_flash/wb_data_o[12] experiarSoC_flash/wb_data_o[13] experiarSoC_flash/wb_data_o[14]
+ experiarSoC_flash/wb_data_o[15] experiarSoC_flash/wb_data_o[16] experiarSoC_flash/wb_data_o[17]
+ experiarSoC_flash/wb_data_o[18] experiarSoC_flash/wb_data_o[19] experiarSoC_flash/wb_data_o[1]
+ experiarSoC_flash/wb_data_o[20] experiarSoC_flash/wb_data_o[21] experiarSoC_flash/wb_data_o[22]
+ experiarSoC_flash/wb_data_o[23] experiarSoC_flash/wb_data_o[24] experiarSoC_flash/wb_data_o[25]
+ experiarSoC_flash/wb_data_o[26] experiarSoC_flash/wb_data_o[27] experiarSoC_flash/wb_data_o[28]
+ experiarSoC_flash/wb_data_o[29] experiarSoC_flash/wb_data_o[2] experiarSoC_flash/wb_data_o[30]
+ experiarSoC_flash/wb_data_o[31] experiarSoC_flash/wb_data_o[3] experiarSoC_flash/wb_data_o[4]
+ experiarSoC_flash/wb_data_o[5] experiarSoC_flash/wb_data_o[6] experiarSoC_flash/wb_data_o[7]
+ experiarSoC_flash/wb_data_o[8] experiarSoC_flash/wb_data_o[9] experiarSoC_flash/wb_error_o
+ wb_rst_i experiarSoC_flash/wb_sel_i[0] experiarSoC_flash/wb_sel_i[1] experiarSoC_flash/wb_sel_i[2]
+ experiarSoC_flash/wb_sel_i[3] experiarSoC_flash/wb_stall_o experiarSoC_flash/wb_stb_i
+ experiarSoC_flash/wb_we_i Flash
.ends

