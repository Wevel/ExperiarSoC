* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt CaravelHost caravel_uart_rx caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0]
+ caravel_wb_adr_o[10] caravel_wb_adr_o[11] caravel_wb_adr_o[12] caravel_wb_adr_o[13]
+ caravel_wb_adr_o[14] caravel_wb_adr_o[15] caravel_wb_adr_o[16] caravel_wb_adr_o[17]
+ caravel_wb_adr_o[18] caravel_wb_adr_o[19] caravel_wb_adr_o[1] caravel_wb_adr_o[20]
+ caravel_wb_adr_o[21] caravel_wb_adr_o[22] caravel_wb_adr_o[23] caravel_wb_adr_o[24]
+ caravel_wb_adr_o[25] caravel_wb_adr_o[26] caravel_wb_adr_o[27] caravel_wb_adr_o[2]
+ caravel_wb_adr_o[3] caravel_wb_adr_o[4] caravel_wb_adr_o[5] caravel_wb_adr_o[6]
+ caravel_wb_adr_o[7] caravel_wb_adr_o[8] caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0]
+ caravel_wb_data_i[10] caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13]
+ caravel_wb_data_i[14] caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17]
+ caravel_wb_data_i[18] caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20]
+ caravel_wb_data_i[21] caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24]
+ caravel_wb_data_i[25] caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28]
+ caravel_wb_data_i[29] caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31]
+ caravel_wb_data_i[3] caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6]
+ caravel_wb_data_i[7] caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0]
+ caravel_wb_data_o[10] caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13]
+ caravel_wb_data_o[14] caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17]
+ caravel_wb_data_o[18] caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20]
+ caravel_wb_data_o[21] caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24]
+ caravel_wb_data_o[25] caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28]
+ caravel_wb_data_o[29] caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31]
+ caravel_wb_data_o[3] caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6]
+ caravel_wb_data_o[7] caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i
+ caravel_wb_sel_o[0] caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3]
+ caravel_wb_stall_i caravel_wb_stb_o caravel_wb_we_o core0Index[0] core0Index[1]
+ core0Index[2] core0Index[3] core0Index[4] core0Index[5] core0Index[6] core0Index[7]
+ core1Index[0] core1Index[1] core1Index[2] core1Index[3] core1Index[4] core1Index[5]
+ core1Index[6] core1Index[7] manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] vccd1 versionID[0] versionID[1]
+ versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12] wbs_data_i[13] wbs_data_i[14]
+ wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18] wbs_data_i[19] wbs_data_i[1]
+ wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23] wbs_data_i[24] wbs_data_i[25]
+ wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29] wbs_data_i[2] wbs_data_i[30]
+ wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5] wbs_data_i[6] wbs_data_i[7]
+ wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10] wbs_data_o[11] wbs_data_o[12]
+ wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16] wbs_data_o[17] wbs_data_o[18]
+ wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21] wbs_data_o[22] wbs_data_o[23]
+ wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27] wbs_data_o[28] wbs_data_o[29]
+ wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3] wbs_data_o[4] wbs_data_o[5]
+ wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_100_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7963_ _7963_/CLK _7963_/D vssd1 vssd1 vccd1 vccd1 _7963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7894_ _7894_/CLK _7894_/D vssd1 vssd1 vccd1 vccd1 _7894_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2973_ _6082_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2973_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6845_ _6845_/A vssd1 vssd1 vccd1 vccd1 _6845_/X sky130_fd_sc_hd__buf_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3988_ _4368_/A vssd1 vssd1 vccd1 vccd1 _5511_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5727_ _7772_/Q _5547_/A _5735_/S vssd1 vssd1 vccd1 vccd1 _5728_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5658_ _5658_/A vssd1 vssd1 vccd1 vccd1 _7803_/D sky130_fd_sc_hd__clkbuf_1
X_4609_ _6910_/A vssd1 vssd1 vccd1 vccd1 _4609_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5589_ _5589_/A vssd1 vssd1 vccd1 vccd1 _7832_/D sky130_fd_sc_hd__clkbuf_1
X_8377_ _8377_/CLK _8377_/D vssd1 vssd1 vccd1 vccd1 _8377_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3387_ _6944_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3387_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7259_ _7262_/B _7262_/C _7262_/D vssd1 vssd1 vccd1 vccd1 _7259_/X sky130_fd_sc_hd__or3b_1
XFILLER_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6882__450 _6882__450/A vssd1 vssd1 vccd1 vccd1 _8045_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3207_ clkbuf_0__3207_/X vssd1 vssd1 vccd1 vccd1 _6511__282/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6930__484 _6931__485/A vssd1 vssd1 vccd1 vccd1 _8081_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6972__518 _6974__520/A vssd1 vssd1 vccd1 vccd1 _8115_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4960_ _7993_/Q vssd1 vssd1 vccd1 vccd1 _5100_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3911_ _3890_/X _8321_/Q _3911_/S vssd1 vssd1 vccd1 vccd1 _3912_/A sky130_fd_sc_hd__mux2_1
X_4891_ _8038_/Q _4410_/X _4891_/S vssd1 vssd1 vccd1 vccd1 _4892_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3842_ _3842_/A vssd1 vssd1 vccd1 vccd1 _8382_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _7066__93/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6561_ _6561_/A vssd1 vssd1 vccd1 vccd1 _7863_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3342_ clkbuf_0__3342_/X vssd1 vssd1 vccd1 vccd1 _6792_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3773_ _8002_/Q vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5527_/S vssd1 vssd1 vccd1 vccd1 _5521_/S sky130_fd_sc_hd__buf_2
X_8300_ _8300_/CLK _8300_/D vssd1 vssd1 vccd1 vccd1 _8300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8231_ _8231_/CLK _8231_/D vssd1 vssd1 vccd1 vccd1 _8231_/Q sky130_fd_sc_hd__dfxtp_1
X_5443_ _3822_/X _7915_/Q _5449_/S vssd1 vssd1 vccd1 vccd1 _5444_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3241_ _6587_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3241_/X sky130_fd_sc_hd__clkbuf_16
X_5374_ _5374_/A vssd1 vssd1 vccd1 vccd1 _7949_/D sky130_fd_sc_hd__clkbuf_1
X_8162_ _8162_/CLK _8162_/D vssd1 vssd1 vccd1 vccd1 _8162_/Q sky130_fd_sc_hd__dfxtp_1
X_7113_ _8224_/Q vssd1 vssd1 vccd1 vccd1 _7113_/Y sky130_fd_sc_hd__inv_2
X_4325_ _5599_/A _5653_/B vssd1 vssd1 vccd1 vccd1 _4348_/S sky130_fd_sc_hd__or2_2
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8093_ _8093_/CLK _8093_/D vssd1 vssd1 vccd1 vccd1 _8093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4256_ _4211_/X _8176_/Q _4260_/S vssd1 vssd1 vccd1 vccd1 _4257_/A sky130_fd_sc_hd__mux2_1
X_7044_ _7075_/A vssd1 vssd1 vccd1 vccd1 _7044_/X sky130_fd_sc_hd__buf_1
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4187_ _4202_/S vssd1 vssd1 vccd1 vccd1 _4196_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7946_ _7946_/CLK _7946_/D vssd1 vssd1 vccd1 vccd1 _7946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7877_ _7877_/CLK _7877_/D vssd1 vssd1 vccd1 vccd1 _7877_/Q sky130_fd_sc_hd__dfxtp_1
X_6828_ _6834_/A vssd1 vssd1 vccd1 vccd1 _6828_/X sky130_fd_sc_hd__buf_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6759_ _7593_/A _7491_/A vssd1 vssd1 vccd1 vccd1 _7410_/B sky130_fd_sc_hd__xor2_1
X_7186__110 _7186__110/A vssd1 vssd1 vccd1 vccd1 _8209_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6477__255 _6477__255/A vssd1 vssd1 vccd1 vccd1 _7812_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5090_ _5090_/A vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__clkbuf_2
X_4110_ _8261_/Q _3947_/X _4112_/S vssd1 vssd1 vccd1 vccd1 _4111_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4041_ _4041_/A vssd1 vssd1 vccd1 vccd1 _8274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ _6400_/A vssd1 vssd1 vccd1 vccd1 _6006_/S sky130_fd_sc_hd__buf_2
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7800_ _7800_/CLK _7800_/D vssd1 vssd1 vccd1 vccd1 _7800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7731_ _8407_/CLK _7731_/D vssd1 vssd1 vccd1 vccd1 _7731_/Q sky130_fd_sc_hd__dfxtp_1
X_4943_ _4341_/X _8016_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__mux2_1
X_7662_ _7697_/CLK _7662_/D vssd1 vssd1 vccd1 vccd1 _7662_/Q sky130_fd_sc_hd__dfxtp_1
X_6421__210 _6421__210/A vssd1 vssd1 vccd1 vccd1 _7767_/CLK sky130_fd_sc_hd__inv_2
X_4874_ _4874_/A vssd1 vssd1 vccd1 vccd1 _8046_/D sky130_fd_sc_hd__clkbuf_1
X_6613_ _6613_/A vssd1 vssd1 vccd1 vccd1 _6613_/X sky130_fd_sc_hd__buf_1
X_7593_ _7593_/A _7599_/B vssd1 vssd1 vccd1 vccd1 _7593_/Y sky130_fd_sc_hd__nor2_1
X_3825_ _8363_/Q vssd1 vssd1 vccd1 vccd1 _3825_/X sky130_fd_sc_hd__buf_2
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6544_ _5877_/A _7856_/Q _6546_/S vssd1 vssd1 vccd1 vccd1 _6545_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3256_ clkbuf_0__3256_/X vssd1 vssd1 vccd1 vccd1 _6668__360/A sky130_fd_sc_hd__clkbuf_4
X_8214_ _8364_/CLK _8214_/D vssd1 vssd1 vccd1 vccd1 _8214_/Q sky130_fd_sc_hd__dfxtp_1
X_5426_ _5426_/A vssd1 vssd1 vccd1 vccd1 _7923_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3187_ clkbuf_0__3187_/X vssd1 vssd1 vccd1 vccd1 _6422_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8145_ _8145_/CLK _8145_/D vssd1 vssd1 vccd1 vccd1 _8145_/Q sky130_fd_sc_hd__dfxtp_1
X_5357_ _5357_/A vssd1 vssd1 vccd1 vccd1 _7956_/D sky130_fd_sc_hd__clkbuf_1
X_8426__201 vssd1 vssd1 vccd1 vccd1 _8426__201/HI core1Index[1] sky130_fd_sc_hd__conb_1
XFILLER_114_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _5555_/A vssd1 vssd1 vccd1 vccd1 _5288_/X sky130_fd_sc_hd__buf_2
X_4308_ _4308_/A vssd1 vssd1 vccd1 vccd1 _8154_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_4 _5973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8076_ _8076_/CLK _8076_/D vssd1 vssd1 vccd1 vccd1 _8076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4239_ _8183_/Q _4131_/X _4241_/S vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7929_ _7929_/CLK _7929_/D vssd1 vssd1 vccd1 vccd1 _7929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6773__380 _6773__380/A vssd1 vssd1 vccd1 vccd1 _7965_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6895__460 _6895__460/A vssd1 vssd1 vccd1 vccd1 _8055_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3402_ clkbuf_0__3402_/X vssd1 vssd1 vccd1 vccd1 _7019__55/A sky130_fd_sc_hd__clkbuf_16
XFILLER_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4590_ _8029_/Q _7984_/Q _7844_/Q _8212_/Q _4559_/A _4589_/X vssd1 vssd1 vccd1 vccd1
+ _4590_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _7422_/A _6249_/X _6251_/X _6228_/X vssd1 vssd1 vccd1 vccd1 _6260_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6191_ _8229_/Q vssd1 vssd1 vccd1 vccd1 _7258_/B sky130_fd_sc_hd__clkbuf_2
X_5211_ _5019_/X _5200_/X _5203_/X _5210_/X _5002_/X vssd1 vssd1 vccd1 vccd1 _5211_/X
+ sky130_fd_sc_hd__o311a_1
X_5142_ _5265_/B _5120_/X _5124_/X _5141_/X vssd1 vssd1 vccd1 vccd1 _5142_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5073_ _8009_/Q _4955_/X _5031_/X _5072_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _5073_/X
+ sky130_fd_sc_hd__a221o_1
X_6904__467 _6906__469/A vssd1 vssd1 vccd1 vccd1 _8062_/CLK sky130_fd_sc_hd__inv_2
X_4024_ _3890_/X _8281_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4025_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5975_ _6400_/A vssd1 vssd1 vccd1 vccd1 _5989_/S sky130_fd_sc_hd__buf_4
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7714_ _7989_/CLK _7714_/D vssd1 vssd1 vccd1 vccd1 _7714_/Q sky130_fd_sc_hd__dfxtp_1
X_4926_ _8023_/Q _4407_/X _4928_/S vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4857_ _4604_/A _4324_/A _6253_/A _4843_/A vssd1 vssd1 vccd1 vccd1 _4858_/B sky130_fd_sc_hd__a31o_1
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7645_ _7645_/CLK _7645_/D vssd1 vssd1 vccd1 vccd1 _7645_/Q sky130_fd_sc_hd__dfxtp_1
X_3808_ _7746_/Q _7747_/Q _7748_/Q _7749_/Q vssd1 vssd1 vccd1 vccd1 _6341_/B sky130_fd_sc_hd__or4_1
XFILLER_118_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6527_ _6527_/A vssd1 vssd1 vccd1 vccd1 _7848_/D sky130_fd_sc_hd__clkbuf_1
X_4788_ _8116_/Q _4705_/X _4593_/S _4787_/X vssd1 vssd1 vccd1 vccd1 _4789_/C sky130_fd_sc_hd__o211a_1
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6985__528 _6985__528/A vssd1 vssd1 vccd1 vccd1 _8125_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__2972_ clkbuf_0__2972_/X vssd1 vssd1 vccd1 vccd1 _6851_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3239_ clkbuf_0__3239_/X vssd1 vssd1 vccd1 vccd1 _6580__295/A sky130_fd_sc_hd__clkbuf_4
X_6389_ _7856_/Q _7749_/Q _6393_/S vssd1 vssd1 vccd1 vccd1 _6390_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _7930_/Q _4514_/X _5413_/S vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3207_ _6509_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3207_/X sky130_fd_sc_hd__clkbuf_16
X_8128_ _8128_/CLK _8128_/D vssd1 vssd1 vccd1 vccd1 _8128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8059_ _8059_/CLK _8059_/D vssd1 vssd1 vccd1 vccd1 _8059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7072__98 _7073__99/A vssd1 vssd1 vccd1 vccd1 _8195_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3590_ clkbuf_0__3590_/X vssd1 vssd1 vccd1 vccd1 _7357_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5760_ _5760_/A vssd1 vssd1 vccd1 vccd1 _7757_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _7788_/Q _5573_/X _5699_/S vssd1 vssd1 vccd1 vccd1 _5692_/A sky130_fd_sc_hd__mux2_1
X_4711_ _7792_/Q _4676_/X _4710_/X _4715_/A vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__o22a_1
XFILLER_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7430_ _7430_/A _7430_/B _7430_/C vssd1 vssd1 vccd1 vccd1 _7430_/X sky130_fd_sc_hd__and3_1
X_4642_ _4642_/A vssd1 vssd1 vccd1 vccd1 _4664_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _8049_/Q _4573_/B vssd1 vssd1 vccd1 vccd1 _4584_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6312_ _6312_/A vssd1 vssd1 vccd1 vccd1 _6326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6243_ _6289_/B vssd1 vssd1 vccd1 vccd1 _6243_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174_ _7629_/A _7697_/Q _6174_/S vssd1 vssd1 vccd1 vccd1 _6175_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5056_ _8379_/Q _7949_/Q _7882_/Q _8371_/Q _5198_/S _4971_/X vssd1 vssd1 vccd1 vccd1
+ _5056_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4007_ _4286_/B _4120_/C _4286_/A vssd1 vssd1 vccd1 vccd1 _4204_/B sky130_fd_sc_hd__or3b_4
Xclkbuf_1_0_0__3240_ clkbuf_0__3240_/X vssd1 vssd1 vccd1 vccd1 _6586__300/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _7861_/Q _5964_/B vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__and2_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _4909_/A vssd1 vssd1 vccd1 vccd1 _8031_/D sky130_fd_sc_hd__clkbuf_1
X_5889_ _5889_/A vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7628_ _7626_/Y _7627_/B _7627_/Y _6151_/X vssd1 vssd1 vccd1 vccd1 _8402_/D sky130_fd_sc_hd__a211oi_1
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6846__421 _6847__422/A vssd1 vssd1 vccd1 vccd1 _8016_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3369_ clkbuf_0__3369_/X vssd1 vssd1 vccd1 vccd1 _6864__435/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8407_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6792_ _6792_/A vssd1 vssd1 vccd1 vccd1 _6792_/X sky130_fd_sc_hd__buf_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5812_ _5812_/A vssd1 vssd1 vccd1 vccd1 _7645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5743_ _5743_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5759_/S sky130_fd_sc_hd__nor2_2
X_5674_ _5674_/A vssd1 vssd1 vccd1 vccd1 _7796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7413_ _7167_/A _6699_/B _6714_/B _7615_/A vssd1 vssd1 vccd1 vccd1 _7413_/Y sky130_fd_sc_hd__a22oi_1
X_8393_ _8399_/CLK _8393_/D vssd1 vssd1 vccd1 vccd1 _8393_/Q sky130_fd_sc_hd__dfxtp_1
X_4625_ _8201_/Q _7819_/Q _7803_/Q _7787_/Q _4595_/A _4559_/A vssd1 vssd1 vccd1 vccd1
+ _4625_/X sky130_fd_sc_hd__mux4_1
X_4556_ _4556_/A vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7275_ _8235_/Q _7277_/B vssd1 vssd1 vccd1 vccd1 _7275_/X sky130_fd_sc_hd__or2_1
X_4487_ _4487_/A vssd1 vssd1 vccd1 vccd1 _8083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6226_ _6237_/A _6226_/B _6226_/C _6309_/A vssd1 vssd1 vccd1 vccd1 _6285_/B sky130_fd_sc_hd__or4b_2
X_6157_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _8385_/Q _5108_/B vssd1 vssd1 vccd1 vccd1 _5108_/X sky130_fd_sc_hd__or2_1
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5039_ _8185_/Q _8177_/Q _7899_/Q _7915_/Q _5037_/X _5207_/S vssd1 vssd1 vccd1 vccd1
+ _5039_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6208__195 _6208__195/A vssd1 vssd1 vccd1 vccd1 _7707_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput97 _5935_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4410_ _7985_/Q vssd1 vssd1 vccd1 vccd1 _4410_/X sky130_fd_sc_hd__clkbuf_2
X_5390_ _5390_/A vssd1 vssd1 vccd1 vccd1 _7939_/D sky130_fd_sc_hd__clkbuf_1
X_4341_ _7987_/Q vssd1 vssd1 vccd1 vccd1 _4341_/X sky130_fd_sc_hd__buf_2
X_4272_ _8169_/Q _4125_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4273_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6011_ _6011_/A vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7962_ _7962_/CLK _7962_/D vssd1 vssd1 vccd1 vccd1 _7962_/Q sky130_fd_sc_hd__dfxtp_1
X_7018__54 _7019__55/A vssd1 vssd1 vccd1 vccd1 _8151_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6913_ _6913_/A vssd1 vssd1 vccd1 vccd1 _6913_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__2972_ _6081_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2972_/X sky130_fd_sc_hd__clkbuf_16
X_7893_ _7893_/CLK _7893_/D vssd1 vssd1 vccd1 vccd1 _7893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3987_ _3987_/A vssd1 vssd1 vccd1 vccd1 _8297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5726_ _5741_/S vssd1 vssd1 vccd1 vccd1 _5735_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5657_ _5552_/X _7803_/Q _5663_/S vssd1 vssd1 vccd1 vccd1 _5658_/A sky130_fd_sc_hd__mux2_1
X_4608_ _6801_/A vssd1 vssd1 vccd1 vccd1 _6910_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5588_ _7832_/Q _5587_/X _5588_/S vssd1 vssd1 vccd1 vccd1 _5589_/A sky130_fd_sc_hd__mux2_1
X_8376_ _8376_/CLK _8376_/D vssd1 vssd1 vccd1 vccd1 _8376_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3386_ _6938_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3386_/X sky130_fd_sc_hd__clkbuf_16
X_4539_ _8066_/Q vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__inv_2
XFILLER_7_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6470__250 _6470__250/A vssd1 vssd1 vccd1 vccd1 _7807_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7258_ _8230_/Q _7258_/B vssd1 vssd1 vccd1 vccd1 _7262_/D sky130_fd_sc_hd__nand2_1
XFILLER_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _6209_/A vssd1 vssd1 vccd1 vccd1 _6209_/X sky130_fd_sc_hd__buf_1
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3206_ clkbuf_0__3206_/X vssd1 vssd1 vccd1 vccd1 _6508__280/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7575__47 _7578__50/A vssd1 vssd1 vccd1 vccd1 _8386_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8443__218 vssd1 vssd1 vccd1 vccd1 _8443__218/HI manufacturerID[10] sky130_fd_sc_hd__conb_1
XFILLER_67_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7315__136 _7316__137/A vssd1 vssd1 vccd1 vccd1 _8263_/CLK sky130_fd_sc_hd__inv_2
X_6640__342 _6641__343/A vssd1 vssd1 vccd1 vccd1 _7923_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3910_ _3910_/A vssd1 vssd1 vccd1 vccd1 _8322_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3410_ clkbuf_0__3410_/X vssd1 vssd1 vccd1 vccd1 _7062__90/A sky130_fd_sc_hd__clkbuf_4
X_4890_ _4890_/A vssd1 vssd1 vccd1 vccd1 _8039_/D sky130_fd_sc_hd__clkbuf_1
X_3841_ _8382_/Q _3840_/X _3841_/S vssd1 vssd1 vccd1 vccd1 _3842_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6560_ _7863_/Q _5893_/A _6564_/S vssd1 vssd1 vccd1 vccd1 _6561_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3772_ _8365_/Q vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__buf_2
X_5511_ _5511_/A _5511_/B vssd1 vssd1 vccd1 vccd1 _5527_/S sky130_fd_sc_hd__nor2_2
XFILLER_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8230_ _8231_/CLK _8230_/D vssd1 vssd1 vccd1 vccd1 _8230_/Q sky130_fd_sc_hd__dfxtp_1
X_5442_ _5442_/A vssd1 vssd1 vccd1 vccd1 _7916_/D sky130_fd_sc_hd__clkbuf_1
X_5373_ _7949_/Q _4514_/X _5377_/S vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__mux2_1
X_8161_ _8161_/CLK _8161_/D vssd1 vssd1 vccd1 vccd1 _8161_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3240_ _6581_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3240_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7112_ _7237_/A _7134_/A _7125_/C _7119_/C vssd1 vssd1 vccd1 vccd1 _7238_/A sky130_fd_sc_hd__or4b_2
X_8092_ _8092_/CLK _8092_/D vssd1 vssd1 vccd1 vccd1 _8092_/Q sky130_fd_sc_hd__dfxtp_1
X_4324_ _4324_/A _4324_/B _4843_/A vssd1 vssd1 vccd1 vccd1 _5653_/B sky130_fd_sc_hd__or3b_4
X_4255_ _4255_/A vssd1 vssd1 vccd1 vccd1 _8177_/D sky130_fd_sc_hd__clkbuf_1
X_4186_ _4912_/A _5689_/B vssd1 vssd1 vccd1 vccd1 _4202_/S sky130_fd_sc_hd__nor2_2
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7945_ _7945_/CLK _7945_/D vssd1 vssd1 vccd1 vccd1 _7945_/Q sky130_fd_sc_hd__dfxtp_1
X_7876_ _7876_/CLK _7876_/D vssd1 vssd1 vccd1 vccd1 _7876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6758_ _8346_/Q _7416_/C _6757_/X vssd1 vssd1 vccd1 vccd1 _7491_/A sky130_fd_sc_hd__a21oi_2
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6689_ _8340_/Q _8339_/Q vssd1 vssd1 vccd1 vccd1 _6702_/A sky130_fd_sc_hd__and2_1
X_5709_ _7780_/Q _5573_/X _5717_/S vssd1 vssd1 vccd1 vccd1 _5710_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8359_ _8359_/CLK _8359_/D vssd1 vssd1 vccd1 vccd1 _8359_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__3369_ _6859_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3369_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4040_ _8274_/Q _3959_/X _4042_/S vssd1 vssd1 vccd1 vccd1 _4041_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5991_ _7718_/Q input31/X _5991_/S vssd1 vssd1 vccd1 vccd1 _5991_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7730_ _7991_/CLK _7730_/D vssd1 vssd1 vccd1 vccd1 _7730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _4942_/A vssd1 vssd1 vccd1 vccd1 _8017_/D sky130_fd_sc_hd__clkbuf_1
X_7661_ _6081_/A _7661_/D vssd1 vssd1 vccd1 vccd1 _7661_/Q sky130_fd_sc_hd__dfxtp_1
X_4873_ _6907_/C _4873_/B _4873_/C vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__and3_1
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7592_ _7602_/A vssd1 vssd1 vccd1 vccd1 _7599_/B sky130_fd_sc_hd__clkbuf_2
X_3824_ _3824_/A vssd1 vssd1 vccd1 vccd1 _8388_/D sky130_fd_sc_hd__clkbuf_1
X_6543_ _6543_/A vssd1 vssd1 vccd1 vccd1 _7855_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3255_ clkbuf_0__3255_/X vssd1 vssd1 vccd1 vccd1 _6655__354/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8213_ _8223_/CLK _8213_/D vssd1 vssd1 vccd1 vccd1 _8213_/Q sky130_fd_sc_hd__dfxtp_1
X_5425_ _7923_/Q _4511_/X _5431_/S vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__mux2_1
X_8144_ _8144_/CLK _8144_/D vssd1 vssd1 vccd1 vccd1 _8144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5356_ _3828_/X _7956_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5357_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_5 _5982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5287_ _7990_/Q vssd1 vssd1 vccd1 vccd1 _5555_/A sky130_fd_sc_hd__buf_2
X_4307_ _8154_/Q _4229_/X _4315_/S vssd1 vssd1 vccd1 vccd1 _4308_/A sky130_fd_sc_hd__mux2_1
X_6686__375 _6686__375/A vssd1 vssd1 vccd1 vccd1 _7959_/CLK sky130_fd_sc_hd__inv_2
X_8075_ _8075_/CLK _8075_/D vssd1 vssd1 vccd1 vccd1 _8075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4238_ _4238_/A vssd1 vssd1 vccd1 vccd1 _8184_/D sky130_fd_sc_hd__clkbuf_1
X_7026_ _7026_/A vssd1 vssd1 vccd1 vccd1 _7026_/X sky130_fd_sc_hd__buf_1
X_6647__348 _6647__348/A vssd1 vssd1 vccd1 vccd1 _7929_/CLK sky130_fd_sc_hd__inv_2
X_4169_ _8212_/Q _4044_/X _4177_/S vssd1 vssd1 vccd1 vccd1 _4170_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7928_ _7928_/CLK _7928_/D vssd1 vssd1 vccd1 vccd1 _7928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7859_ _8349_/CLK _7859_/D vssd1 vssd1 vccd1 vccd1 _7859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6483__260 _6483__260/A vssd1 vssd1 vccd1 vccd1 _7817_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7387__20 _7387__20/A vssd1 vssd1 vccd1 vccd1 _8322_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8449__224 vssd1 vssd1 vccd1 vccd1 _8449__224/HI partID[12] sky130_fd_sc_hd__conb_1
X_5210_ _5267_/A _5210_/B _5210_/C vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__or3_1
X_6190_ _6190_/A vssd1 vssd1 vccd1 vccd1 _7702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5141_ _5124_/A _5129_/X _5133_/X _5002_/A _5140_/X vssd1 vssd1 vccd1 vccd1 _5141_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5072_ _5002_/X _5059_/X _5063_/X _5071_/X vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__a31o_2
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6943__495 _6943__495/A vssd1 vssd1 vccd1 vccd1 _8092_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4023_ _4023_/A vssd1 vssd1 vccd1 vccd1 _8282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _7546_/A vssd1 vssd1 vccd1 vccd1 _6400_/A sky130_fd_sc_hd__buf_4
X_7713_ _7989_/CLK _7713_/D vssd1 vssd1 vccd1 vccd1 _7713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4925_ _4925_/A vssd1 vssd1 vccd1 vccd1 _8024_/D sky130_fd_sc_hd__clkbuf_1
X_7644_ _8397_/CLK _7644_/D vssd1 vssd1 vccd1 vccd1 _7644_/Q sky130_fd_sc_hd__dfxtp_1
X_4856_ _4856_/A vssd1 vssd1 vccd1 vccd1 _8053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3807_ _7733_/Q _6341_/A _6342_/B _7732_/Q vssd1 vssd1 vccd1 vccd1 _3812_/A sky130_fd_sc_hd__or4b_1
X_6526_ _7605_/B _7848_/Q _6528_/S vssd1 vssd1 vccd1 vccd1 _6527_/A sky130_fd_sc_hd__mux2_1
X_4787_ _7790_/Q _4676_/A _4786_/X _4729_/X vssd1 vssd1 vccd1 vccd1 _4787_/X sky130_fd_sc_hd__o22a_1
X_6653__352 _6655__354/A vssd1 vssd1 vccd1 vccd1 _7933_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6388_ _6388_/A vssd1 vssd1 vccd1 vccd1 _7748_/D sky130_fd_sc_hd__clkbuf_1
X_5408_ _5408_/A vssd1 vssd1 vccd1 vccd1 _7931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3206_ _6503_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3206_/X sky130_fd_sc_hd__clkbuf_16
X_5339_ _5296_/X _7964_/Q _5339_/S vssd1 vssd1 vccd1 vccd1 _5340_/A sky130_fd_sc_hd__mux2_1
X_8127_ _8127_/CLK _8127_/D vssd1 vssd1 vccd1 vccd1 _8127_/Q sky130_fd_sc_hd__dfxtp_1
X_8058_ _8058_/CLK _8058_/D vssd1 vssd1 vccd1 vccd1 _8058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3385_ clkbuf_0__3385_/X vssd1 vssd1 vccd1 vccd1 _6936__489/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6596__306 _6597__307/A vssd1 vssd1 vccd1 vccd1 _7887_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4716_/A _7888_/Q _7832_/Q _4717_/A vssd1 vssd1 vccd1 vccd1 _4710_/X sky130_fd_sc_hd__a22o_1
X_5690_ _5705_/S vssd1 vssd1 vccd1 vccd1 _5699_/S sky130_fd_sc_hd__buf_2
XFILLER_15_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4641_ _4641_/A vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4572_ _8021_/Q _7876_/Q _7780_/Q _7764_/Q _4569_/X _4571_/X vssd1 vssd1 vccd1 vccd1
+ _4572_/X sky130_fd_sc_hd__mux4_1
X_6311_ _6332_/C vssd1 vssd1 vccd1 vccd1 _6322_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6242_ _6237_/A _6241_/Y _6254_/B vssd1 vssd1 vccd1 vccd1 _6289_/B sky130_fd_sc_hd__o21a_1
XFILLER_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6173_ _6173_/A vssd1 vssd1 vccd1 vccd1 _7696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5124_ _5124_/A _5124_/B vssd1 vssd1 vccd1 vccd1 _5124_/X sky130_fd_sc_hd__or2_1
X_5055_ _3872_/X _5029_/X _5054_/X _5027_/X vssd1 vssd1 vccd1 vccd1 _8010_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4006_ _4006_/A vssd1 vssd1 vccd1 vccd1 _8289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6991__533 _6991__533/A vssd1 vssd1 vccd1 vccd1 _8130_/CLK sky130_fd_sc_hd__inv_2
X_5957_ _5957_/A vssd1 vssd1 vccd1 vccd1 _5957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4908_ _8031_/Q _4407_/X _4910_/S vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__mux2_1
X_5888_ _5888_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__or2_1
X_7627_ _8402_/Q _7627_/B vssd1 vssd1 vccd1 vccd1 _7627_/Y sky130_fd_sc_hd__nor2_1
X_4839_ _8056_/Q _4604_/A _4836_/X _4838_/Y vssd1 vssd1 vccd1 vccd1 _8056_/D sky130_fd_sc_hd__o211a_1
X_7381__15 _7381__15/A vssd1 vssd1 vccd1 vccd1 _8317_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7489_ _7489_/A vssd1 vssd1 vccd1 vccd1 _7527_/B sky130_fd_sc_hd__clkbuf_2
X_6509_ _6575_/A vssd1 vssd1 vccd1 vccd1 _6509_/X sky130_fd_sc_hd__buf_1
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7079__103 _7080__104/A vssd1 vssd1 vccd1 vccd1 _8200_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6584__298 _6586__300/A vssd1 vssd1 vccd1 vccd1 _7879_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3368_ clkbuf_0__3368_/X vssd1 vssd1 vccd1 vccd1 _6857__429/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6604__313 _6606__315/A vssd1 vssd1 vccd1 vccd1 _7894_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5811_ _4099_/X _7645_/Q _5811_/S vssd1 vssd1 vccd1 vccd1 _5812_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5742_ _5742_/A vssd1 vssd1 vccd1 vccd1 _7765_/D sky130_fd_sc_hd__clkbuf_1
X_5673_ _7796_/Q _5573_/X _5681_/S vssd1 vssd1 vccd1 vccd1 _5674_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4624_ _7651_/Q _7659_/Q _7710_/Q _7811_/Q _4595_/X _4596_/X vssd1 vssd1 vccd1 vccd1
+ _4624_/X sky130_fd_sc_hd__mux4_2
X_7412_ _7612_/A _7412_/B vssd1 vssd1 vccd1 vccd1 _7412_/X sky130_fd_sc_hd__xor2_1
X_8392_ _8399_/CLK _8392_/D vssd1 vssd1 vccd1 vccd1 _8392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4555_ _4641_/A vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__clkbuf_4
X_7274_ _8006_/Q _7266_/X _7273_/X _7269_/X vssd1 vssd1 vccd1 vccd1 _8234_/D sky130_fd_sc_hd__o211a_1
X_4486_ _4347_/X _8083_/Q _4486_/S vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6225_ _7732_/Q _6909_/A _6342_/B vssd1 vssd1 vccd1 vccd1 _6226_/C sky130_fd_sc_hd__or3_2
X_6156_ _7863_/Q _6151_/X _6152_/X _6154_/X _7687_/Q vssd1 vssd1 vccd1 vccd1 _7687_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5151_/A vssd1 vssd1 vccd1 vccd1 _5108_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5038_ _5204_/S vssd1 vssd1 vccd1 vccd1 _5207_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6505__277 _6507__279/A vssd1 vssd1 vccd1 vccd1 _7834_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput98 _5937_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998__539 _6998__539/A vssd1 vssd1 vccd1 vccd1 _8136_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7050__80 _7050__80/A vssd1 vssd1 vccd1 vccd1 _8177_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4340_ _4340_/A vssd1 vssd1 vccd1 vccd1 _8142_/D sky130_fd_sc_hd__clkbuf_1
X_4271_ _4271_/A vssd1 vssd1 vccd1 vccd1 _8170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _7672_/Q _6008_/X _6023_/S vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__mux2_4
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7961_ _7961_/CLK _7961_/D vssd1 vssd1 vccd1 vccd1 _7961_/Q sky130_fd_sc_hd__dfxtp_1
X_7892_ _7892_/CLK _7892_/D vssd1 vssd1 vccd1 vccd1 _7892_/Q sky130_fd_sc_hd__dfxtp_1
X_6774_ _6786_/A vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__buf_1
X_3986_ _8297_/Q _3963_/X _3986_/S vssd1 vssd1 vccd1 vccd1 _3987_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5725_ _5725_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _5741_/S sky130_fd_sc_hd__nor2_2
XFILLER_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _5656_/A vssd1 vssd1 vccd1 vccd1 _7804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4607_ _4844_/A vssd1 vssd1 vccd1 vccd1 _6801_/A sky130_fd_sc_hd__buf_2
XFILLER_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5587_ _7988_/Q vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__clkbuf_2
X_8375_ _8375_/CLK _8375_/D vssd1 vssd1 vccd1 vccd1 _8375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4538_ _4538_/A vssd1 vssd1 vccd1 vccd1 _4538_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__3385_ _6932_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3385_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7326_ _7326_/A vssd1 vssd1 vccd1 vccd1 _7326_/X sky130_fd_sc_hd__buf_1
XFILLER_117_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7257_ _7257_/A vssd1 vssd1 vccd1 vccd1 _8229_/D sky130_fd_sc_hd__clkbuf_1
X_4469_ _4469_/A vssd1 vssd1 vccd1 vccd1 _8091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6139_ _6136_/X _7853_/Q _6134_/X _6137_/X _7677_/Q vssd1 vssd1 vccd1 vccd1 _7677_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_100_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3205_ clkbuf_0__3205_/X vssd1 vssd1 vccd1 vccd1 _6575_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3840_ _8358_/Q vssd1 vssd1 vccd1 vccd1 _3840_/X sky130_fd_sc_hd__buf_2
X_5510_ _5510_/A vssd1 vssd1 vccd1 vccd1 _7885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6490_ _6496_/A vssd1 vssd1 vccd1 vccd1 _6490_/X sky130_fd_sc_hd__buf_1
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5441_ _3772_/X _7916_/Q _5449_/S vssd1 vssd1 vccd1 vccd1 _5442_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5372_ _5372_/A vssd1 vssd1 vccd1 vccd1 _7950_/D sky130_fd_sc_hd__clkbuf_1
X_8160_ _8160_/CLK _8160_/D vssd1 vssd1 vccd1 vccd1 _8160_/Q sky130_fd_sc_hd__dfxtp_1
X_4323_ _7992_/Q vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__clkbuf_2
X_7111_ _8222_/Q _8221_/Q vssd1 vssd1 vccd1 vccd1 _7119_/C sky130_fd_sc_hd__and2_1
X_8091_ _8091_/CLK _8091_/D vssd1 vssd1 vccd1 vccd1 _8091_/Q sky130_fd_sc_hd__dfxtp_1
X_6866__436 _6868__438/A vssd1 vssd1 vccd1 vccd1 _8031_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4254_ _4208_/X _8177_/Q _4260_/S vssd1 vssd1 vccd1 vccd1 _4255_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4185_ _4414_/A _4413_/A _4387_/B vssd1 vssd1 vccd1 vccd1 _5689_/B sky130_fd_sc_hd__or3b_4
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7944_ _7944_/CLK _7944_/D vssd1 vssd1 vccd1 vccd1 _7944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ _7875_/CLK _7875_/D vssd1 vssd1 vccd1 vccd1 _7875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6757_ _8346_/Q _8345_/Q _8344_/Q _6757_/D vssd1 vssd1 vccd1 vccd1 _6757_/X sky130_fd_sc_hd__and4b_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5708_ _5723_/S vssd1 vssd1 vccd1 vccd1 _5717_/S sky130_fd_sc_hd__buf_2
X_3969_ _5475_/A vssd1 vssd1 vccd1 vccd1 _5367_/B sky130_fd_sc_hd__buf_4
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6688_ _3814_/X _6287_/X _7531_/C _6118_/A vssd1 vssd1 vccd1 vccd1 _7519_/A sky130_fd_sc_hd__a31oi_4
X_5639_ _7811_/Q _5578_/X _5645_/S vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__mux2_1
X_8358_ _8359_/CLK _8358_/D vssd1 vssd1 vccd1 vccd1 _8358_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3368_ _6853_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3368_/X sky130_fd_sc_hd__clkbuf_16
X_8289_ _8289_/CLK _8289_/D vssd1 vssd1 vccd1 vccd1 _8289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7321__141 _7322__142/A vssd1 vssd1 vccd1 vccd1 _8268_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5990_ _5990_/A vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__clkbuf_1
X_4941_ _4338_/X _8017_/Q _4941_/S vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__mux2_1
X_7660_ _7660_/CLK _7660_/D vssd1 vssd1 vccd1 vccd1 _7660_/Q sky130_fd_sc_hd__dfxtp_1
X_4872_ _4872_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4873_/C sky130_fd_sc_hd__nand2_1
X_3823_ _8388_/Q _3822_/X _3832_/S vssd1 vssd1 vccd1 vccd1 _3824_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7591_ _7595_/A _7591_/B vssd1 vssd1 vccd1 vccd1 _7591_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6542_ _5875_/A _7855_/Q _6546_/S vssd1 vssd1 vccd1 vccd1 _6543_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_9_wb_clk_i _7717_/CLK vssd1 vssd1 vccd1 vccd1 _7747_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1_0__3254_ clkbuf_0__3254_/X vssd1 vssd1 vccd1 vccd1 _6675_/A sky130_fd_sc_hd__clkbuf_4
X_8212_ _8212_/CLK _8212_/D vssd1 vssd1 vccd1 vccd1 _8212_/Q sky130_fd_sc_hd__dfxtp_1
X_5424_ _5424_/A vssd1 vssd1 vccd1 vccd1 _7924_/D sky130_fd_sc_hd__clkbuf_1
X_8143_ _8143_/CLK _8143_/D vssd1 vssd1 vccd1 vccd1 _8143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5355_ _5355_/A vssd1 vssd1 vccd1 vccd1 _7957_/D sky130_fd_sc_hd__clkbuf_1
X_5286_ _5286_/A vssd1 vssd1 vccd1 vccd1 _7983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_6 _5982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8074_ _8074_/CLK _8074_/D vssd1 vssd1 vccd1 vccd1 _8074_/Q sky130_fd_sc_hd__dfxtp_1
X_4306_ _4321_/S vssd1 vssd1 vccd1 vccd1 _4315_/S sky130_fd_sc_hd__buf_2
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4237_ _8184_/Q _4128_/X _4241_/S vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4168_ _4183_/S vssd1 vssd1 vccd1 vccd1 _4177_/S sky130_fd_sc_hd__clkbuf_4
X_4099_ _7985_/Q vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__buf_2
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7927_ _7927_/CLK _7927_/D vssd1 vssd1 vccd1 vccd1 _7927_/Q sky130_fd_sc_hd__dfxtp_1
X_6955__504 _6955__504/A vssd1 vssd1 vccd1 vccd1 _8101_/CLK sky130_fd_sc_hd__inv_2
X_7858_ _8349_/CLK _7858_/D vssd1 vssd1 vccd1 vccd1 _7858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6809_ _6809_/A vssd1 vssd1 vccd1 vccd1 _7990_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7789_ _7789_/CLK _7789_/D vssd1 vssd1 vccd1 vccd1 _7789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3599_ clkbuf_0__3599_/X vssd1 vssd1 vccd1 vccd1 _7379__13/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _5243_/A _5140_/B _5140_/C vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__or3_1
X_5071_ _5065_/X _5067_/X _5070_/X _5019_/X _5095_/A vssd1 vssd1 vccd1 vccd1 _5071_/X
+ sky130_fd_sc_hd__o221a_1
X_4022_ _3887_/X _8282_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5973_ _7713_/Q input14/X _6052_/A vssd1 vssd1 vccd1 vccd1 _5973_/X sky130_fd_sc_hd__mux2_4
XFILLER_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7712_ _7989_/CLK _7712_/D vssd1 vssd1 vccd1 vccd1 _7712_/Q sky130_fd_sc_hd__dfxtp_1
X_4924_ _8024_/Q _4404_/X _4928_/S vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7643_ _7643_/A vssd1 vssd1 vccd1 vccd1 _8407_/D sky130_fd_sc_hd__clkbuf_1
X_4855_ _6907_/C _4855_/B _4855_/C vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__and3_1
X_3806_ _7740_/Q _7741_/Q vssd1 vssd1 vccd1 vccd1 _6342_/B sky130_fd_sc_hd__or2_1
X_4786_ _4730_/X _7886_/Q _7830_/Q _4698_/A vssd1 vssd1 vccd1 vccd1 _4786_/X sky130_fd_sc_hd__a22o_1
X_6525_ _6525_/A vssd1 vssd1 vccd1 vccd1 _7847_/D sky130_fd_sc_hd__clkbuf_1
X_7328__147 _7329__148/A vssd1 vssd1 vccd1 vccd1 _8274_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6387_ _7855_/Q _7748_/Q _6393_/S vssd1 vssd1 vccd1 vccd1 _6388_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5407_ _7931_/Q _4511_/X _5413_/S vssd1 vssd1 vccd1 vccd1 _5408_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5338_ _5338_/A vssd1 vssd1 vccd1 vccd1 _7965_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3205_ _6502_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3205_/X sky130_fd_sc_hd__clkbuf_16
X_8126_ _8126_/CLK _8126_/D vssd1 vssd1 vccd1 vccd1 _8126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8057_ _8057_/CLK _8057_/D vssd1 vssd1 vccd1 vccd1 _8057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5269_ _5269_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3384_ clkbuf_0__3384_/X vssd1 vssd1 vccd1 vccd1 _6928__482/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8409__231 vssd1 vssd1 vccd1 vccd1 partID[0] _8409__231/LO sky130_fd_sc_hd__conb_1
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4557_/A _4637_/X _4639_/X vssd1 vssd1 vccd1 vccd1 _4640_/X sky130_fd_sc_hd__a21o_1
X_6310_ _6337_/B vssd1 vssd1 vccd1 vccd1 _6326_/B sky130_fd_sc_hd__clkbuf_1
X_4571_ _4571_/A vssd1 vssd1 vccd1 vccd1 _4571_/X sky130_fd_sc_hd__buf_2
XFILLER_115_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6241_ _7734_/Q _6350_/C _6343_/B _6241_/D vssd1 vssd1 vccd1 vccd1 _6241_/Y sky130_fd_sc_hd__nand4_1
X_6172_ _7538_/B _7696_/Q _6174_/S vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__mux2_1
X_5123_ _5121_/X _5122_/X _5123_/S vssd1 vssd1 vccd1 vccd1 _5124_/B sky130_fd_sc_hd__mux2_2
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _8010_/Q _4955_/X _5031_/X _5053_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _5054_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4005_ _8289_/Q _3963_/X _4005_/S vssd1 vssd1 vccd1 vccd1 _4006_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7334__151 _7336__153/A vssd1 vssd1 vccd1 vccd1 _8278_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5956_ _7860_/Q _5964_/B vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__and2_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5887_ _5887_/A vssd1 vssd1 vccd1 vccd1 _5887_/X sky130_fd_sc_hd__clkbuf_1
X_4907_ _4907_/A vssd1 vssd1 vccd1 vccd1 _8032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7626_ _7626_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7626_/Y sky130_fd_sc_hd__nand2_1
X_4838_ _4853_/B vssd1 vssd1 vccd1 vccd1 _4838_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4769_ _7971_/Q _4681_/A _4642_/A _4768_/X vssd1 vssd1 vccd1 vccd1 _4770_/C sky130_fd_sc_hd__o211a_1
XFILLER_119_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7488_ _7488_/A _7488_/B vssd1 vssd1 vccd1 vccd1 _8345_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8109_ _8109_/CLK _8109_/D vssd1 vssd1 vccd1 vccd1 _8109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3367_ clkbuf_0__3367_/X vssd1 vssd1 vccd1 vccd1 _6871_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7366__2 _7366__2/A vssd1 vssd1 vccd1 vccd1 _8304_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8334_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5810_ _5810_/A vssd1 vssd1 vccd1 vccd1 _7646_/D sky130_fd_sc_hd__clkbuf_1
X_5741_ _7765_/Q _5570_/A _5741_/S vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__mux2_1
X_7411_ _7411_/A _7411_/B vssd1 vssd1 vccd1 vccd1 _7412_/B sky130_fd_sc_hd__nand2_1
X_6793__396 _6796__399/A vssd1 vssd1 vccd1 vccd1 _7981_/CLK sky130_fd_sc_hd__inv_2
X_5672_ _5687_/S vssd1 vssd1 vccd1 vccd1 _5681_/S sky130_fd_sc_hd__clkbuf_4
X_4623_ _4619_/X _4620_/X _4650_/S vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__mux2_1
X_8391_ _8391_/CLK _8391_/D vssd1 vssd1 vccd1 vccd1 _8391_/Q sky130_fd_sc_hd__dfxtp_1
X_4554_ _4573_/B _4675_/A vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__or2_1
X_7273_ _8234_/Q _7277_/B vssd1 vssd1 vccd1 vccd1 _7273_/X sky130_fd_sc_hd__or2_1
XFILLER_104_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6224_ _7733_/Q vssd1 vssd1 vccd1 vccd1 _6909_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4485_ _4485_/A vssd1 vssd1 vccd1 vccd1 _8084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6155_ _7862_/Q _6151_/X _6152_/X _6154_/X _7686_/Q vssd1 vssd1 vccd1 vccd1 _7686_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_106_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5115_/A vssd1 vssd1 vccd1 vccd1 _5151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _7000_/A vssd1 vssd1 vccd1 vccd1 _6988_/X sky130_fd_sc_hd__buf_1
X_5939_ _5939_/A vssd1 vssd1 vccd1 vccd1 _5939_/X sky130_fd_sc_hd__clkbuf_1
X_7609_ _6754_/A _7608_/Y _7615_/B vssd1 vssd1 vccd1 vccd1 _7610_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3599_ _7376_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3599_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput99 _5939_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__buf_2
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6820__404 _6820__404/A vssd1 vssd1 vccd1 vccd1 _7997_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _8170_/Q _4229_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7960_ _8364_/CLK _7960_/D vssd1 vssd1 vccd1 vccd1 _7960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7891_ _7891_/CLK _7891_/D vssd1 vssd1 vccd1 vccd1 _7891_/Q sky130_fd_sc_hd__dfxtp_1
X_6911_ _6911_/A vssd1 vssd1 vccd1 vccd1 _8066_/D sky130_fd_sc_hd__clkbuf_1
X_6842_ _6842_/A vssd1 vssd1 vccd1 vccd1 _8013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _3985_/A vssd1 vssd1 vccd1 vccd1 _8298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5724_ _5724_/A vssd1 vssd1 vccd1 vccd1 _7773_/D sky130_fd_sc_hd__clkbuf_1
X_5655_ _5547_/X _7804_/Q _5663_/S vssd1 vssd1 vccd1 vccd1 _5656_/A sky130_fd_sc_hd__mux2_1
X_4606_ _4540_/X _8064_/Q _4869_/A _4603_/X _4605_/X vssd1 vssd1 vccd1 vccd1 _4606_/X
+ sky130_fd_sc_hd__a221o_1
X_8374_ _8374_/CLK _8374_/D vssd1 vssd1 vccd1 vccd1 _8374_/Q sky130_fd_sc_hd__dfxtp_1
X_5586_ _5586_/A vssd1 vssd1 vccd1 vccd1 _7833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3384_ _6926_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3384_/X sky130_fd_sc_hd__clkbuf_16
X_4537_ _4604_/A _4604_/B _4604_/C vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__nand3_2
X_7256_ _7254_/X _7285_/S _7256_/C vssd1 vssd1 vccd1 vccd1 _7257_/A sky130_fd_sc_hd__and3b_1
X_4468_ _3840_/X _8091_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4469_/A sky130_fd_sc_hd__mux2_1
X_7187_ _7187_/A vssd1 vssd1 vccd1 vccd1 _7187_/X sky130_fd_sc_hd__buf_1
X_6138_ _6136_/X _7852_/Q _6134_/X _6137_/X _7676_/Q vssd1 vssd1 vccd1 vccd1 _7676_/D
+ sky130_fd_sc_hd__o32a_1
X_4399_ _8119_/Q _4398_/X _4402_/S vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__mux2_1
X_6511__282 _6511__282/A vssd1 vssd1 vccd1 vccd1 _7839_/CLK sky130_fd_sc_hd__inv_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _7691_/Q _6061_/X _6039_/A _6068_/X vssd1 vssd1 vccd1 vccd1 _6069_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3204_ clkbuf_0__3204_/X vssd1 vssd1 vccd1 vccd1 _6500__274/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7024__59 _7025__60/A vssd1 vssd1 vccd1 vccd1 _8156_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _5455_/S vssd1 vssd1 vccd1 vccd1 _5449_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6454__236 _6458__240/A vssd1 vssd1 vccd1 vccd1 _7793_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5371_ _7950_/Q _4511_/X _5377_/S vssd1 vssd1 vccd1 vccd1 _5372_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8090_ _8090_/CLK _8090_/D vssd1 vssd1 vccd1 vccd1 _8090_/Q sky130_fd_sc_hd__dfxtp_1
X_7110_ _8220_/Q _8219_/Q _7110_/C _7129_/A vssd1 vssd1 vccd1 vccd1 _7125_/C sky130_fd_sc_hd__nand4_1
X_4322_ _4322_/A vssd1 vssd1 vccd1 vccd1 _8147_/D sky130_fd_sc_hd__clkbuf_1
X_4253_ _4253_/A vssd1 vssd1 vccd1 vccd1 _8178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4184_ _4184_/A vssd1 vssd1 vccd1 vccd1 _8205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7943_ _8391_/CLK _7943_/D vssd1 vssd1 vccd1 vccd1 _7943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7874_ _7874_/CLK _7874_/D vssd1 vssd1 vccd1 vccd1 _7874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6756_ _6747_/X _6749_/Y _6751_/Y _6754_/Y _6755_/X vssd1 vssd1 vccd1 vccd1 _6763_/B
+ sky130_fd_sc_hd__o2111a_1
X_3968_ _5261_/A _3968_/B _6838_/A _3867_/A vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__or4bb_4
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5707_ _5725_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5723_/S sky130_fd_sc_hd__nor2_2
X_6687_ _6687_/A _6687_/B _7546_/C vssd1 vssd1 vccd1 vccd1 _7531_/C sky130_fd_sc_hd__and3_2
X_3899_ _3872_/X _8327_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3900_/A sky130_fd_sc_hd__mux2_1
X_6617__324 _6618__325/A vssd1 vssd1 vccd1 vccd1 _7905_/CLK sky130_fd_sc_hd__inv_2
X_5638_ _5638_/A vssd1 vssd1 vccd1 vccd1 _7812_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3399_ clkbuf_0__3399_/X vssd1 vssd1 vccd1 vccd1 _7010__549/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8357_ _8399_/CLK _8357_/D vssd1 vssd1 vccd1 vccd1 _8357_/Q sky130_fd_sc_hd__dfxtp_1
X_5569_ _5569_/A vssd1 vssd1 vccd1 vccd1 _7838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3367_ _6852_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3367_/X sky130_fd_sc_hd__clkbuf_16
X_7308_ _7326_/A vssd1 vssd1 vccd1 vccd1 _7308_/X sky130_fd_sc_hd__buf_1
X_8288_ _8288_/CLK _8288_/D vssd1 vssd1 vccd1 vccd1 _8288_/Q sky130_fd_sc_hd__dfxtp_1
X_7239_ _7237_/X _7238_/Y _7251_/A vssd1 vssd1 vccd1 vccd1 _8223_/D sky130_fd_sc_hd__a21oi_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _4940_/A vssd1 vssd1 vccd1 vccd1 _8018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4871_ _4872_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4873_/B sky130_fd_sc_hd__or2_1
X_6872__441 _6873__442/A vssd1 vssd1 vccd1 vccd1 _8036_/CLK sky130_fd_sc_hd__inv_2
X_7590_ _7615_/B vssd1 vssd1 vccd1 vccd1 _7590_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3822_ _8364_/Q vssd1 vssd1 vccd1 vccd1 _3822_/X sky130_fd_sc_hd__buf_2
X_6541_ _6541_/A vssd1 vssd1 vccd1 vccd1 _7854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6472_ _6478_/A vssd1 vssd1 vccd1 vccd1 _6472_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3253_ clkbuf_0__3253_/X vssd1 vssd1 vccd1 vccd1 _6647__348/A sky130_fd_sc_hd__clkbuf_4
X_8211_ _8211_/CLK _8211_/D vssd1 vssd1 vccd1 vccd1 _8211_/Q sky130_fd_sc_hd__dfxtp_1
X_5423_ _7924_/Q _5366_/X _5431_/S vssd1 vssd1 vccd1 vccd1 _5424_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5354_ _3825_/X _7957_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__mux2_1
X_8142_ _8142_/CLK _8142_/D vssd1 vssd1 vccd1 vccd1 _8142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _5385_/A _4368_/B vssd1 vssd1 vccd1 vccd1 _4321_/S sky130_fd_sc_hd__nor2_4
X_5285_ _5284_/X _7983_/Q _5297_/S vssd1 vssd1 vccd1 vccd1 _5286_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_7 _7285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8073_ _8073_/CLK _8073_/D vssd1 vssd1 vccd1 vccd1 _8073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _4236_/A vssd1 vssd1 vccd1 vccd1 _8185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4167_ _5635_/A _5548_/A vssd1 vssd1 vccd1 vccd1 _4183_/S sky130_fd_sc_hd__nor2_2
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4098_ _4098_/A vssd1 vssd1 vccd1 vccd1 _8266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7926_ _7926_/CLK _7926_/D vssd1 vssd1 vccd1 vccd1 _7926_/Q sky130_fd_sc_hd__dfxtp_1
X_7857_ _8348_/CLK _7857_/D vssd1 vssd1 vccd1 vccd1 _7857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6808_ _8355_/Q _6810_/B vssd1 vssd1 vccd1 vccd1 _6809_/A sky130_fd_sc_hd__and2_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7788_ _7788_/CLK _7788_/D vssd1 vssd1 vccd1 vccd1 _7788_/Q sky130_fd_sc_hd__dfxtp_1
X_8433__208 vssd1 vssd1 vccd1 vccd1 _8433__208/HI manufacturerID[0] sky130_fd_sc_hd__conb_1
XFILLER_109_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6739_ _8403_/Q _7432_/B vssd1 vssd1 vccd1 vccd1 _6739_/X sky130_fd_sc_hd__xor2_1
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3598_ clkbuf_0__3598_/X vssd1 vssd1 vccd1 vccd1 _7374__9/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5070_ _5068_/X _5069_/X _5089_/S vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__mux2_2
X_4021_ _4021_/A vssd1 vssd1 vccd1 vccd1 _8283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _5972_/A vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__clkbuf_1
X_7711_ _7711_/CLK _7711_/D vssd1 vssd1 vccd1 vccd1 _7711_/Q sky130_fd_sc_hd__dfxtp_1
X_4923_ _4923_/A vssd1 vssd1 vccd1 vccd1 _8025_/D sky130_fd_sc_hd__clkbuf_1
X_7642_ _7642_/A _7642_/B vssd1 vssd1 vccd1 vccd1 _7643_/A sky130_fd_sc_hd__or2_1
X_4854_ _4930_/C _4854_/B vssd1 vssd1 vccd1 vccd1 _4855_/C sky130_fd_sc_hd__or2_1
X_7393__25 _7393__25/A vssd1 vssd1 vccd1 vccd1 _8327_/CLK sky130_fd_sc_hd__inv_2
X_3805_ _7755_/Q _7754_/Q vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__nor2_2
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4785_ _4750_/X _4783_/X _4784_/X vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__o21a_1
X_7573_ _7573_/A vssd1 vssd1 vccd1 vccd1 _7573_/X sky130_fd_sc_hd__buf_1
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6524_ _7608_/B _7847_/Q _6528_/S vssd1 vssd1 vccd1 vccd1 _6525_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6386_ _6386_/A vssd1 vssd1 vccd1 vccd1 _7747_/D sky130_fd_sc_hd__clkbuf_1
X_5406_ _5406_/A vssd1 vssd1 vccd1 vccd1 _7932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5337_ _5292_/X _7965_/Q _5339_/S vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3204_ _6496_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3204_/X sky130_fd_sc_hd__clkbuf_16
X_8125_ _8125_/CLK _8125_/D vssd1 vssd1 vccd1 vccd1 _8125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5268_ _7996_/Q _5265_/A _5267_/Y _5178_/X vssd1 vssd1 vccd1 vccd1 _7996_/D sky130_fd_sc_hd__o211a_1
X_8056_ _8056_/CLK _8056_/D vssd1 vssd1 vccd1 vccd1 _8056_/Q sky130_fd_sc_hd__dfxtp_1
X_4219_ _4219_/A vssd1 vssd1 vccd1 vccd1 _8190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5199_ _8282_/Q _5098_/X _5183_/X _8274_/Q vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__o22a_1
X_6879__447 _6879__447/A vssd1 vssd1 vccd1 vccd1 _8042_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3383_ clkbuf_0__3383_/X vssd1 vssd1 vccd1 vccd1 _6925__480/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6660__358 _6661__359/A vssd1 vssd1 vccd1 vccd1 _7939_/CLK sky130_fd_sc_hd__inv_2
X_7909_ _7909_/CLK _7909_/D vssd1 vssd1 vccd1 vccd1 _7909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6411__201 _6413__203/A vssd1 vssd1 vccd1 vccd1 _7758_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _4682_/A vssd1 vssd1 vccd1 vccd1 _4571_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6240_ _6232_/Y _6235_/X _6254_/B vssd1 vssd1 vccd1 vccd1 _6240_/Y sky130_fd_sc_hd__o21ai_1
X_6171_ _6171_/A vssd1 vssd1 vccd1 vccd1 _7695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5122_ _8150_/Q _8134_/Q _8126_/Q _8158_/Q _5043_/A _5037_/X vssd1 vssd1 vccd1 vccd1
+ _5122_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5053_ _5002_/X _5035_/X _5041_/X _5052_/X vssd1 vssd1 vccd1 vccd1 _5053_/X sky130_fd_sc_hd__a31o_2
X_4004_ _4004_/A vssd1 vssd1 vccd1 vccd1 _8290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5955_ _5955_/A vssd1 vssd1 vccd1 vccd1 _5964_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5886_ _5886_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__or2_1
X_4906_ _8032_/Q _4404_/X _4910_/S vssd1 vssd1 vccd1 vccd1 _4907_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7625_ _7625_/A vssd1 vssd1 vccd1 vccd1 _8401_/D sky130_fd_sc_hd__clkbuf_1
X_4837_ _4843_/C vssd1 vssd1 vccd1 vccd1 _4853_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4768_ _8032_/Q _4676_/A _4767_/X _4750_/A vssd1 vssd1 vccd1 vccd1 _4768_/X sky130_fd_sc_hd__o22a_1
X_7487_ _7416_/B _7416_/C _7446_/Y _7458_/X _8345_/Q vssd1 vssd1 vccd1 vccd1 _7488_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4699_ _4699_/A vssd1 vssd1 vccd1 vccd1 _4699_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6885__451 _6889__455/A vssd1 vssd1 vccd1 vccd1 _8046_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6369_ _5927_/A _7740_/Q _6371_/S vssd1 vssd1 vccd1 vccd1 _6370_/A sky130_fd_sc_hd__mux2_1
X_8108_ _8108_/CLK _8108_/D vssd1 vssd1 vccd1 vccd1 _8108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8039_ _8039_/CLK _8039_/D vssd1 vssd1 vccd1 vccd1 _8039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8439__214 vssd1 vssd1 vccd1 vccd1 _8439__214/HI manufacturerID[6] sky130_fd_sc_hd__conb_1
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3366_ clkbuf_0__3366_/X vssd1 vssd1 vccd1 vccd1 _6981_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7062__90 _7062__90/A vssd1 vssd1 vccd1 vccd1 _8187_/CLK sky130_fd_sc_hd__inv_2
X_6968__515 _6968__515/A vssd1 vssd1 vccd1 vccd1 _8112_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5740_ _5740_/A vssd1 vssd1 vccd1 vccd1 _7766_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7410_ _7410_/A _7410_/B _7410_/C _7410_/D vssd1 vssd1 vccd1 vccd1 _7496_/B sky130_fd_sc_hd__and4_1
X_5671_ _5743_/A _5671_/B vssd1 vssd1 vccd1 vccd1 _5687_/S sky130_fd_sc_hd__nor2_2
X_8390_ _8397_/CLK _8390_/D vssd1 vssd1 vccd1 vccd1 _8390_/Q sky130_fd_sc_hd__dfxtp_1
X_6418__207 _6418__207/A vssd1 vssd1 vccd1 vccd1 _7764_/CLK sky130_fd_sc_hd__inv_2
X_4622_ _4622_/A vssd1 vssd1 vccd1 vccd1 _4650_/S sky130_fd_sc_hd__clkbuf_2
X_4553_ _4682_/A _4682_/B _8048_/Q vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__a21oi_1
XFILLER_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7272_ _8005_/Q _7266_/X _7271_/X _7269_/X vssd1 vssd1 vccd1 vccd1 _8233_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6611__319 _6611__319/A vssd1 vssd1 vccd1 vccd1 _7900_/CLK sky130_fd_sc_hd__inv_2
X_4484_ _4344_/X _8084_/Q _4486_/S vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__mux2_1
X_6223_ _7618_/A vssd1 vssd1 vccd1 vccd1 _6839_/C sky130_fd_sc_hd__buf_2
X_6154_ _6154_/A vssd1 vssd1 vccd1 vccd1 _6154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _8324_/Q _8070_/Q _5224_/S vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__mux2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _7939_/Q _7931_/Q _7923_/Q _7958_/Q _4978_/X _4995_/X vssd1 vssd1 vccd1 vccd1
+ _5036_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5938_ _7852_/Q _5942_/B vssd1 vssd1 vccd1 vccd1 _5939_/A sky130_fd_sc_hd__and2_1
XFILLER_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5869_ _7591_/B _5877_/B vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__or2_1
XFILLER_21_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7608_ _7608_/A _7608_/B vssd1 vssd1 vccd1 vccd1 _7608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7539_ _7539_/A vssd1 vssd1 vccd1 vccd1 _8361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3598_ _7370_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3598_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7890_ _7890_/CLK _7890_/D vssd1 vssd1 vccd1 vccd1 _7890_/Q sky130_fd_sc_hd__dfxtp_1
X_6910_ _6910_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__and2_1
X_6841_ _8240_/Q _7547_/A _6841_/C _7170_/A vssd1 vssd1 vccd1 vccd1 _6842_/A sky130_fd_sc_hd__and4b_1
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6086__177 _6087__178/A vssd1 vssd1 vccd1 vccd1 _7646_/CLK sky130_fd_sc_hd__inv_2
X_3984_ _8298_/Q _3959_/X _3986_/S vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__mux2_1
X_5723_ _7773_/Q _5596_/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__mux2_1
X_5654_ _5669_/S vssd1 vssd1 vccd1 vccd1 _5663_/S sky130_fd_sc_hd__clkbuf_4
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _4605_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8373_ _8373_/CLK _8373_/D vssd1 vssd1 vccd1 vccd1 _8373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5585_ _7833_/Q _5584_/X _5588_/S vssd1 vssd1 vccd1 vccd1 _5586_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4536_ _4536_/A _4536_/B _4536_/C _4536_/D vssd1 vssd1 vccd1 vccd1 _4604_/C sky130_fd_sc_hd__and4_1
Xclkbuf_0__3383_ _6920_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3383_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7255_ _8204_/Q _7202_/B _7252_/Y _7258_/B vssd1 vssd1 vccd1 vccd1 _7256_/C sky130_fd_sc_hd__a31o_1
X_4467_ _4467_/A vssd1 vssd1 vccd1 vccd1 _8092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4398_ _7989_/Q vssd1 vssd1 vccd1 vccd1 _4398_/X sky130_fd_sc_hd__buf_2
XFILLER_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6137_ _6154_/A vssd1 vssd1 vccd1 vccd1 _6137_/X sky130_fd_sc_hd__clkbuf_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6068_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__and2_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5019_ _5090_/A vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__buf_2
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3203_ clkbuf_0__3203_/X vssd1 vssd1 vccd1 vccd1 _6492__267/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7347__162 _7350__165/A vssd1 vssd1 vccd1 vccd1 _8289_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6939__491 _6941__493/A vssd1 vssd1 vccd1 vccd1 _8088_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _5370_/A vssd1 vssd1 vccd1 vccd1 _7951_/D sky130_fd_sc_hd__clkbuf_1
X_4321_ _8147_/Q _4143_/X _4321_/S vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4252_ _4249_/X _8178_/Q _4260_/S vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _8205_/Q _4099_/X _4183_/S vssd1 vssd1 vccd1 vccd1 _4184_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7942_ _8391_/CLK _7942_/D vssd1 vssd1 vccd1 vccd1 _7942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7873_ _7873_/CLK _7873_/D vssd1 vssd1 vccd1 vccd1 _7873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6755_ _7599_/A _7420_/B vssd1 vssd1 vccd1 vccd1 _6755_/X sky130_fd_sc_hd__or2_1
X_3967_ _3967_/A vssd1 vssd1 vccd1 vccd1 _6838_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5706_ _5706_/A vssd1 vssd1 vccd1 vccd1 _7781_/D sky130_fd_sc_hd__clkbuf_1
X_3898_ _3898_/A vssd1 vssd1 vccd1 vccd1 _8328_/D sky130_fd_sc_hd__clkbuf_1
X_5637_ _7812_/Q _5573_/X _5645_/S vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3398_ clkbuf_0__3398_/X vssd1 vssd1 vccd1 vccd1 _7005__545/A sky130_fd_sc_hd__clkbuf_4
X_8356_ _8397_/CLK _8356_/D vssd1 vssd1 vccd1 vccd1 _8356_/Q sky130_fd_sc_hd__dfxtp_1
X_5568_ _5567_/X _7838_/Q _5571_/S vssd1 vssd1 vccd1 vccd1 _5569_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3366_ _6851_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3366_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4519_ _4519_/A vssd1 vssd1 vccd1 vccd1 _8071_/D sky130_fd_sc_hd__clkbuf_1
X_8287_ _8287_/CLK _8287_/D vssd1 vssd1 vccd1 vccd1 _8287_/Q sky130_fd_sc_hd__dfxtp_1
X_5499_ _5288_/X _7890_/Q _5503_/S vssd1 vssd1 vccd1 vccd1 _5500_/A sky130_fd_sc_hd__mux2_1
X_7238_ _7238_/A _7238_/B _7238_/C vssd1 vssd1 vccd1 vccd1 _7238_/Y sky130_fd_sc_hd__nand3_1
X_7169_ _7173_/B _7173_/C _7173_/D vssd1 vssd1 vccd1 vccd1 _7202_/B sky130_fd_sc_hd__and3_2
XFILLER_86_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6624__329 _6625__330/A vssd1 vssd1 vccd1 vccd1 _7910_/CLK sky130_fd_sc_hd__inv_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4870_ _4562_/X _4865_/A _4869_/Y _4836_/X vssd1 vssd1 vccd1 vccd1 _8047_/D sky130_fd_sc_hd__o211a_1
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6460__241 _6462__243/A vssd1 vssd1 vccd1 vccd1 _7798_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ _3821_/A vssd1 vssd1 vccd1 vccd1 _8389_/D sky130_fd_sc_hd__clkbuf_1
X_6540_ _7579_/B _7854_/Q _6546_/S vssd1 vssd1 vccd1 vccd1 _6541_/A sky130_fd_sc_hd__mux2_1
X_6833__415 _6833__415/A vssd1 vssd1 vccd1 vccd1 _8008_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3252_ clkbuf_0__3252_/X vssd1 vssd1 vccd1 vccd1 _6643__345/A sky130_fd_sc_hd__clkbuf_4
X_6471_ _6471_/A vssd1 vssd1 vccd1 vccd1 _6471_/X sky130_fd_sc_hd__buf_1
XFILLER_9_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8210_ _8210_/CLK _8210_/D vssd1 vssd1 vccd1 vccd1 _8210_/Q sky130_fd_sc_hd__dfxtp_1
X_5422_ _5437_/S vssd1 vssd1 vccd1 vccd1 _5431_/S sky130_fd_sc_hd__buf_2
XFILLER_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5353_ _5353_/A vssd1 vssd1 vccd1 vccd1 _7958_/D sky130_fd_sc_hd__clkbuf_1
X_8141_ _8141_/CLK _8141_/D vssd1 vssd1 vccd1 vccd1 _8141_/Q sky130_fd_sc_hd__dfxtp_1
X_4304_ _4304_/A vssd1 vssd1 vccd1 vccd1 _8155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _5552_/A vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__buf_2
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8072_ _8072_/CLK _8072_/D vssd1 vssd1 vccd1 vccd1 _8072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_8 _8327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4235_ _8185_/Q _4125_/X _4241_/S vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _4414_/A _4387_/B _4413_/A vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__or3b_4
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4097_ _8266_/Q _4096_/X _4100_/S vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__mux2_1
X_7925_ _7925_/CLK _7925_/D vssd1 vssd1 vccd1 vccd1 _7925_/Q sky130_fd_sc_hd__dfxtp_1
X_7856_ _8348_/CLK _7856_/D vssd1 vssd1 vccd1 vccd1 _7856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6807_ _6807_/A vssd1 vssd1 vccd1 vccd1 _7989_/D sky130_fd_sc_hd__clkbuf_1
X_7787_ _7787_/CLK _7787_/D vssd1 vssd1 vccd1 vccd1 _7787_/Q sky130_fd_sc_hd__dfxtp_1
X_4999_ _4990_/X _4996_/X _5230_/A vssd1 vssd1 vccd1 vccd1 _4999_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6738_ _8335_/Q _6738_/B vssd1 vssd1 vccd1 vccd1 _7432_/B sky130_fd_sc_hd__xnor2_2
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6669_ _6675_/A vssd1 vssd1 vccd1 vccd1 _6669_/X sky130_fd_sc_hd__buf_1
X_8339_ _8342_/CLK _8339_/D vssd1 vssd1 vccd1 vccd1 _8339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3597_ clkbuf_0__3597_/X vssd1 vssd1 vccd1 vccd1 _7366__2/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8348_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4020_ _3884_/X _8283_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5971_ _7661_/Q _5968_/X _6079_/D vssd1 vssd1 vccd1 vccd1 _5972_/A sky130_fd_sc_hd__mux2_8
X_7710_ _7710_/CLK _7710_/D vssd1 vssd1 vccd1 vccd1 _7710_/Q sky130_fd_sc_hd__dfxtp_1
X_4922_ _8025_/Q _4401_/X _4922_/S vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__mux2_1
X_7378__12 _7381__15/A vssd1 vssd1 vccd1 vccd1 _8314_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7641_ _7143_/A _7531_/C _7641_/S vssd1 vssd1 vccd1 vccd1 _7642_/B sky130_fd_sc_hd__mux2_1
X_4853_ _4853_/A _4853_/B vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__nand2_1
X_3804_ _6234_/A _6343_/B vssd1 vssd1 vccd1 vccd1 _6285_/A sky130_fd_sc_hd__nand2_2
X_4784_ _8206_/Q _4703_/A _8023_/Q _4705_/A _4622_/A vssd1 vssd1 vccd1 vccd1 _4784_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6523_ _6523_/A vssd1 vssd1 vccd1 vccd1 _7846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ _7932_/Q _5366_/X _5413_/S vssd1 vssd1 vccd1 vccd1 _5406_/A sky130_fd_sc_hd__mux2_1
X_6385_ _7854_/Q _7747_/Q _6393_/S vssd1 vssd1 vccd1 vccd1 _6386_/A sky130_fd_sc_hd__mux2_1
X_5336_ _5336_/A vssd1 vssd1 vccd1 vccd1 _7966_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3203_ _6490_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3203_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8124_ _8124_/CLK _8124_/D vssd1 vssd1 vccd1 vccd1 _8124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5267_ _5267_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5267_/Y sky130_fd_sc_hd__nand2_1
X_8055_ _8055_/CLK _8055_/D vssd1 vssd1 vccd1 vccd1 _8055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4218_ _4217_/X _8190_/Q _4218_/S vssd1 vssd1 vccd1 vccd1 _4219_/A sky130_fd_sc_hd__mux2_1
X_7006_ _7006_/A vssd1 vssd1 vccd1 vccd1 _7006_/X sky130_fd_sc_hd__buf_1
X_6467__247 _6467__247/A vssd1 vssd1 vccd1 vccd1 _7804_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5198_ _8188_/Q _8258_/Q _5198_/S vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4149_ _4164_/S vssd1 vssd1 vccd1 vccd1 _4158_/S sky130_fd_sc_hd__buf_4
Xclkbuf_1_0_0__3382_ clkbuf_0__3382_/X vssd1 vssd1 vccd1 vccd1 _6944_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7908_ _7908_/CLK _7908_/D vssd1 vssd1 vccd1 vccd1 _7908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7839_ _7839_/CLK _7839_/D vssd1 vssd1 vccd1 vccd1 _7839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6676__366 _6677__367/A vssd1 vssd1 vccd1 vccd1 _7950_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6170_ _7536_/B _7695_/Q _6174_/S vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5121_ _8252_/Q _8166_/Q _7904_/Q _8094_/Q _5037_/A _5227_/S vssd1 vssd1 vccd1 vccd1
+ _5121_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _5045_/X _5047_/X _5051_/X _5019_/X _5095_/A vssd1 vssd1 vccd1 vccd1 _5052_/X
+ sky130_fd_sc_hd__o221a_1
X_4003_ _8290_/Q _3959_/X _4005_/S vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5954_ _5954_/A vssd1 vssd1 vccd1 vccd1 _5954_/X sky130_fd_sc_hd__clkbuf_1
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__clkbuf_1
X_4905_ _4905_/A vssd1 vssd1 vccd1 vccd1 _8033_/D sky130_fd_sc_hd__clkbuf_1
X_7624_ _7642_/A _7624_/B vssd1 vssd1 vccd1 vccd1 _7625_/A sky130_fd_sc_hd__or2_1
X_4836_ _6801_/A vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7555_ _7561_/A vssd1 vssd1 vccd1 vccd1 _7555_/X sky130_fd_sc_hd__buf_1
XFILLER_119_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4767_ _4696_/A _7963_/Q _7767_/Q _4731_/A vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__a22o_1
X_7486_ _7488_/A _7486_/B vssd1 vssd1 vccd1 vccd1 _8344_/D sky130_fd_sc_hd__nor2_1
X_6473__251 _6474__252/A vssd1 vssd1 vccd1 vccd1 _7808_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4698_ _4698_/A vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6368_ _6368_/A vssd1 vssd1 vccd1 vccd1 _7739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7341__157 _7341__157/A vssd1 vssd1 vccd1 vccd1 _8284_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5319_ _5292_/X _7973_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5320_/A sky130_fd_sc_hd__mux2_1
X_8107_ _8107_/CLK _8107_/D vssd1 vssd1 vccd1 vccd1 _8107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6299_ _7942_/Q _6301_/B _6231_/X _6244_/X vssd1 vssd1 vccd1 vccd1 _6299_/X sky130_fd_sc_hd__a31o_1
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8038_ _8038_/CLK _8038_/D vssd1 vssd1 vccd1 vccd1 _8038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3365_ clkbuf_0__3365_/X vssd1 vssd1 vccd1 vccd1 _6847__422/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6933__486 _6936__489/A vssd1 vssd1 vccd1 vccd1 _8083_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5670_ _5670_/A vssd1 vssd1 vccd1 vccd1 _7797_/D sky130_fd_sc_hd__clkbuf_1
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__clkbuf_4
X_4552_ _8046_/Q vssd1 vssd1 vccd1 vccd1 _4682_/B sky130_fd_sc_hd__buf_2
X_7271_ _8233_/Q _7277_/B vssd1 vssd1 vccd1 vccd1 _7271_/X sky130_fd_sc_hd__or2_1
X_4483_ _4483_/A vssd1 vssd1 vccd1 vccd1 _8085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6222_ _8407_/Q vssd1 vssd1 vccd1 vccd1 _7143_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6153_ _7861_/Q _6151_/X _6152_/X _6146_/X _7685_/Q vssd1 vssd1 vccd1 vccd1 _7685_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_58_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6096_/A vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__buf_1
X_5104_ _5240_/S vssd1 vssd1 vccd1 vccd1 _5224_/S sky130_fd_sc_hd__clkbuf_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _4988_/X _5032_/X _5034_/X vssd1 vssd1 vccd1 vccd1 _5035_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7036__69 _7037__70/A vssd1 vssd1 vccd1 vccd1 _8166_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5937_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7189__112 _7190__113/A vssd1 vssd1 vccd1 vccd1 _8211_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5877_/B sky130_fd_sc_hd__clkbuf_1
X_7607_ _7590_/X _7605_/Y _7606_/Y _7600_/X vssd1 vssd1 vccd1 vccd1 _8396_/D sky130_fd_sc_hd__a211oi_1
X_5799_ _4081_/X _7651_/Q _5805_/S vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4819_ _4819_/A _4819_/B _4819_/C vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__or3_1
X_7538_ _7595_/A _7538_/B _7549_/C vssd1 vssd1 vccd1 vccd1 _7539_/A sky130_fd_sc_hd__and3_1
Xclkbuf_0__3597_ _7364_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3597_/X sky130_fd_sc_hd__clkbuf_16
X_7469_ _7430_/B _7430_/C _7446_/Y _7458_/X _8337_/Q vssd1 vssd1 vccd1 vccd1 _7470_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6974__520 _6974__520/A vssd1 vssd1 vccd1 vccd1 _8117_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6424__212 _6424__212/A vssd1 vssd1 vccd1 vccd1 _7769_/CLK sky130_fd_sc_hd__inv_2
X_6840_ _6840_/A vssd1 vssd1 vccd1 vccd1 _8012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5722_ _5722_/A vssd1 vssd1 vccd1 vccd1 _7774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3983_ _3983_/A vssd1 vssd1 vccd1 vccd1 _8299_/D sky130_fd_sc_hd__clkbuf_1
X_5653_ _5689_/B _5653_/B vssd1 vssd1 vccd1 vccd1 _5669_/S sky130_fd_sc_hd__or2_2
XFILLER_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5584_ _7989_/Q vssd1 vssd1 vccd1 vccd1 _5584_/X sky130_fd_sc_hd__buf_2
X_4604_ _4604_/A _4604_/B _4604_/C vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__and3_1
X_8372_ _8372_/CLK _8372_/D vssd1 vssd1 vccd1 vccd1 _8372_/Q sky130_fd_sc_hd__dfxtp_1
X_4535_ _4843_/B _4717_/A _4056_/Y vssd1 vssd1 vccd1 vccd1 _4604_/B sky130_fd_sc_hd__o21a_1
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3382_ _6919_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3382_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7254_ _7258_/B _7254_/B vssd1 vssd1 vccd1 vccd1 _7254_/X sky130_fd_sc_hd__and2_1
X_4466_ _3837_/X _8092_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4467_/A sky130_fd_sc_hd__mux2_1
X_4397_ _4397_/A vssd1 vssd1 vccd1 vccd1 _8120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6136_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _7690_/Q _6061_/X _6039_/A _6066_/X vssd1 vssd1 vccd1 vccd1 _6067_/X sky130_fd_sc_hd__o22a_4
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5018_ _5015_/X _5016_/X _5084_/A vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__mux2_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3202_ clkbuf_0__3202_/X vssd1 vssd1 vccd1 vccd1 _6489__265/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6969_ _6975_/A vssd1 vssd1 vccd1 vccd1 _6969_/X sky130_fd_sc_hd__buf_1
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6776__382 _6777__383/A vssd1 vssd1 vccd1 vccd1 _7967_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7002__542 _7004__544/A vssd1 vssd1 vccd1 vccd1 _8139_/CLK sky130_fd_sc_hd__inv_2
X_6898__462 _6898__462/A vssd1 vssd1 vccd1 vccd1 _8057_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4320_ _4320_/A vssd1 vssd1 vccd1 vccd1 _8148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4251_ _4266_/S vssd1 vssd1 vccd1 vccd1 _4260_/S sky130_fd_sc_hd__buf_2
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6092__182 _6093__183/A vssd1 vssd1 vccd1 vccd1 _7651_/CLK sky130_fd_sc_hd__inv_2
X_4182_ _4182_/A vssd1 vssd1 vccd1 vccd1 _8206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7941_ _8359_/CLK _7941_/D vssd1 vssd1 vccd1 vccd1 _7941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8424__199 vssd1 vssd1 vccd1 vccd1 _8424__199/HI core0Index[6] sky130_fd_sc_hd__conb_1
X_7872_ _7872_/CLK _7872_/D vssd1 vssd1 vccd1 vccd1 _7872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6754_ _6754_/A _7418_/B vssd1 vssd1 vccd1 vccd1 _6754_/Y sky130_fd_sc_hd__xnor2_1
X_3966_ _8365_/Q vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__clkbuf_4
X_5705_ _7781_/Q _5596_/X _5705_/S vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__mux2_1
X_5636_ _5651_/S vssd1 vssd1 vccd1 vccd1 _5645_/S sky130_fd_sc_hd__clkbuf_4
X_3897_ _3865_/X _8328_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3397_ clkbuf_0__3397_/X vssd1 vssd1 vccd1 vccd1 _6999__540/A sky130_fd_sc_hd__clkbuf_4
X_8355_ _8397_/CLK _8355_/D vssd1 vssd1 vccd1 vccd1 _8355_/Q sky130_fd_sc_hd__dfxtp_1
X_5567_ _5567_/A vssd1 vssd1 vccd1 vccd1 _5567_/X sky130_fd_sc_hd__clkbuf_2
X_5498_ _5498_/A vssd1 vssd1 vccd1 vccd1 _7891_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3365_ _6845_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3365_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4518_ _8071_/Q _4517_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__mux2_1
X_8286_ _8286_/CLK _8286_/D vssd1 vssd1 vccd1 vccd1 _8286_/Q sky130_fd_sc_hd__dfxtp_1
X_7237_ _7237_/A _7237_/B vssd1 vssd1 vccd1 vccd1 _7237_/X sky130_fd_sc_hd__or2_1
X_4449_ _4449_/A vssd1 vssd1 vccd1 vccd1 _8100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7168_ _7155_/Y _7156_/X _7163_/X _7164_/Y _7167_/X vssd1 vssd1 vccd1 vccd1 _7173_/D
+ sky130_fd_sc_hd__o2111a_1
X_6119_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6119_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7099_ _7150_/B vssd1 vssd1 vccd1 vccd1 _7119_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3820_ _8389_/Q _3772_/X _3832_/S vssd1 vssd1 vccd1 vccd1 _3821_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3251_ clkbuf_0__3251_/X vssd1 vssd1 vccd1 vccd1 _6635__338/A sky130_fd_sc_hd__clkbuf_4
X_6987__530 _6987__530/A vssd1 vssd1 vccd1 vccd1 _8127_/CLK sky130_fd_sc_hd__inv_2
X_5421_ _5511_/B _5421_/B vssd1 vssd1 vccd1 vccd1 _5437_/S sky130_fd_sc_hd__nor2_2
X_5352_ _3822_/X _7958_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5353_/A sky130_fd_sc_hd__mux2_1
X_8140_ _8140_/CLK _8140_/D vssd1 vssd1 vccd1 vccd1 _8140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7009__548 _7010__549/A vssd1 vssd1 vccd1 vccd1 _8145_/CLK sky130_fd_sc_hd__inv_2
X_8071_ _8071_/CLK _8071_/D vssd1 vssd1 vccd1 vccd1 _8071_/Q sky130_fd_sc_hd__dfxtp_1
X_4303_ _4226_/X _8155_/Q _4303_/S vssd1 vssd1 vccd1 vccd1 _4304_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5283_ _7991_/Q vssd1 vssd1 vccd1 vccd1 _5552_/A sky130_fd_sc_hd__buf_2
XFILLER_4_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7296__121 _7298__123/A vssd1 vssd1 vccd1 vccd1 _8248_/CLK sky130_fd_sc_hd__inv_2
X_4234_ _4234_/A vssd1 vssd1 vccd1 vccd1 _8186_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_9 _8328_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4165_ _4165_/A vssd1 vssd1 vccd1 vccd1 _8241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _7986_/Q vssd1 vssd1 vccd1 vccd1 _4096_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7924_ _7924_/CLK _7924_/D vssd1 vssd1 vccd1 vccd1 _7924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7855_ _8348_/CLK _7855_/D vssd1 vssd1 vccd1 vccd1 _7855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6806_ _8354_/Q _6810_/B vssd1 vssd1 vccd1 vccd1 _6807_/A sky130_fd_sc_hd__and2_1
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7786_ _7786_/CLK _7786_/D vssd1 vssd1 vccd1 vccd1 _7786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4998_ _5090_/A vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__buf_2
X_6737_ _7135_/A _7426_/B vssd1 vssd1 vccd1 vccd1 _6737_/X sky130_fd_sc_hd__xor2_1
X_3949_ _3949_/A vssd1 vssd1 vccd1 vccd1 _8309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8407_ _8407_/CLK _8407_/D vssd1 vssd1 vccd1 vccd1 _8407_/Q sky130_fd_sc_hd__dfxtp_1
X_5619_ _5547_/X _7820_/Q _5627_/S vssd1 vssd1 vccd1 vccd1 _5620_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8338_ _8341_/CLK _8338_/D vssd1 vssd1 vccd1 vccd1 _8338_/Q sky130_fd_sc_hd__dfxtp_1
X_6099__188 _6101__190/A vssd1 vssd1 vccd1 vccd1 _7657_/CLK sky130_fd_sc_hd__inv_2
X_7305__128 _7306__129/A vssd1 vssd1 vccd1 vccd1 _8255_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6630__334 _6631__335/A vssd1 vssd1 vccd1 vccd1 _7915_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8269_ _8269_/CLK _8269_/D vssd1 vssd1 vccd1 vccd1 _8269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3596_ clkbuf_0__3596_/X vssd1 vssd1 vccd1 vccd1 _7388_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _7546_/A vssd1 vssd1 vccd1 vccd1 _6079_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4921_ _4921_/A vssd1 vssd1 vccd1 vccd1 _8026_/D sky130_fd_sc_hd__clkbuf_1
X_7640_ _7640_/A vssd1 vssd1 vccd1 vccd1 _8406_/D sky130_fd_sc_hd__clkbuf_1
X_4852_ _4852_/A vssd1 vssd1 vccd1 vccd1 _8054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3803_ _7735_/Q _3803_/B vssd1 vssd1 vccd1 vccd1 _6343_/B sky130_fd_sc_hd__nor2_2
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4783_ _4697_/A _7978_/Q _7838_/Q _4699_/A vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6522_ _7611_/B _7846_/Q _6528_/S vssd1 vssd1 vccd1 vccd1 _6523_/A sky130_fd_sc_hd__mux2_1
X_6453_ _6453_/A vssd1 vssd1 vccd1 vccd1 _6453_/X sky130_fd_sc_hd__buf_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7183__107 _7184__108/A vssd1 vssd1 vccd1 vccd1 _8206_/CLK sky130_fd_sc_hd__inv_2
X_5404_ _5419_/S vssd1 vssd1 vccd1 vccd1 _5413_/S sky130_fd_sc_hd__buf_2
X_6384_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6393_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3202_ _6484_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3202_/X sky130_fd_sc_hd__clkbuf_16
X_8123_ _8123_/CLK _8123_/D vssd1 vssd1 vccd1 vccd1 _8123_/Q sky130_fd_sc_hd__dfxtp_1
X_5335_ _5288_/X _7966_/Q _5339_/S vssd1 vssd1 vccd1 vccd1 _5336_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5266_ _7997_/Q _5265_/A _5265_/Y _5178_/X vssd1 vssd1 vccd1 vccd1 _7997_/D sky130_fd_sc_hd__o211a_1
X_8054_ _8054_/CLK _8054_/D vssd1 vssd1 vccd1 vccd1 _8054_/Q sky130_fd_sc_hd__dfxtp_1
X_4217_ _4217_/A vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5197_ _5019_/X _5185_/X _5189_/X _5265_/B _5196_/X vssd1 vssd1 vccd1 vccd1 _5197_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4148_ _5599_/A _4912_/A vssd1 vssd1 vccd1 vccd1 _4164_/S sky130_fd_sc_hd__nor2_2
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3381_ clkbuf_0__3381_/X vssd1 vssd1 vccd1 vccd1 _6918__475/A sky130_fd_sc_hd__clkbuf_4
X_4079_ _8272_/Q _4044_/X _4091_/S vssd1 vssd1 vccd1 vccd1 _4080_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7907_ _7907_/CLK _7907_/D vssd1 vssd1 vccd1 vccd1 _7907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7838_ _7838_/CLK _7838_/D vssd1 vssd1 vccd1 vccd1 _7838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7769_ _7769_/CLK _7769_/D vssd1 vssd1 vccd1 vccd1 _7769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8416__238 vssd1 vssd1 vccd1 vccd1 partID[14] _8416__238/LO sky130_fd_sc_hd__conb_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ _4990_/X _5109_/X _5118_/X _5267_/A vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__a211o_1
X_5051_ _5049_/X _5050_/X _5089_/S vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__mux2_2
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4002_/A vssd1 vssd1 vccd1 vccd1 _8291_/D sky130_fd_sc_hd__clkbuf_1
X_7048__78 _7048__78/A vssd1 vssd1 vccd1 vccd1 _8175_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ _7859_/Q _5953_/B vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__and2_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _5884_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__or2_1
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4904_ _8033_/Q _4401_/X _4904_/S vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7623_ _6719_/A _7547_/C _7635_/S vssd1 vssd1 vccd1 vccd1 _7624_/B sky130_fd_sc_hd__mux2_1
X_4835_ _4347_/X _4538_/A _4834_/X _4774_/X vssd1 vssd1 vccd1 vccd1 _8057_/D sky130_fd_sc_hd__o211a_1
X_4766_ _4729_/X _4764_/X _4765_/X vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7485_ _8344_/Q _7466_/A _7474_/X _7420_/B vssd1 vssd1 vccd1 vccd1 _7486_/B sky130_fd_sc_hd__o2bb2a_1
X_6770__377 _6772__379/A vssd1 vssd1 vccd1 vccd1 _7962_/CLK sky130_fd_sc_hd__inv_2
X_4697_ _4697_/A vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6367_ _5925_/A _7739_/Q _6371_/S vssd1 vssd1 vccd1 vccd1 _6368_/A sky130_fd_sc_hd__mux2_1
X_5318_ _5318_/A vssd1 vssd1 vccd1 vccd1 _7974_/D sky130_fd_sc_hd__clkbuf_1
X_8106_ _8106_/CLK _8106_/D vssd1 vssd1 vccd1 vccd1 _8106_/Q sky130_fd_sc_hd__dfxtp_1
X_6298_ _6221_/X _6296_/X _6297_/X _6292_/X vssd1 vssd1 vccd1 vccd1 _7719_/D sky130_fd_sc_hd__a211o_1
X_8037_ _8037_/CLK _8037_/D vssd1 vssd1 vccd1 vccd1 _8037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5249_ _5347_/B _5249_/B _5261_/B vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8365_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6892__457 _6893__458/A vssd1 vssd1 vccd1 vccd1 _8052_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6682__371 _6683__372/A vssd1 vssd1 vccd1 vccd1 _7955_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _8028_/Q _7983_/Q _7843_/Q _8211_/Q _4579_/A _4589_/X vssd1 vssd1 vccd1 vccd1
+ _4620_/X sky130_fd_sc_hd__mux4_1
X_4551_ _8047_/Q vssd1 vssd1 vccd1 vccd1 _4682_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7270_ _8004_/Q _7266_/X _7268_/X _7269_/X vssd1 vssd1 vccd1 vccd1 _8232_/D sky130_fd_sc_hd__o211a_1
X_4482_ _4341_/X _8085_/Q _4486_/S vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__mux2_1
X_6221_ _6270_/A vssd1 vssd1 vccd1 vccd1 _6221_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6152_ _6188_/A vssd1 vssd1 vccd1 vccd1 _6152_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5148_/A vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__clkbuf_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6471_/A vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__buf_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _4965_/A _5033_/X _5230_/A vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _5936_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__and2_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5867_ _5867_/A vssd1 vssd1 vccd1 vccd1 _5867_/X sky130_fd_sc_hd__clkbuf_1
X_7606_ _8396_/Q _7615_/B vssd1 vssd1 vccd1 vccd1 _7606_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5798_ _5798_/A vssd1 vssd1 vccd1 vccd1 _7652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4818_ _4750_/X _4816_/X _4817_/X vssd1 vssd1 vccd1 vccd1 _4819_/C sky130_fd_sc_hd__o21a_1
X_7537_ _7537_/A vssd1 vssd1 vccd1 vccd1 _8360_/D sky130_fd_sc_hd__clkbuf_1
X_4749_ _4743_/X _4745_/X _4865_/B _4748_/X vssd1 vssd1 vccd1 vccd1 _4749_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_0__3596_ _7363_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3596_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7468_ _7470_/A _7468_/B vssd1 vssd1 vccd1 vccd1 _8336_/D sky130_fd_sc_hd__nor2_1
X_7399_ _7399_/A input1/X vssd1 vssd1 vccd1 vccd1 _7529_/A sky130_fd_sc_hd__nor2_1
X_8445__220 vssd1 vssd1 vccd1 vccd1 _8445__220/HI partID[3] sky130_fd_sc_hd__conb_1
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3347_ clkbuf_0__3347_/X vssd1 vssd1 vccd1 vccd1 _6796__399/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6900__464 _6901__465/A vssd1 vssd1 vccd1 vccd1 _8059_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7290__116 _7291__117/A vssd1 vssd1 vccd1 vccd1 _8243_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3982_ _8299_/Q _3955_/X _3986_/S vssd1 vssd1 vccd1 vccd1 _3983_/A sky130_fd_sc_hd__mux2_1
X_5721_ _7774_/Q _5593_/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7041__73 _7041__73/A vssd1 vssd1 vccd1 vccd1 _8170_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5652_ _5652_/A vssd1 vssd1 vccd1 vccd1 _7805_/D sky130_fd_sc_hd__clkbuf_1
X_5583_ _5583_/A vssd1 vssd1 vccd1 vccd1 _7834_/D sky130_fd_sc_hd__clkbuf_1
X_4603_ _4549_/X _4577_/X _4587_/X _4602_/X vssd1 vssd1 vccd1 vccd1 _4603_/X sky130_fd_sc_hd__a31o_1
X_8371_ _8371_/CLK _8371_/D vssd1 vssd1 vccd1 vccd1 _8371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4534_ _4698_/A vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3381_ _6913_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3381_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7253_ _7262_/B _7202_/B _7252_/Y _7192_/Y vssd1 vssd1 vccd1 vccd1 _7254_/B sky130_fd_sc_hd__o211a_1
X_4465_ _4465_/A vssd1 vssd1 vccd1 vccd1 _8093_/D sky130_fd_sc_hd__clkbuf_1
X_8429__204 vssd1 vssd1 vccd1 vccd1 _8429__204/HI core1Index[4] sky130_fd_sc_hd__conb_1
X_4396_ _8120_/Q _4395_/X _4402_/S vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__mux2_1
X_6204_ _8204_/Q _6196_/X _6198_/X _7219_/A vssd1 vssd1 vccd1 vccd1 _7703_/D sky130_fd_sc_hd__a211o_1
X_6135_ _6128_/X _7851_/Q _6134_/X _6129_/X _7675_/Q vssd1 vssd1 vccd1 vccd1 _7675_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6066_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__and2_1
XFILLER_97_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5017_ _5017_/A vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__buf_2
XFILLER_85_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3201_ clkbuf_0__3201_/X vssd1 vssd1 vccd1 vccd1 _6482__259/A sky130_fd_sc_hd__clkbuf_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5919_ _5919_/A vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6486__262 _6487__263/A vssd1 vssd1 vccd1 vccd1 _7819_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7354__168 _7355__169/A vssd1 vssd1 vccd1 vccd1 _8295_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4368_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _4266_/S sky130_fd_sc_hd__or2_2
X_6649__350 _6649__350/A vssd1 vssd1 vccd1 vccd1 _7931_/CLK sky130_fd_sc_hd__inv_2
X_6946__497 _6949__500/A vssd1 vssd1 vccd1 vccd1 _8094_/CLK sky130_fd_sc_hd__inv_2
X_4181_ _8206_/Q _4096_/X _4183_/S vssd1 vssd1 vccd1 vccd1 _4182_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7940_ _7940_/CLK _7940_/D vssd1 vssd1 vccd1 vccd1 _7940_/Q sky130_fd_sc_hd__dfxtp_1
X_7871_ _7871_/CLK _7871_/D vssd1 vssd1 vccd1 vccd1 _7871_/Q sky130_fd_sc_hd__dfxtp_1
X_6822_ _6845_/A vssd1 vssd1 vccd1 vccd1 _6822_/X sky130_fd_sc_hd__buf_1
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3603_ clkbuf_0__3603_/X vssd1 vssd1 vccd1 vccd1 _7553__29/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6753_ _8341_/Q _6753_/B vssd1 vssd1 vccd1 vccd1 _7418_/B sky130_fd_sc_hd__xor2_4
X_3965_ _3965_/A vssd1 vssd1 vccd1 vccd1 _8305_/D sky130_fd_sc_hd__clkbuf_1
X_5704_ _5704_/A vssd1 vssd1 vccd1 vccd1 _7782_/D sky130_fd_sc_hd__clkbuf_1
X_3896_ _3911_/S vssd1 vssd1 vccd1 vccd1 _3905_/S sky130_fd_sc_hd__buf_2
X_5635_ _5635_/A _5795_/B vssd1 vssd1 vccd1 vccd1 _5651_/S sky130_fd_sc_hd__nor2_2
X_8354_ _8399_/CLK _8354_/D vssd1 vssd1 vccd1 vccd1 _8354_/Q sky130_fd_sc_hd__dfxtp_1
X_5566_ _5566_/A vssd1 vssd1 vccd1 vccd1 _7839_/D sky130_fd_sc_hd__clkbuf_1
X_5497_ _5284_/X _7891_/Q _5503_/S vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__mux2_1
X_4517_ _8362_/Q vssd1 vssd1 vccd1 vccd1 _4517_/X sky130_fd_sc_hd__clkbuf_2
X_8285_ _8285_/CLK _8285_/D vssd1 vssd1 vccd1 vccd1 _8285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7236_ _7233_/X _7234_/X _7251_/A vssd1 vssd1 vccd1 vccd1 _8222_/D sky130_fd_sc_hd__a21oi_1
X_4448_ _4223_/X _8100_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__mux2_1
X_7167_ _7167_/A _7167_/B vssd1 vssd1 vccd1 vccd1 _7167_/X sky130_fd_sc_hd__xor2_1
X_4379_ _4379_/A vssd1 vssd1 vccd1 vccd1 _8126_/D sky130_fd_sc_hd__clkbuf_1
X_6118_ _6118_/A vssd1 vssd1 vccd1 vccd1 _6157_/A sky130_fd_sc_hd__clkbuf_4
X_7098_ _7098_/A _7098_/B _7134_/A vssd1 vssd1 vccd1 vccd1 _7216_/A sky130_fd_sc_hd__or3_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6049_/X sky130_fd_sc_hd__and2_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7571__44 _7572__45/A vssd1 vssd1 vccd1 vccd1 _8383_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3250_ clkbuf_0__3250_/X vssd1 vssd1 vccd1 vccd1 _6628__332/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5420_ _5420_/A vssd1 vssd1 vccd1 vccd1 _7925_/D sky130_fd_sc_hd__clkbuf_1
X_5351_ _5351_/A vssd1 vssd1 vccd1 vccd1 _7959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5282_ _5282_/A vssd1 vssd1 vccd1 vccd1 _7984_/D sky130_fd_sc_hd__clkbuf_1
X_4302_ _4302_/A vssd1 vssd1 vccd1 vccd1 _8156_/D sky130_fd_sc_hd__clkbuf_1
X_8070_ _8070_/CLK _8070_/D vssd1 vssd1 vccd1 vccd1 _8070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4233_ _8186_/Q _4229_/X _4241_/S vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _8241_/Q _4099_/X _4164_/S vssd1 vssd1 vccd1 vccd1 _4165_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4095_ _4095_/A vssd1 vssd1 vccd1 vccd1 _8267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7923_ _7923_/CLK _7923_/D vssd1 vssd1 vccd1 vccd1 _7923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7854_ _7854_/CLK _7854_/D vssd1 vssd1 vccd1 vccd1 _7854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6805_ _6805_/A vssd1 vssd1 vccd1 vccd1 _7988_/D sky130_fd_sc_hd__clkbuf_1
X_7785_ _7785_/CLK _7785_/D vssd1 vssd1 vccd1 vccd1 _7785_/Q sky130_fd_sc_hd__dfxtp_1
X_6736_ _8334_/Q _7423_/B vssd1 vssd1 vccd1 vccd1 _7426_/B sky130_fd_sc_hd__xor2_2
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _5020_/B _4997_/B vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__nor2_2
X_3948_ _8309_/Q _3947_/X _3952_/S vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__mux2_1
X_6667_ _6667_/A vssd1 vssd1 vccd1 vccd1 _7943_/D sky130_fd_sc_hd__clkbuf_1
X_3879_ _3878_/X _8370_/Q _3882_/S vssd1 vssd1 vccd1 vccd1 _3880_/A sky130_fd_sc_hd__mux2_1
X_6437__223 _6437__223/A vssd1 vssd1 vccd1 vccd1 _7780_/CLK sky130_fd_sc_hd__inv_2
X_8406_ _8407_/CLK _8406_/D vssd1 vssd1 vccd1 vccd1 _8406_/Q sky130_fd_sc_hd__dfxtp_2
X_5618_ _5633_/S vssd1 vssd1 vccd1 vccd1 _5627_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8337_ _8341_/CLK _8337_/D vssd1 vssd1 vccd1 vccd1 _8337_/Q sky130_fd_sc_hd__dfxtp_1
X_6849__424 _6850__425/A vssd1 vssd1 vccd1 vccd1 _8019_/CLK sky130_fd_sc_hd__inv_2
X_5549_ _5571_/S vssd1 vssd1 vccd1 vccd1 _5562_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_117_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3347_ _6792_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3347_/X sky130_fd_sc_hd__clkbuf_16
X_8268_ _8268_/CLK _8268_/D vssd1 vssd1 vccd1 vccd1 _8268_/Q sky130_fd_sc_hd__dfxtp_1
X_8199_ _8199_/CLK _8199_/D vssd1 vssd1 vccd1 vccd1 _8199_/Q sky130_fd_sc_hd__dfxtp_1
X_7219_ _7219_/A vssd1 vssd1 vccd1 vccd1 _7244_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3595_ clkbuf_0__3595_/X vssd1 vssd1 vccd1 vccd1 _7362__175/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7369__5 _7369__5/A vssd1 vssd1 vccd1 vccd1 _8307_/CLK sky130_fd_sc_hd__inv_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6856__428 _6857__429/A vssd1 vssd1 vccd1 vccd1 _8023_/CLK sky130_fd_sc_hd__inv_2
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6789__393 _6790__394/A vssd1 vssd1 vccd1 vccd1 _7978_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8239_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2973_ clkbuf_0__2973_/X vssd1 vssd1 vccd1 vccd1 _6471_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4920_ _8026_/Q _4398_/X _4922_/S vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4851_ _6907_/C _4851_/B _4851_/C vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__and3_1
XFILLER_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3802_ _7736_/Q _7737_/Q _7738_/Q _7739_/Q vssd1 vssd1 vccd1 vccd1 _3803_/B sky130_fd_sc_hd__or4_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _4776_/X _4778_/X _4865_/B _4781_/X vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__a211o_1
X_6521_ _6521_/A vssd1 vssd1 vccd1 vccd1 _7845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3387_ clkbuf_0__3387_/X vssd1 vssd1 vccd1 vccd1 _6949__500/A sky130_fd_sc_hd__clkbuf_16
XFILLER_118_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5403_ _5475_/A _5421_/B vssd1 vssd1 vccd1 vccd1 _5419_/S sky130_fd_sc_hd__nor2_2
X_6383_ _6383_/A vssd1 vssd1 vccd1 vccd1 _7746_/D sky130_fd_sc_hd__clkbuf_1
X_8122_ _8122_/CLK _8122_/D vssd1 vssd1 vccd1 vccd1 _8122_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3201_ _6478_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3201_/X sky130_fd_sc_hd__clkbuf_16
X_5334_ _5334_/A vssd1 vssd1 vccd1 vccd1 _7967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5265_ _5265_/A _5265_/B vssd1 vssd1 vccd1 vccd1 _5265_/Y sky130_fd_sc_hd__nand2_1
X_8053_ _8053_/CLK _8053_/D vssd1 vssd1 vccd1 vccd1 _8053_/Q sky130_fd_sc_hd__dfxtp_1
X_5196_ _5191_/X _5192_/X _5267_/A _5195_/X vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__a211o_1
X_4216_ _4216_/A vssd1 vssd1 vccd1 vccd1 _8191_/D sky130_fd_sc_hd__clkbuf_1
X_4147_ _5795_/A vssd1 vssd1 vccd1 vccd1 _4912_/A sky130_fd_sc_hd__buf_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4100_/S vssd1 vssd1 vccd1 vccd1 _4091_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7906_ _7906_/CLK _7906_/D vssd1 vssd1 vccd1 vccd1 _7906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7837_ _7837_/CLK _7837_/D vssd1 vssd1 vccd1 vccd1 _7837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7384__17 _7385__18/A vssd1 vssd1 vccd1 vccd1 _8319_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7311__133 _7311__133/A vssd1 vssd1 vccd1 vccd1 _8260_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7768_ _7768_/CLK _7768_/D vssd1 vssd1 vccd1 vccd1 _7768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7699_ _7846_/CLK _7699_/D vssd1 vssd1 vccd1 vccd1 _7699_/Q sky130_fd_sc_hd__dfxtp_1
X_6719_ _6719_/A _7430_/B _7430_/C vssd1 vssd1 vccd1 vccd1 _6719_/X sky130_fd_sc_hd__and3_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7371__6 _7372__7/A vssd1 vssd1 vccd1 vccd1 _8308_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3241_ clkbuf_0__3241_/X vssd1 vssd1 vccd1 vccd1 _6650_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5050_ _8153_/Q _8137_/Q _8129_/Q _8161_/Q _5204_/S _5037_/X vssd1 vssd1 vccd1 vccd1
+ _5050_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4001_ _8291_/Q _3955_/X _4005_/S vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5952_ _5952_/A vssd1 vssd1 vccd1 vccd1 _5952_/X sky130_fd_sc_hd__clkbuf_1
X_4903_ _4903_/A vssd1 vssd1 vccd1 vccd1 _8034_/D sky130_fd_sc_hd__clkbuf_1
X_5883_ _5883_/A vssd1 vssd1 vccd1 vccd1 _5883_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7622_ _7617_/Y _7627_/B _7621_/Y _7600_/X vssd1 vssd1 vccd1 vccd1 _8400_/D sky130_fd_sc_hd__a211oi_1
X_4834_ _4540_/A _8057_/Q _4872_/B _4833_/X _4605_/A vssd1 vssd1 vccd1 vccd1 _4834_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4765_ _4724_/A _7759_/Q _4725_/A _8016_/Q _4726_/A vssd1 vssd1 vccd1 vccd1 _4765_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7484_ _7488_/A _7484_/B vssd1 vssd1 vccd1 vccd1 _8343_/D sky130_fd_sc_hd__nor2_1
X_4696_ _4696_/A vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6366_ _6366_/A vssd1 vssd1 vccd1 vccd1 _7738_/D sky130_fd_sc_hd__clkbuf_1
X_5317_ _5288_/X _7974_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5318_/A sky130_fd_sc_hd__mux2_1
X_8105_ _8105_/CLK _8105_/D vssd1 vssd1 vccd1 vccd1 _8105_/Q sky130_fd_sc_hd__dfxtp_1
X_8036_ _8036_/CLK _8036_/D vssd1 vssd1 vccd1 vccd1 _8036_/Q sky130_fd_sc_hd__dfxtp_1
X_6297_ _7719_/Q _7546_/C vssd1 vssd1 vccd1 vccd1 _6297_/X sky130_fd_sc_hd__and2_1
XFILLER_29_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5248_ _8003_/Q _8012_/Q _3968_/B _5178_/X vssd1 vssd1 vccd1 vccd1 _8003_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5179_ _3884_/X _5029_/X _5177_/X _5178_/X vssd1 vssd1 vccd1 vccd1 _8006_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6480__257 _6482__259/A vssd1 vssd1 vccd1 vccd1 _7814_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7318__139 _7319__140/A vssd1 vssd1 vccd1 vccd1 _8266_/CLK sky130_fd_sc_hd__inv_2
X_6643__345 _6643__345/A vssd1 vssd1 vccd1 vccd1 _7926_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7053__82 _7055__84/A vssd1 vssd1 vccd1 vccd1 _8179_/CLK sky130_fd_sc_hd__inv_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4564_/A vssd1 vssd1 vccd1 vccd1 _4573_/B sky130_fd_sc_hd__clkbuf_2
X_4481_ _4481_/A vssd1 vssd1 vccd1 vccd1 _8086_/D sky130_fd_sc_hd__clkbuf_1
X_6220_ _7540_/B vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6151_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6151_/X sky130_fd_sc_hd__clkbuf_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6851_/A vssd1 vssd1 vccd1 vccd1 _6082_/X sky130_fd_sc_hd__buf_1
XFILLER_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _8279_/Q _8263_/Q _8193_/Q _8287_/Q _5231_/S _5010_/X vssd1 vssd1 vccd1 vccd1
+ _5033_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5935_ _5935_/A vssd1 vssd1 vccd1 vccd1 _5935_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5866_ _7595_/B _5866_/B vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__or2_1
X_7605_ _7614_/A _7605_/B vssd1 vssd1 vccd1 vccd1 _7605_/Y sky130_fd_sc_hd__nand2_1
X_4817_ _8205_/Q _4724_/X _8022_/Q _4681_/A _4622_/A vssd1 vssd1 vccd1 vccd1 _4817_/X
+ sky130_fd_sc_hd__o221a_1
X_5797_ _4044_/X _7652_/Q _5805_/S vssd1 vssd1 vccd1 vccd1 _5798_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7536_ _7595_/A _7536_/B _7549_/C vssd1 vssd1 vccd1 vccd1 _7537_/A sky130_fd_sc_hd__and3_1
Xclkbuf_0__3595_ _7357_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3595_/X sky130_fd_sc_hd__clkbuf_16
X_4748_ _4869_/B _4746_/X _4747_/X vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__o21a_1
X_7467_ _8336_/Q _7466_/X _7461_/X _7429_/Y vssd1 vssd1 vccd1 vccd1 _7468_/B sky130_fd_sc_hd__o2bb2a_1
X_4679_ _4704_/A vssd1 vssd1 vccd1 vccd1 _4725_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7398_ _7450_/A _7450_/B vssd1 vssd1 vccd1 vccd1 _7447_/B sky130_fd_sc_hd__nand2_2
X_6349_ _6349_/A _6687_/A _6349_/C _6349_/D vssd1 vssd1 vccd1 vccd1 _6350_/D sky130_fd_sc_hd__nand4_2
XFILLER_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8019_ _8019_/CLK _8019_/D vssd1 vssd1 vccd1 vccd1 _8019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3346_ clkbuf_0__3346_/X vssd1 vssd1 vccd1 vccd1 _6790__394/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3361_ clkbuf_0__3361_/X vssd1 vssd1 vccd1 vccd1 _6837__418/A sky130_fd_sc_hd__clkbuf_16
XFILLER_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6829__411 _6830__412/A vssd1 vssd1 vccd1 vccd1 _8004_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _3981_/A vssd1 vssd1 vccd1 vccd1 _8300_/D sky130_fd_sc_hd__clkbuf_1
X_5720_ _5720_/A vssd1 vssd1 vccd1 vccd1 _7775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _7805_/Q _5596_/X _5651_/S vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__mux2_1
X_5582_ _7834_/Q _5581_/X _5588_/S vssd1 vssd1 vccd1 vccd1 _5583_/A sky130_fd_sc_hd__mux2_1
X_4602_ _4588_/X _4593_/X _4600_/X _4674_/A vssd1 vssd1 vccd1 vccd1 _4602_/X sky130_fd_sc_hd__o211a_1
X_8370_ _8370_/CLK _8370_/D vssd1 vssd1 vccd1 vccd1 _8370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4533_ _4731_/A vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__clkbuf_2
X_7252_ _7262_/C _7252_/B vssd1 vssd1 vccd1 vccd1 _7252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6203_ _7235_/A vssd1 vssd1 vccd1 vccd1 _7219_/A sky130_fd_sc_hd__buf_2
X_6431__218 _6432__219/A vssd1 vssd1 vccd1 vccd1 _7775_/CLK sky130_fd_sc_hd__inv_2
X_4464_ _3834_/X _8093_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__mux2_1
X_4395_ _7990_/Q vssd1 vssd1 vccd1 vccd1 _4395_/X sky130_fd_sc_hd__buf_2
X_6134_ _6188_/A vssd1 vssd1 vccd1 vccd1 _6134_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6843__419 _6844__420/A vssd1 vssd1 vccd1 vccd1 _8014_/CLK sky130_fd_sc_hd__inv_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _7689_/Q _6061_/X _6039_/A _6064_/X vssd1 vssd1 vccd1 vccd1 _6065_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5016_ _8256_/Q _8170_/Q _7908_/Q _8098_/Q _4995_/A _5181_/A vssd1 vssd1 vccd1 vccd1
+ _5016_/X sky130_fd_sc_hd__mux4_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3200_ clkbuf_0__3200_/X vssd1 vssd1 vccd1 vccd1 _6474__252/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6958__506 _6962__510/A vssd1 vssd1 vccd1 vccd1 _8103_/CLK sky130_fd_sc_hd__inv_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5918_ _5918_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__and2_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5849_ _7546_/B _5855_/B vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__or2_1
X_6592__303 _6592__303/A vssd1 vssd1 vccd1 vccd1 _7884_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7519_ _7519_/A vssd1 vssd1 vccd1 vccd1 _7519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6783__388 _6785__390/A vssd1 vssd1 vccd1 vccd1 _7973_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4180_ _4180_/A vssd1 vssd1 vccd1 vccd1 _8207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7870_ _7870_/CLK _7870_/D vssd1 vssd1 vccd1 vccd1 _7870_/Q sky130_fd_sc_hd__dfxtp_1
X_6580__295 _6580__295/A vssd1 vssd1 vccd1 vccd1 _7876_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3602_ clkbuf_0__3602_/X vssd1 vssd1 vccd1 vccd1 _7561_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6752_ _8397_/Q vssd1 vssd1 vccd1 vccd1 _6754_/A sky130_fd_sc_hd__inv_2
X_3964_ _8305_/Q _3963_/X _3964_/S vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__mux2_1
X_3895_ _4507_/A _4368_/A vssd1 vssd1 vccd1 vccd1 _3911_/S sky130_fd_sc_hd__or2_4
X_5703_ _7782_/Q _5593_/X _5705_/S vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__mux2_1
X_5634_ _5634_/A vssd1 vssd1 vccd1 vccd1 _7813_/D sky130_fd_sc_hd__clkbuf_1
X_6656__355 _6656__355/A vssd1 vssd1 vccd1 vccd1 _7936_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8353_ _8399_/CLK _8353_/D vssd1 vssd1 vccd1 vccd1 _8353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5565_ _5564_/X _7839_/Q _5571_/S vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5496_ _5496_/A vssd1 vssd1 vccd1 vccd1 _7892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4516_ _4516_/A vssd1 vssd1 vccd1 vccd1 _8072_/D sky130_fd_sc_hd__clkbuf_1
X_8284_ _8284_/CLK _8284_/D vssd1 vssd1 vccd1 vccd1 _8284_/Q sky130_fd_sc_hd__dfxtp_1
X_7235_ _7235_/A vssd1 vssd1 vccd1 vccd1 _7251_/A sky130_fd_sc_hd__clkbuf_2
X_4447_ _4447_/A vssd1 vssd1 vccd1 vccd1 _8101_/D sky130_fd_sc_hd__clkbuf_1
X_7166_ _7166_/A _7165_/X vssd1 vssd1 vccd1 vccd1 _7167_/B sky130_fd_sc_hd__or2b_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6117_ _6104_/X _7697_/Q _6116_/X _6111_/X _7665_/Q vssd1 vssd1 vccd1 vccd1 _7665_/D
+ sky130_fd_sc_hd__o32a_1
X_4378_ _4217_/X _8126_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__mux2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7097_ _7221_/A _7221_/B _7096_/A vssd1 vssd1 vccd1 vccd1 _7104_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6048_ _6079_/D vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__buf_2
XFILLER_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6600__310 _6600__310/A vssd1 vssd1 vccd1 vccd1 _7891_/CLK sky130_fd_sc_hd__inv_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _7999_/CLK _7999_/D vssd1 vssd1 vccd1 vccd1 _7999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7556__31 _7559__34/A vssd1 vssd1 vccd1 vccd1 _8370_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7360__173 _7362__175/A vssd1 vssd1 vccd1 vccd1 _8300_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6599__309 _6600__310/A vssd1 vssd1 vccd1 vccd1 _7890_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5350_ _3772_/X _7959_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5351_/A sky130_fd_sc_hd__mux2_1
X_5281_ _5278_/X _7984_/Q _5297_/S vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4301_ _4223_/X _8156_/Q _4303_/S vssd1 vssd1 vccd1 vccd1 _4302_/A sky130_fd_sc_hd__mux2_1
X_7020_ _7038_/A vssd1 vssd1 vccd1 vccd1 _7020_/X sky130_fd_sc_hd__buf_1
X_4232_ _4247_/S vssd1 vssd1 vccd1 vccd1 _4241_/S sky130_fd_sc_hd__clkbuf_4
X_4163_ _4163_/A vssd1 vssd1 vccd1 vccd1 _8242_/D sky130_fd_sc_hd__clkbuf_1
X_4094_ _8267_/Q _4093_/X _4100_/S vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7922_ _7922_/CLK _7922_/D vssd1 vssd1 vccd1 vccd1 _7922_/Q sky130_fd_sc_hd__dfxtp_1
X_6211__197 _6213__199/A vssd1 vssd1 vccd1 vccd1 _7709_/CLK sky130_fd_sc_hd__inv_2
X_7853_ _7854_/CLK _7853_/D vssd1 vssd1 vccd1 vccd1 _7853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7396__26 _7554__30/A vssd1 vssd1 vccd1 vccd1 _8328_/CLK sky130_fd_sc_hd__inv_2
X_6804_ _8353_/Q _6810_/B vssd1 vssd1 vccd1 vccd1 _6805_/A sky130_fd_sc_hd__and2_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7784_ _7784_/CLK _7784_/D vssd1 vssd1 vccd1 vccd1 _7784_/Q sky130_fd_sc_hd__dfxtp_1
X_4996_ _8280_/Q _8264_/Q _8194_/Q _8288_/Q _5227_/S _4995_/X vssd1 vssd1 vccd1 vccd1
+ _4996_/X sky130_fd_sc_hd__mux4_1
X_6735_ _6727_/X _6729_/Y _6731_/Y _6733_/Y _6734_/X vssd1 vssd1 vccd1 vccd1 _6735_/X
+ sky130_fd_sc_hd__o2111a_1
X_3947_ _4214_/A vssd1 vssd1 vccd1 vccd1 _3947_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6666_ _6536_/A _7943_/Q _6666_/S vssd1 vssd1 vccd1 vccd1 _6667_/A sky130_fd_sc_hd__mux2_1
X_3878_ _8362_/Q vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__clkbuf_4
X_8405_ _8407_/CLK _8405_/D vssd1 vssd1 vccd1 vccd1 _8405_/Q sky130_fd_sc_hd__dfxtp_1
X_5617_ _5689_/B _5617_/B vssd1 vssd1 vccd1 vccd1 _5633_/S sky130_fd_sc_hd__or2_2
X_8336_ _8341_/CLK _8336_/D vssd1 vssd1 vccd1 vccd1 _8336_/Q sky130_fd_sc_hd__dfxtp_1
X_5548_ _5548_/A _5617_/B vssd1 vssd1 vccd1 vccd1 _5571_/S sky130_fd_sc_hd__or2_2
Xclkbuf_0__3346_ _6786_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3346_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8267_ _8267_/CLK _8267_/D vssd1 vssd1 vccd1 vccd1 _8267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7218_ _7218_/A _7218_/B vssd1 vssd1 vccd1 vccd1 _8218_/D sky130_fd_sc_hd__nor2_1
X_5479_ _7899_/Q _4208_/A _5485_/S vssd1 vssd1 vccd1 vccd1 _5480_/A sky130_fd_sc_hd__mux2_1
X_8198_ _8198_/CLK _8198_/D vssd1 vssd1 vccd1 vccd1 _8198_/Q sky130_fd_sc_hd__dfxtp_1
X_7149_ _8226_/Q vssd1 vssd1 vccd1 vccd1 _7151_/B sky130_fd_sc_hd__inv_2
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3594_ clkbuf_0__3594_/X vssd1 vssd1 vccd1 vccd1 _7355__169/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6444__228 _6446__230/A vssd1 vssd1 vccd1 vccd1 _7785_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4850_ _4604_/A _4853_/A _6253_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _4851_/C sky130_fd_sc_hd__a31o_1
XFILLER_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3801_ _7734_/Q vssd1 vssd1 vccd1 vccd1 _6234_/A sky130_fd_sc_hd__inv_2
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6499__273 _6500__274/A vssd1 vssd1 vccd1 vccd1 _7830_/CLK sky130_fd_sc_hd__inv_2
X_6520_ _7614_/B _7845_/Q _6528_/S vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__mux2_1
X_4781_ _4869_/B _4779_/X _4780_/X vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3386_ clkbuf_0__3386_/X vssd1 vssd1 vccd1 vccd1 _6943__495/A sky130_fd_sc_hd__clkbuf_16
X_6382_ _7853_/Q _7746_/Q _6382_/S vssd1 vssd1 vccd1 vccd1 _6383_/A sky130_fd_sc_hd__mux2_1
X_5402_ _5402_/A vssd1 vssd1 vccd1 vccd1 _7933_/D sky130_fd_sc_hd__clkbuf_1
X_5333_ _5284_/X _7967_/Q _5339_/S vssd1 vssd1 vccd1 vccd1 _5334_/A sky130_fd_sc_hd__mux2_1
X_8121_ _8121_/CLK _8121_/D vssd1 vssd1 vccd1 vccd1 _8121_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3200_ _6472_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3200_/X sky130_fd_sc_hd__clkbuf_16
X_5264_ _5274_/B vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8052_ _8052_/CLK _8052_/D vssd1 vssd1 vccd1 vccd1 _8052_/Q sky130_fd_sc_hd__dfxtp_1
X_5195_ _5191_/A _5193_/X _5194_/X _4990_/X vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__o211a_1
X_4215_ _4214_/X _8191_/Q _4218_/S vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4146_ _4324_/B _4843_/A _4843_/B vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__or3b_4
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _5599_/A _5635_/A vssd1 vssd1 vccd1 vccd1 _4100_/S sky130_fd_sc_hd__nor2_2
XFILLER_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7905_ _7905_/CLK _7905_/D vssd1 vssd1 vccd1 vccd1 _7905_/Q sky130_fd_sc_hd__dfxtp_1
X_7836_ _7836_/CLK _7836_/D vssd1 vssd1 vccd1 vccd1 _7836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _8186_/Q _8178_/Q _7900_/Q _7916_/Q _4971_/A _4978_/X vssd1 vssd1 vccd1 vccd1
+ _4979_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7767_ _7767_/CLK _7767_/D vssd1 vssd1 vccd1 vccd1 _7767_/Q sky130_fd_sc_hd__dfxtp_1
X_7698_ _7846_/CLK _7698_/D vssd1 vssd1 vccd1 vccd1 _7698_/Q sky130_fd_sc_hd__dfxtp_1
X_6718_ _7430_/B _7430_/C _6719_/A vssd1 vssd1 vccd1 vccd1 _6718_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8319_ _8319_/CLK _8319_/D vssd1 vssd1 vccd1 vccd1 _8319_/Q sky130_fd_sc_hd__dfxtp_1
X_6862__433 _6863__434/A vssd1 vssd1 vccd1 vccd1 _8028_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6823__406 _6827__410/A vssd1 vssd1 vccd1 vccd1 _7999_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _8292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5951_ _7858_/Q _5953_/B vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__and2_1
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4902_ _8034_/Q _4398_/X _4904_/S vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5882_ _5882_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__or2_1
X_7621_ _7621_/A _7627_/B vssd1 vssd1 vccd1 vccd1 _7621_/Y sky130_fd_sc_hd__nor2_1
X_4833_ _4863_/B _4812_/X _4819_/X _4832_/X vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__a31o_2
X_4764_ _4730_/X _7871_/Q _7775_/Q _4731_/X vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7483_ _8343_/Q _7466_/X _7474_/X _6706_/B vssd1 vssd1 vccd1 vccd1 _7484_/B sky130_fd_sc_hd__o2bb2a_1
X_6503_ _6575_/A vssd1 vssd1 vccd1 vccd1 _6503_/X sky130_fd_sc_hd__buf_1
X_6434_ _6434_/A vssd1 vssd1 vccd1 vccd1 _6434_/X sky130_fd_sc_hd__buf_1
X_4695_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4869_/B sky130_fd_sc_hd__clkbuf_4
X_6365_ _5923_/A _7738_/Q _6371_/S vssd1 vssd1 vccd1 vccd1 _6366_/A sky130_fd_sc_hd__mux2_1
X_5316_ _5316_/A vssd1 vssd1 vccd1 vccd1 _7975_/D sky130_fd_sc_hd__clkbuf_1
X_6296_ _7621_/A _6839_/C _6312_/A _6289_/X _6295_/X vssd1 vssd1 vccd1 vccd1 _6296_/X
+ sky130_fd_sc_hd__a32o_1
X_8104_ _8104_/CLK _8104_/D vssd1 vssd1 vccd1 vccd1 _8104_/Q sky130_fd_sc_hd__dfxtp_1
X_8035_ _8035_/CLK _8035_/D vssd1 vssd1 vccd1 vccd1 _8035_/Q sky130_fd_sc_hd__dfxtp_1
X_5247_ _3890_/X _5029_/A _5246_/X _5178_/X vssd1 vssd1 vccd1 vccd1 _8004_/D sky130_fd_sc_hd__o211a_1
X_5178_ _7533_/A vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__buf_2
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4129_ _8254_/Q _4128_/X _4135_/S vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7819_ _7819_/CLK _7819_/D vssd1 vssd1 vccd1 vccd1 _7819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6869__439 _6870__440/A vssd1 vssd1 vccd1 vccd1 _8034_/CLK sky130_fd_sc_hd__inv_2
X_4480_ _4338_/X _8086_/Q _4480_/S vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__mux2_1
X_6150_ _6145_/X _7860_/Q _6142_/X _6146_/X _7684_/Q vssd1 vssd1 vccd1 vccd1 _7684_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5115_/A _5101_/B vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__nand2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A vssd1 vssd1 vccd1 vccd1 _6081_/X sky130_fd_sc_hd__buf_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _8380_/Q _7950_/Q _7883_/Q _8372_/Q _5198_/S _4971_/X vssd1 vssd1 vccd1 vccd1
+ _5032_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_10_wb_clk_i _7717_/CLK vssd1 vssd1 vccd1 vccd1 _8391_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5934_ _5934_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__and2_1
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5865_ _5865_/A vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__clkbuf_1
X_7604_ _6032_/X _5862_/A _7590_/X _7603_/X vssd1 vssd1 vccd1 vccd1 _8395_/D sky130_fd_sc_hd__a31o_1
X_4816_ _4697_/A _7977_/Q _7837_/Q _4699_/A vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__a22o_1
X_5796_ _5811_/S vssd1 vssd1 vccd1 vccd1 _5805_/S sky130_fd_sc_hd__clkbuf_4
X_7535_ _7535_/A vssd1 vssd1 vccd1 vccd1 _7549_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__3594_ _7351_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3594_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4747_ _4703_/X _7807_/Q _7647_/Q _4705_/X _4669_/S vssd1 vssd1 vccd1 vccd1 _4747_/X
+ sky130_fd_sc_hd__o221a_1
X_7466_ _7466_/A vssd1 vssd1 vccd1 vccd1 _7466_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4678_ _4682_/A _8046_/Q vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__or2_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7397_ _8329_/Q vssd1 vssd1 vccd1 vccd1 _7450_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6348_ _7731_/Q _6405_/B _6347_/Y _6251_/X vssd1 vssd1 vccd1 vccd1 _7731_/D sky130_fd_sc_hd__o211a_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6279_ _8062_/Q _6231_/A _6201_/X _6235_/X vssd1 vssd1 vccd1 vccd1 _6279_/X sky130_fd_sc_hd__a31o_1
X_8018_ _8018_/CLK _8018_/D vssd1 vssd1 vccd1 vccd1 _8018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3414_ clkbuf_0__3414_/X vssd1 vssd1 vccd1 vccd1 _7081__105/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3345_ clkbuf_0__3345_/X vssd1 vssd1 vccd1 vccd1 _6782__387/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7324__144 _7325__145/A vssd1 vssd1 vccd1 vccd1 _8271_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _8300_/Q _3951_/X _3980_/S vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5650_ _5650_/A vssd1 vssd1 vccd1 vccd1 _7806_/D sky130_fd_sc_hd__clkbuf_1
X_4601_ _8050_/Q _4601_/B vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__xnor2_4
X_6916__473 _6918__475/A vssd1 vssd1 vccd1 vccd1 _8070_/CLK sky130_fd_sc_hd__inv_2
X_5581_ _7990_/Q vssd1 vssd1 vccd1 vccd1 _5581_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _8065_/Q vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7320_ _7320_/A vssd1 vssd1 vccd1 vccd1 _7320_/X sky130_fd_sc_hd__buf_1
X_7251_ _7251_/A _7251_/B vssd1 vssd1 vccd1 vccd1 _8228_/D sky130_fd_sc_hd__nor2_1
X_4463_ _4463_/A vssd1 vssd1 vccd1 vccd1 _8094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _3814_/X _7533_/B _6201_/X _6144_/A vssd1 vssd1 vccd1 vccd1 _7235_/A sky130_fd_sc_hd__a31o_1
X_4394_ _4394_/A vssd1 vssd1 vccd1 vccd1 _8121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6133_ _6128_/X _7850_/Q _6126_/X _6129_/X _7674_/Q vssd1 vssd1 vccd1 vccd1 _7674_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6064_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6064_/X sky130_fd_sc_hd__and2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5015_ _8154_/Q _8138_/Q _8130_/Q _8162_/Q _5204_/S _4971_/A vssd1 vssd1 vccd1 vccd1
+ _5015_/X sky130_fd_sc_hd__mux4_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5917_ _5917_/A vssd1 vssd1 vccd1 vccd1 _5917_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5848_ _5848_/A vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__clkbuf_1
X_5779_ _7660_/Q _5547_/A _5785_/S vssd1 vssd1 vccd1 vccd1 _5780_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7518_ _8353_/Q _7523_/B _7513_/X vssd1 vssd1 vccd1 vccd1 _7518_/X sky130_fd_sc_hd__or3b_1
XFILLER_107_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7449_ _7447_/A _7446_/Y _7447_/Y _7448_/X vssd1 vssd1 vccd1 vccd1 _8331_/D sky130_fd_sc_hd__o211a_1
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6493__268 _6495__270/A vssd1 vssd1 vccd1 vccd1 _7825_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3601_ clkbuf_0__3601_/X vssd1 vssd1 vccd1 vccd1 _7390__22/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6751_ _7599_/A _7420_/B vssd1 vssd1 vccd1 vccd1 _6751_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8435__210 vssd1 vssd1 vccd1 vccd1 _8435__210/HI manufacturerID[2] sky130_fd_sc_hd__conb_1
X_3963_ _4226_/A vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__buf_2
XFILLER_16_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_3894_ _3967_/A _3894_/B vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__nand2_2
X_5702_ _5702_/A vssd1 vssd1 vccd1 vccd1 _7783_/D sky130_fd_sc_hd__clkbuf_1
X_5633_ _5570_/X _7813_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3394_ clkbuf_0__3394_/X vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__clkbuf_4
X_8352_ _8399_/CLK _8352_/D vssd1 vssd1 vccd1 vccd1 _8352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5564_ _5564_/A vssd1 vssd1 vccd1 vccd1 _5564_/X sky130_fd_sc_hd__buf_2
X_4515_ _8072_/Q _4514_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5495_ _5278_/X _7892_/Q _5503_/S vssd1 vssd1 vccd1 vccd1 _5496_/A sky130_fd_sc_hd__mux2_1
X_6964__511 _6966__513/A vssd1 vssd1 vccd1 vccd1 _8108_/CLK sky130_fd_sc_hd__inv_2
X_8283_ _8283_/CLK _8283_/D vssd1 vssd1 vccd1 vccd1 _8283_/Q sky130_fd_sc_hd__dfxtp_1
X_7234_ _7234_/A _7234_/B _7238_/C vssd1 vssd1 vccd1 vccd1 _7234_/X sky130_fd_sc_hd__or3b_1
X_4446_ _4220_/X _8101_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7165_ _7159_/A _7159_/B _7150_/D _8225_/Q vssd1 vssd1 vccd1 vccd1 _7165_/X sky130_fd_sc_hd__a31o_1
X_4377_ _4377_/A vssd1 vssd1 vccd1 vccd1 _8127_/D sky130_fd_sc_hd__clkbuf_1
X_6116_ _6116_/A vssd1 vssd1 vccd1 vccd1 _6116_/X sky130_fd_sc_hd__buf_4
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/A _7221_/A _7221_/B vssd1 vssd1 vccd1 vccd1 _7104_/A sky130_fd_sc_hd__and3_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _7682_/Q _6032_/X _6039_/X _6046_/X vssd1 vssd1 vccd1 vccd1 _6047_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7998_ _7998_/CLK _7998_/D vssd1 vssd1 vccd1 vccd1 _7998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6501__275 _6501__275/A vssd1 vssd1 vccd1 vccd1 _7832_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5280_ _5309_/S vssd1 vssd1 vccd1 vccd1 _5297_/S sky130_fd_sc_hd__buf_4
X_4300_ _4300_/A vssd1 vssd1 vccd1 vccd1 _8157_/D sky130_fd_sc_hd__clkbuf_1
X_4231_ _5385_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _4247_/S sky130_fd_sc_hd__nor2_2
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4162_ _8242_/Q _4096_/X _4164_/S vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4093_ _7987_/Q vssd1 vssd1 vccd1 vccd1 _4093_/X sky130_fd_sc_hd__buf_2
X_7337__154 _7338__155/A vssd1 vssd1 vccd1 vccd1 _8281_/CLK sky130_fd_sc_hd__inv_2
X_7921_ _7921_/CLK _7921_/D vssd1 vssd1 vccd1 vccd1 _7921_/Q sky130_fd_sc_hd__dfxtp_1
X_7852_ _7854_/CLK _7852_/D vssd1 vssd1 vccd1 vccd1 _7852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6803_ _6803_/A vssd1 vssd1 vccd1 vccd1 _7987_/D sky130_fd_sc_hd__clkbuf_1
X_7783_ _7783_/CLK _7783_/D vssd1 vssd1 vccd1 vccd1 _7783_/Q sky130_fd_sc_hd__dfxtp_1
X_4995_ _4995_/A vssd1 vssd1 vccd1 vccd1 _4995_/X sky130_fd_sc_hd__buf_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6734_ _8407_/Q _7447_/A vssd1 vssd1 vccd1 vccd1 _6734_/X sky130_fd_sc_hd__or2_1
X_3946_ _8362_/Q vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__buf_2
X_6665_ _6665_/A vssd1 vssd1 vccd1 vccd1 _7942_/D sky130_fd_sc_hd__clkbuf_1
X_8404_ _8407_/CLK _8404_/D vssd1 vssd1 vccd1 vccd1 _8404_/Q sky130_fd_sc_hd__dfxtp_1
X_3877_ _3877_/A vssd1 vssd1 vccd1 vccd1 _8371_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3377_ clkbuf_0__3377_/X vssd1 vssd1 vccd1 vccd1 _6906__469/A sky130_fd_sc_hd__clkbuf_4
X_5616_ _5616_/A vssd1 vssd1 vccd1 vccd1 _7821_/D sky130_fd_sc_hd__clkbuf_1
X_5547_ _5547_/A vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__buf_2
X_8335_ _8335_/CLK _8335_/D vssd1 vssd1 vccd1 vccd1 _8335_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__3414_ _7076_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3414_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__3345_ _6780_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3345_/X sky130_fd_sc_hd__clkbuf_16
X_8266_ _8266_/CLK _8266_/D vssd1 vssd1 vccd1 vccd1 _8266_/Q sky130_fd_sc_hd__dfxtp_1
X_5478_ _5478_/A vssd1 vssd1 vccd1 vccd1 _7900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7217_ _6198_/X _7216_/Y _7198_/X _7194_/X _7098_/A vssd1 vssd1 vccd1 vccd1 _7218_/B
+ sky130_fd_sc_hd__o32a_1
X_4429_ _4429_/A vssd1 vssd1 vccd1 vccd1 _8109_/D sky130_fd_sc_hd__clkbuf_1
X_6929__483 _6931__485/A vssd1 vssd1 vccd1 vccd1 _8080_/CLK sky130_fd_sc_hd__inv_2
X_8197_ _8197_/CLK _8197_/D vssd1 vssd1 vccd1 vccd1 _8197_/Q sky130_fd_sc_hd__dfxtp_1
X_7148_ _8227_/Q vssd1 vssd1 vccd1 vccd1 _7151_/A sky130_fd_sc_hd__inv_2
XFILLER_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3593_ clkbuf_0__3593_/X vssd1 vssd1 vccd1 vccd1 _7350__165/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6796__399 _6796__399/A vssd1 vssd1 vccd1 vccd1 _7984_/CLK sky130_fd_sc_hd__inv_2
X_3800_ _7755_/Q _7754_/Q vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__or2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _4703_/X _7806_/Q _7646_/Q _4705_/X _4726_/X vssd1 vssd1 vccd1 vccd1 _4780_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6381_ _6381_/A vssd1 vssd1 vccd1 vccd1 _7745_/D sky130_fd_sc_hd__clkbuf_1
X_5401_ _7933_/Q _4529_/X _5401_/S vssd1 vssd1 vccd1 vccd1 _5402_/A sky130_fd_sc_hd__mux2_1
X_5332_ _5332_/A vssd1 vssd1 vccd1 vccd1 _7968_/D sky130_fd_sc_hd__clkbuf_1
X_8120_ _8120_/CLK _8120_/D vssd1 vssd1 vccd1 vccd1 _8120_/Q sky130_fd_sc_hd__dfxtp_1
X_5263_ _5263_/A vssd1 vssd1 vccd1 vccd1 _7998_/D sky130_fd_sc_hd__clkbuf_1
X_8051_ _8051_/CLK _8051_/D vssd1 vssd1 vccd1 vccd1 _8051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5194_ _8100_/Q _5098_/X _5125_/X _8383_/Q vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__o22a_1
X_4214_ _4214_/A vssd1 vssd1 vccd1 vccd1 _4214_/X sky130_fd_sc_hd__clkbuf_4
X_4145_ _4145_/A vssd1 vssd1 vccd1 vccd1 _8249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4076_ _5743_/A vssd1 vssd1 vccd1 vccd1 _5635_/A sky130_fd_sc_hd__buf_4
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7904_ _7904_/CLK _7904_/D vssd1 vssd1 vccd1 vccd1 _7904_/Q sky130_fd_sc_hd__dfxtp_1
X_7835_ _7835_/CLK _7835_/D vssd1 vssd1 vccd1 vccd1 _7835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _5149_/S vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7766_ _7766_/CLK _7766_/D vssd1 vssd1 vccd1 vccd1 _7766_/Q sky130_fd_sc_hd__dfxtp_1
X_6717_ _6738_/B _6720_/B _8337_/Q vssd1 vssd1 vccd1 vccd1 _7430_/C sky130_fd_sc_hd__a21o_1
X_3929_ _3929_/A vssd1 vssd1 vccd1 vccd1 _8315_/D sky130_fd_sc_hd__clkbuf_1
X_7697_ _7697_/CLK _7697_/D vssd1 vssd1 vccd1 vccd1 _7697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8318_ _8318_/CLK _8318_/D vssd1 vssd1 vccd1 vccd1 _8318_/Q sky130_fd_sc_hd__dfxtp_1
X_6450__233 _6451__234/A vssd1 vssd1 vccd1 vccd1 _7790_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8249_ _8249_/CLK _8249_/D vssd1 vssd1 vccd1 vccd1 _8249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7065__92 _7066__93/A vssd1 vssd1 vccd1 vccd1 _8189_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5950_/A vssd1 vssd1 vccd1 vccd1 _5950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4901_ _4901_/A vssd1 vssd1 vccd1 vccd1 _8035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5881_ _5881_/A vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__clkbuf_1
X_7620_ _7635_/S vssd1 vssd1 vccd1 vccd1 _7627_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4832_ _4757_/A _4822_/X _4825_/X _4831_/X _4549_/A vssd1 vssd1 vccd1 vccd1 _4832_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _4686_/X _4761_/X _4762_/X vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__o21a_1
X_7482_ _7482_/A _7482_/B vssd1 vssd1 vccd1 vccd1 _8342_/D sky130_fd_sc_hd__nor2_1
X_4694_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__buf_2
X_6502_ _6502_/A vssd1 vssd1 vccd1 vccd1 _6502_/X sky130_fd_sc_hd__buf_1
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6364_ _6364_/A vssd1 vssd1 vccd1 vccd1 _7737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5315_ _5284_/X _7975_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5316_/A sky130_fd_sc_hd__mux2_1
X_6514__285 _6514__285/A vssd1 vssd1 vccd1 vccd1 _7842_/CLK sky130_fd_sc_hd__inv_2
X_6295_ _8064_/Q _6231_/X _6287_/X _6244_/X vssd1 vssd1 vccd1 vccd1 _6295_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8103_ _8103_/CLK _8103_/D vssd1 vssd1 vccd1 vccd1 _8103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8034_ _8034_/CLK _8034_/D vssd1 vssd1 vccd1 vccd1 _8034_/Q sky130_fd_sc_hd__dfxtp_1
X_5246_ _8004_/Q _4956_/A _5274_/B _5245_/X _4953_/A vssd1 vssd1 vccd1 vccd1 _5246_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5177_ _8006_/Q _4956_/A _5031_/X _5176_/X _4953_/A vssd1 vssd1 vccd1 vccd1 _5177_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _8363_/Q vssd1 vssd1 vccd1 vccd1 _4128_/X sky130_fd_sc_hd__buf_2
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4059_ _8051_/Q _4059_/B vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7818_ _7818_/CLK _7818_/D vssd1 vssd1 vccd1 vccd1 _7818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7749_ _8348_/CLK _7749_/D vssd1 vssd1 vccd1 vccd1 _7749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6457__239 _6457__239/A vssd1 vssd1 vccd1 vccd1 _7796_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6080_ _6080_/A vssd1 vssd1 vccd1 vccd1 _7644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _5101_/B sky130_fd_sc_hd__nand2_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5031_ _5274_/B vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6982_ _7000_/A vssd1 vssd1 vccd1 vccd1 _6982_/X sky130_fd_sc_hd__buf_1
X_5933_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5942_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5864_ _7598_/B _5866_/B vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__or2_1
X_7603_ _7167_/A _7602_/Y _6246_/X vssd1 vssd1 vccd1 vccd1 _7603_/X sky130_fd_sc_hd__a21o_1
X_4815_ _7789_/Q _4683_/A _4814_/X vssd1 vssd1 vccd1 vccd1 _4819_/B sky130_fd_sc_hd__o21a_1
X_7534_ _7534_/A vssd1 vssd1 vccd1 vccd1 _8359_/D sky130_fd_sc_hd__clkbuf_1
X_5795_ _5795_/A _5795_/B vssd1 vssd1 vccd1 vccd1 _5811_/S sky130_fd_sc_hd__or2_2
X_4746_ _4697_/X _7706_/Q _7655_/Q _4699_/X vssd1 vssd1 vccd1 vccd1 _4746_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_0__3593_ _7345_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3593_/X sky130_fd_sc_hd__clkbuf_16
X_7465_ _7470_/A _7465_/B vssd1 vssd1 vccd1 vccd1 _8335_/D sky130_fd_sc_hd__nor2_1
X_4677_ _7784_/Q _4573_/B _4676_/X vssd1 vssd1 vccd1 vccd1 _4677_/X sky130_fd_sc_hd__a21o_1
X_6416_ _6434_/A vssd1 vssd1 vccd1 vccd1 _6416_/X sky130_fd_sc_hd__buf_1
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6347_ _6309_/A _6237_/A _6144_/A vssd1 vssd1 vccd1 vccd1 _6347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6278_ _8402_/Q _6249_/X _6301_/B _6228_/X vssd1 vssd1 vccd1 vccd1 _6278_/X sky130_fd_sc_hd__a31o_1
X_5229_ _5103_/X _5227_/X _5228_/X vssd1 vssd1 vccd1 vccd1 _5230_/C sky130_fd_sc_hd__o21a_1
X_8017_ _8017_/CLK _8017_/D vssd1 vssd1 vccd1 vccd1 _8017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3413_ clkbuf_0__3413_/X vssd1 vssd1 vccd1 vccd1 _7187_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3344_ clkbuf_0__3344_/X vssd1 vssd1 vccd1 vccd1 _6779__385/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8452__227 vssd1 vssd1 vccd1 vccd1 _8452__227/HI versionID[1] sky130_fd_sc_hd__conb_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6836__417 _6837__418/A vssd1 vssd1 vccd1 vccd1 _8010_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875__444 _6876__445/A vssd1 vssd1 vccd1 vccd1 _8039_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4600_ _4594_/X _4597_/X _4599_/X vssd1 vssd1 vccd1 vccd1 _4600_/X sky130_fd_sc_hd__a21o_1
X_5580_ _5580_/A vssd1 vssd1 vccd1 vccd1 _7835_/D sky130_fd_sc_hd__clkbuf_1
X_4531_ _4531_/A vssd1 vssd1 vccd1 vccd1 _8067_/D sky130_fd_sc_hd__clkbuf_1
X_7250_ _7202_/A _7153_/B _7222_/A _7233_/A _7152_/A vssd1 vssd1 vccd1 vccd1 _7251_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4462_ _3831_/X _8094_/Q _4462_/S vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6201_ _7618_/A vssd1 vssd1 vccd1 vccd1 _6201_/X sky130_fd_sc_hd__clkbuf_2
X_4393_ _8121_/Q _4392_/X _4402_/S vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__mux2_1
X_7181_ _7187_/A vssd1 vssd1 vccd1 vccd1 _7181_/X sky130_fd_sc_hd__buf_1
X_6132_ _6128_/X _7849_/Q _6126_/X _6129_/X _7673_/Q vssd1 vssd1 vccd1 vccd1 _7673_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _7688_/Q _6061_/X _6051_/X _6062_/X vssd1 vssd1 vccd1 vccd1 _6063_/X sky130_fd_sc_hd__o22a_4
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6923__478 _6925__480/A vssd1 vssd1 vccd1 vccd1 _8075_/CLK sky130_fd_sc_hd__inv_2
X_5014_ _5240_/S vssd1 vssd1 vccd1 vccd1 _5204_/S sky130_fd_sc_hd__buf_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7568__41 _7569__42/A vssd1 vssd1 vccd1 vccd1 _8380_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _5916_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__and2_1
XFILLER_81_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6896_ _6896_/A vssd1 vssd1 vccd1 vccd1 _6896_/X sky130_fd_sc_hd__buf_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5847_ _7626_/A _5855_/B vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__or2_1
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5778_ _5778_/A vssd1 vssd1 vccd1 vccd1 _7704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7517_ _8351_/Q _7511_/X _7516_/X _7448_/X vssd1 vssd1 vccd1 vccd1 _8351_/D sky130_fd_sc_hd__o211a_1
X_4729_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7448_ _7493_/A vssd1 vssd1 vccd1 vccd1 _7448_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3189_ clkbuf_0__3189_/X vssd1 vssd1 vccd1 vccd1 _6421__210/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3600_ clkbuf_0__3600_/X vssd1 vssd1 vccd1 vccd1 _7387__20/A sky130_fd_sc_hd__clkbuf_4
X_6750_ _8344_/Q _6757_/D vssd1 vssd1 vccd1 vccd1 _7420_/B sky130_fd_sc_hd__xnor2_4
X_5701_ _7783_/Q _5590_/X _5705_/S vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__mux2_1
X_3962_ _8358_/Q vssd1 vssd1 vccd1 vccd1 _4226_/A sky130_fd_sc_hd__clkbuf_4
X_3893_ _3893_/A _3968_/B vssd1 vssd1 vccd1 vccd1 _3894_/B sky130_fd_sc_hd__nor2_1
X_6681_ _6681_/A vssd1 vssd1 vccd1 vccd1 _6681_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3393_ clkbuf_0__3393_/X vssd1 vssd1 vccd1 vccd1 _6980__525/A sky130_fd_sc_hd__clkbuf_4
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _7814_/D sky130_fd_sc_hd__clkbuf_1
X_8351_ _8407_/CLK _8351_/D vssd1 vssd1 vccd1 vccd1 _8351_/Q sky130_fd_sc_hd__dfxtp_2
X_5563_ _5563_/A vssd1 vssd1 vccd1 vccd1 _7840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4514_ _8363_/Q vssd1 vssd1 vccd1 vccd1 _4514_/X sky130_fd_sc_hd__clkbuf_2
X_7302_ _7320_/A vssd1 vssd1 vccd1 vccd1 _7302_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3361_ _6834_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3361_/X sky130_fd_sc_hd__clkbuf_16
X_8282_ _8282_/CLK _8282_/D vssd1 vssd1 vccd1 vccd1 _8282_/Q sky130_fd_sc_hd__dfxtp_1
X_5494_ _5509_/S vssd1 vssd1 vccd1 vccd1 _5503_/S sky130_fd_sc_hd__buf_4
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7233_ _7233_/A _8222_/Q vssd1 vssd1 vccd1 vccd1 _7233_/X sky130_fd_sc_hd__or2b_1
X_4445_ _4445_/A vssd1 vssd1 vccd1 vccd1 _8102_/D sky130_fd_sc_hd__clkbuf_1
X_7164_ _7599_/A _7164_/B vssd1 vssd1 vccd1 vccd1 _7164_/Y sky130_fd_sc_hd__nand2_1
X_4376_ _4214_/X _8127_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6115_ _6104_/X _7696_/Q _6107_/X _6111_/X _7664_/Q vssd1 vssd1 vccd1 vccd1 _7664_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7110_/C _7129_/A _7150_/B _8219_/Q vssd1 vssd1 vccd1 vccd1 _7221_/B sky130_fd_sc_hd__a31o_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6046_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__and2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _7997_/CLK _7997_/D vssd1 vssd1 vccd1 vccd1 _7997_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6414__204 _6415__205/A vssd1 vssd1 vccd1 vccd1 _7761_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7562__36 _7564__38/A vssd1 vssd1 vccd1 vccd1 _8375_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4230_ _5347_/C _5347_/B _4230_/C vssd1 vssd1 vccd1 vccd1 _5475_/B sky130_fd_sc_hd__nand3_4
X_4161_ _4161_/A vssd1 vssd1 vccd1 vccd1 _8243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4092_ _4092_/A vssd1 vssd1 vccd1 vccd1 _8268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7920_ _7920_/CLK _7920_/D vssd1 vssd1 vccd1 vccd1 _7920_/Q sky130_fd_sc_hd__dfxtp_1
X_7851_ _7854_/CLK _7851_/D vssd1 vssd1 vccd1 vccd1 _7851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6802_ _8352_/Q _6810_/B vssd1 vssd1 vccd1 vccd1 _6803_/A sky130_fd_sc_hd__and2_1
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7782_ _7782_/CLK _7782_/D vssd1 vssd1 vccd1 vccd1 _7782_/Q sky130_fd_sc_hd__dfxtp_1
X_4994_ _5100_/A vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6733_ _7143_/A _7447_/A vssd1 vssd1 vccd1 vccd1 _6733_/Y sky130_fd_sc_hd__nand2_1
X_3945_ _3945_/A vssd1 vssd1 vccd1 vccd1 _8310_/D sky130_fd_sc_hd__clkbuf_1
X_6664_ _6518_/A _6322_/C _6666_/S vssd1 vssd1 vccd1 vccd1 _6665_/A sky130_fd_sc_hd__mux2_1
X_8403_ _8407_/CLK _8403_/D vssd1 vssd1 vccd1 vccd1 _8403_/Q sky130_fd_sc_hd__dfxtp_2
X_3876_ _3875_/X _8371_/Q _3882_/S vssd1 vssd1 vccd1 vccd1 _3877_/A sky130_fd_sc_hd__mux2_1
X_5615_ _5570_/X _7821_/Q _5615_/S vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3376_ clkbuf_0__3376_/X vssd1 vssd1 vccd1 vccd1 _6901__465/A sky130_fd_sc_hd__clkbuf_4
X_6595_ _6601_/A vssd1 vssd1 vccd1 vccd1 _6595_/X sky130_fd_sc_hd__buf_1
XFILLER_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8334_ _8334_/CLK _8334_/D vssd1 vssd1 vccd1 vccd1 _8334_/Q sky130_fd_sc_hd__dfxtp_1
X_6888__454 _6888__454/A vssd1 vssd1 vccd1 vccd1 _8049_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3413_ _7075_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3413_/X sky130_fd_sc_hd__clkbuf_16
X_5546_ _5546_/A vssd1 vssd1 vccd1 vccd1 _7869_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3344_ _6774_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3344_/X sky130_fd_sc_hd__clkbuf_16
X_5477_ _7900_/Q _5025_/A _5485_/S vssd1 vssd1 vccd1 vccd1 _5478_/A sky130_fd_sc_hd__mux2_1
X_8265_ _8265_/CLK _8265_/D vssd1 vssd1 vccd1 vccd1 _8265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7216_ _7216_/A _7216_/B vssd1 vssd1 vccd1 vccd1 _7216_/Y sky130_fd_sc_hd__nand2_1
X_4428_ _8109_/Q _4404_/X _4432_/S vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__mux2_1
X_8196_ _8196_/CLK _8196_/D vssd1 vssd1 vccd1 vccd1 _8196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7147_ _8228_/Q vssd1 vssd1 vccd1 vccd1 _7152_/A sky130_fd_sc_hd__inv_2
XFILLER_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4359_ _4359_/A vssd1 vssd1 vccd1 vccd1 _8135_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3592_ clkbuf_0__3592_/X vssd1 vssd1 vccd1 vccd1 _7344__160/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i _7717_/CLK vssd1 vssd1 vccd1 vccd1 _7846_/CLK sky130_fd_sc_hd__clkbuf_16
X_6029_ _7729_/Q input11/X _6029_/S vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6639__341 _6641__343/A vssd1 vssd1 vccd1 vccd1 _7922_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6380_ _7852_/Q _7745_/Q _6382_/S vssd1 vssd1 vccd1 vccd1 _6381_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5400_ _5400_/A vssd1 vssd1 vccd1 vccd1 _7934_/D sky130_fd_sc_hd__clkbuf_1
X_5331_ _5278_/X _7968_/Q _5339_/S vssd1 vssd1 vccd1 vccd1 _5332_/A sky130_fd_sc_hd__mux2_1
X_8050_ _8050_/CLK _8050_/D vssd1 vssd1 vccd1 vccd1 _8050_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5262_ _5262_/A _7547_/A _5262_/C vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__and3_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5193_ _8322_/Q _8068_/Q _5207_/S vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__mux2_1
X_4213_ _4213_/A vssd1 vssd1 vccd1 vccd1 _8192_/D sky130_fd_sc_hd__clkbuf_1
X_4144_ _8249_/Q _4143_/X _4144_/S vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4075_ _4843_/A _4324_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _5743_/A sky130_fd_sc_hd__or3_4
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7903_ _7903_/CLK _7903_/D vssd1 vssd1 vccd1 vccd1 _7903_/Q sky130_fd_sc_hd__dfxtp_1
X_7834_ _7834_/CLK _7834_/D vssd1 vssd1 vccd1 vccd1 _7834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7765_ _7765_/CLK _7765_/D vssd1 vssd1 vccd1 vccd1 _7765_/Q sky130_fd_sc_hd__dfxtp_1
X_6716_ _6716_/A vssd1 vssd1 vccd1 vccd1 _7430_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4977_ _5240_/S vssd1 vssd1 vccd1 vccd1 _5149_/S sky130_fd_sc_hd__buf_4
X_3928_ _3884_/X _8315_/Q _3932_/S vssd1 vssd1 vccd1 vccd1 _3929_/A sky130_fd_sc_hd__mux2_1
X_7696_ _7697_/CLK _7696_/D vssd1 vssd1 vccd1 vccd1 _7696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3859_ _3859_/A vssd1 vssd1 vccd1 vccd1 _8376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3359_ clkbuf_0__3359_/X vssd1 vssd1 vccd1 vccd1 _6827__410/A sky130_fd_sc_hd__clkbuf_4
X_8317_ _8317_/CLK _8317_/D vssd1 vssd1 vccd1 vccd1 _8317_/Q sky130_fd_sc_hd__dfxtp_1
X_5529_ _5761_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _5545_/S sky130_fd_sc_hd__or2_2
X_8248_ _8248_/CLK _8248_/D vssd1 vssd1 vccd1 vccd1 _8248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8179_ _8179_/CLK _8179_/D vssd1 vssd1 vccd1 vccd1 _8179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3189_ _6416_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3189_/X sky130_fd_sc_hd__clkbuf_16
X_6977__522 _6977__522/A vssd1 vssd1 vccd1 vccd1 _8119_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8420__195 vssd1 vssd1 vccd1 vccd1 _8420__195/HI core0Index[2] sky130_fd_sc_hd__conb_1
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5880_ _5880_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__or2_1
X_4900_ _8035_/Q _4395_/X _4904_/S vssd1 vssd1 vccd1 vccd1 _4901_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4831_ _4664_/A _4827_/X _4830_/X _4575_/X vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7550_ _7550_/A vssd1 vssd1 vccd1 vccd1 _8365_/D sky130_fd_sc_hd__clkbuf_1
X_4762_ _8109_/Q _4724_/X _4725_/X _8085_/Q _4726_/X vssd1 vssd1 vccd1 vccd1 _4762_/X
+ sky130_fd_sc_hd__o221a_1
X_7481_ _8342_/Q _7466_/X _7474_/X _6699_/B vssd1 vssd1 vccd1 vccd1 _7482_/B sky130_fd_sc_hd__o2bb2a_1
X_4693_ _8198_/Q _4681_/X _4686_/X _4692_/X vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6363_ _5920_/A _7737_/Q _6371_/S vssd1 vssd1 vccd1 vccd1 _6364_/A sky130_fd_sc_hd__mux2_1
X_8102_ _8102_/CLK _8102_/D vssd1 vssd1 vccd1 vccd1 _8102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5314_ _5314_/A vssd1 vssd1 vccd1 vccd1 _7976_/D sky130_fd_sc_hd__clkbuf_1
X_6294_ _8400_/Q vssd1 vssd1 vccd1 vccd1 _7621_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8033_ _8033_/CLK _8033_/D vssd1 vssd1 vccd1 vccd1 _8033_/Q sky130_fd_sc_hd__dfxtp_1
X_5245_ _5265_/B _5223_/X _5230_/X _5244_/X vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5176_ _5265_/B _5154_/X _5161_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_1_0_0__3360_ clkbuf_0__3360_/X vssd1 vssd1 vccd1 vccd1 _6830__412/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4127_ _4127_/A vssd1 vssd1 vccd1 vccd1 _8255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4058_ _8053_/Q _8048_/Q vssd1 vssd1 vccd1 vccd1 _4536_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7817_ _7817_/CLK _7817_/D vssd1 vssd1 vccd1 vccd1 _7817_/Q sky130_fd_sc_hd__dfxtp_1
X_7748_ _8348_/CLK _7748_/D vssd1 vssd1 vccd1 vccd1 _7748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7679_ _8348_/CLK _7679_/D vssd1 vssd1 vccd1 vccd1 _7679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6576__291 _6577__292/A vssd1 vssd1 vccd1 vccd1 _7872_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5274_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6981_ _6981_/A vssd1 vssd1 vccd1 vccd1 _6981_/X sky130_fd_sc_hd__buf_1
X_5932_ _5932_/A vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5863_/A vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7602_ _7602_/A vssd1 vssd1 vccd1 vccd1 _7602_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5794_ _5794_/A vssd1 vssd1 vccd1 vccd1 _7653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4814_ _8115_/Q _4705_/A _4750_/A _4813_/X _4642_/A vssd1 vssd1 vccd1 vccd1 _4814_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7533_ _7533_/A _7533_/B _7547_/B vssd1 vssd1 vccd1 vccd1 _7534_/A sky130_fd_sc_hd__and3_1
X_4745_ _8197_/Q _4681_/X _4715_/X _4744_/X vssd1 vssd1 vccd1 vccd1 _4745_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3592_ _7339_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3592_/X sky130_fd_sc_hd__clkbuf_16
X_7464_ _8335_/Q _7458_/X _7461_/X _7432_/B vssd1 vssd1 vccd1 vccd1 _7465_/B sky130_fd_sc_hd__o2bb2a_1
X_4676_ _4676_/A vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7395_ _7561_/A vssd1 vssd1 vccd1 vccd1 _7395_/X sky130_fd_sc_hd__buf_1
X_6346_ _7170_/A _6346_/B _7547_/B vssd1 vssd1 vccd1 vccd1 _6405_/B sky130_fd_sc_hd__nand3_1
XFILLER_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6277_ _7716_/Q _6216_/X _6276_/X vssd1 vssd1 vccd1 vccd1 _7716_/D sky130_fd_sc_hd__a21o_1
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8016_ _8016_/CLK _8016_/D vssd1 vssd1 vccd1 vccd1 _8016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5228_ _8155_/Q _5187_/A _5151_/X _8147_/Q _5009_/A vssd1 vssd1 vccd1 vccd1 _5228_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0_0__3412_ clkbuf_0__3412_/X vssd1 vssd1 vccd1 vccd1 _7073__99/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5159_ _8157_/Q _5187_/A _5151_/X _8149_/Q _5009_/A vssd1 vssd1 vccd1 vccd1 _5159_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0_0__3343_ clkbuf_0__3343_/X vssd1 vssd1 vccd1 vccd1 _6772__379/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6463__244 _6464__245/A vssd1 vssd1 vccd1 vccd1 _7801_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4530_ _8067_/Q _4529_/X _4530_/S vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__mux2_1
X_6103__191 _6103__191/A vssd1 vssd1 vccd1 vccd1 _7660_/CLK sky130_fd_sc_hd__inv_2
X_4461_ _4461_/A vssd1 vssd1 vccd1 vccd1 _8095_/D sky130_fd_sc_hd__clkbuf_1
X_6200_ _6249_/A _6236_/A vssd1 vssd1 vccd1 vccd1 _7618_/A sky130_fd_sc_hd__and2_1
X_7180_ _7262_/B _7174_/C _7179_/Y vssd1 vssd1 vccd1 vccd1 _8204_/D sky130_fd_sc_hd__a21oi_1
XFILLER_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6131_ _6128_/X _7848_/Q _6126_/X _6129_/X _7672_/Q vssd1 vssd1 vccd1 vccd1 _7672_/D
+ sky130_fd_sc_hd__o32a_1
X_4392_ _7991_/Q vssd1 vssd1 vccd1 vccd1 _4392_/X sky130_fd_sc_hd__buf_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6062_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__and2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5009_/X _5011_/X _5119_/A vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__a21o_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5915_ _5915_/A vssd1 vssd1 vccd1 vccd1 _5915_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5846_ _5903_/B vssd1 vssd1 vccd1 vccd1 _5855_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5777_ _5570_/X _7704_/Q _5777_/S vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__mux2_1
X_7516_ _8352_/Q _7523_/B _7513_/X vssd1 vssd1 vccd1 vccd1 _7516_/X sky130_fd_sc_hd__or3b_1
X_6672__363 _6674__365/A vssd1 vssd1 vccd1 vccd1 _7947_/CLK sky130_fd_sc_hd__inv_2
X_4728_ _4686_/X _4723_/X _4727_/X vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4659_ _7973_/Q _7965_/Q _7769_/Q _8034_/Q _4579_/X _4580_/X vssd1 vssd1 vccd1 vccd1
+ _4659_/X sky130_fd_sc_hd__mux4_1
X_7447_ _7447_/A _7447_/B vssd1 vssd1 vccd1 vccd1 _7447_/Y sky130_fd_sc_hd__nand2_1
X_8412__234 vssd1 vssd1 vccd1 vccd1 partID[6] _8412__234/LO sky130_fd_sc_hd__conb_1
X_6633__336 _6635__338/A vssd1 vssd1 vccd1 vccd1 _7917_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6329_ _7596_/A _6337_/B _6332_/C _6337_/D vssd1 vssd1 vccd1 vccd1 _6329_/X sky130_fd_sc_hd__and4_1
XFILLER_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3188_ clkbuf_0__3188_/X vssd1 vssd1 vccd1 vccd1 _6413__203/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8235_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _8306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5700_ _5700_/A vssd1 vssd1 vccd1 vccd1 _7784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3892_ _3892_/A vssd1 vssd1 vccd1 vccd1 _8366_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3392_ clkbuf_0__3392_/X vssd1 vssd1 vccd1 vccd1 _6971__517/A sky130_fd_sc_hd__clkbuf_4
X_5631_ _5567_/X _7814_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8350_ _8407_/CLK _8350_/D vssd1 vssd1 vccd1 vccd1 _8350_/Q sky130_fd_sc_hd__dfxtp_1
X_5562_ _5561_/X _7840_/Q _5562_/S vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3360_ _6828_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3360_/X sky130_fd_sc_hd__clkbuf_16
X_8281_ _8281_/CLK _8281_/D vssd1 vssd1 vccd1 vccd1 _8281_/Q sky130_fd_sc_hd__dfxtp_1
X_4513_ _4513_/A vssd1 vssd1 vccd1 vccd1 _8073_/D sky130_fd_sc_hd__clkbuf_1
X_7301_ _7332_/A vssd1 vssd1 vccd1 vccd1 _7301_/X sky130_fd_sc_hd__buf_1
X_7232_ _7244_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _8221_/D sky130_fd_sc_hd__nor2_1
X_5493_ _5761_/A _5671_/B vssd1 vssd1 vccd1 vccd1 _5509_/S sky130_fd_sc_hd__or2_2
X_7307__130 _7307__130/A vssd1 vssd1 vccd1 vccd1 _8257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4444_ _4217_/X _8102_/Q _4444_/S vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__mux2_1
X_7163_ _8394_/Q _7164_/B _7161_/X _7162_/Y vssd1 vssd1 vccd1 vccd1 _7163_/X sky130_fd_sc_hd__o22a_1
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _8128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7094_ _8216_/Q _8215_/Q _8214_/Q _8213_/Q vssd1 vssd1 vccd1 vccd1 _7150_/B sky130_fd_sc_hd__and4_1
X_6114_ _6104_/X _7695_/Q _6107_/X _6111_/X _7663_/Q vssd1 vssd1 vccd1 vccd1 _7663_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _7681_/Q _6032_/X _6039_/X _6044_/X vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__o22a_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7996_ _7996_/CLK _7996_/D vssd1 vssd1 vccd1 vccd1 _7996_/Q sky130_fd_sc_hd__dfxtp_2
X_6971__517 _6971__517/A vssd1 vssd1 vccd1 vccd1 _8114_/CLK sky130_fd_sc_hd__inv_2
X_5829_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5909_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7374__9 _7374__9/A vssd1 vssd1 vccd1 vccd1 _8311_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6679__369 _6680__370/A vssd1 vssd1 vccd1 vccd1 _7953_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4160_ _8243_/Q _4093_/X _4164_/S vssd1 vssd1 vccd1 vccd1 _4161_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4091_ _8268_/Q _4090_/X _4091_/S vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7850_ _7991_/CLK _7850_/D vssd1 vssd1 vccd1 vccd1 _7850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6801_ _6801_/A vssd1 vssd1 vccd1 vccd1 _6810_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3513_ clkbuf_0__3513_/X vssd1 vssd1 vccd1 vccd1 _7190__113/A sky130_fd_sc_hd__clkbuf_4
X_7781_ _7781_/CLK _7781_/D vssd1 vssd1 vccd1 vccd1 _7781_/Q sky130_fd_sc_hd__dfxtp_1
X_4993_ _5171_/S vssd1 vssd1 vccd1 vccd1 _5227_/S sky130_fd_sc_hd__buf_4
X_6732_ _8331_/Q vssd1 vssd1 vccd1 vccd1 _7447_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3944_ _8310_/Q _3943_/X _3952_/S vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__mux2_1
X_6663_ _6663_/A vssd1 vssd1 vccd1 vccd1 _7941_/D sky130_fd_sc_hd__clkbuf_1
X_3875_ _8363_/Q vssd1 vssd1 vccd1 vccd1 _3875_/X sky130_fd_sc_hd__clkbuf_4
X_8402_ _8407_/CLK _8402_/D vssd1 vssd1 vccd1 vccd1 _8402_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_1_0__3375_ clkbuf_0__3375_/X vssd1 vssd1 vccd1 vccd1 _6893__458/A sky130_fd_sc_hd__clkbuf_4
X_5614_ _5614_/A vssd1 vssd1 vccd1 vccd1 _7822_/D sky130_fd_sc_hd__clkbuf_1
X_6476__254 _6477__255/A vssd1 vssd1 vccd1 vccd1 _7811_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3412_ _7069_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3412_/X sky130_fd_sc_hd__clkbuf_16
X_8333_ _8334_/CLK _8333_/D vssd1 vssd1 vccd1 vccd1 _8333_/Q sky130_fd_sc_hd__dfxtp_1
X_5545_ _5308_/X _7869_/Q _5545_/S vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3343_ _6768_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3343_/X sky130_fd_sc_hd__clkbuf_16
X_8264_ _8264_/CLK _8264_/D vssd1 vssd1 vccd1 vccd1 _8264_/Q sky130_fd_sc_hd__dfxtp_1
X_5476_ _5491_/S vssd1 vssd1 vccd1 vccd1 _5485_/S sky130_fd_sc_hd__buf_2
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7215_ _7218_/A _7215_/B vssd1 vssd1 vccd1 vccd1 _8217_/D sky130_fd_sc_hd__nor2_1
X_8195_ _8195_/CLK _8195_/D vssd1 vssd1 vccd1 vccd1 _8195_/Q sky130_fd_sc_hd__dfxtp_1
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _8110_/D sky130_fd_sc_hd__clkbuf_1
X_7146_ _7104_/X _7146_/B _7146_/C _7146_/D vssd1 vssd1 vccd1 vccd1 _7173_/B sky130_fd_sc_hd__and4b_1
XFILLER_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4358_ _8135_/Q _4131_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4359_/A sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3591_ clkbuf_0__3591_/X vssd1 vssd1 vccd1 vccd1 _7336__153/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4249_/X _8162_/Q _4297_/S vssd1 vssd1 vccd1 vccd1 _4290_/A sky130_fd_sc_hd__mux2_1
X_6028_ _6028_/A vssd1 vssd1 vccd1 vccd1 _6028_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7979_ _7979_/CLK _7979_/D vssd1 vssd1 vccd1 vccd1 _7979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936__489 _6936__489/A vssd1 vssd1 vccd1 vccd1 _8086_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8425__200 vssd1 vssd1 vccd1 vccd1 _8425__200/HI core0Index[7] sky130_fd_sc_hd__conb_1
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5345_/S vssd1 vssd1 vccd1 vccd1 _5339_/S sky130_fd_sc_hd__clkbuf_4
X_5261_ _5261_/A _5261_/B vssd1 vssd1 vccd1 vccd1 _5262_/C sky130_fd_sc_hd__or2_1
XFILLER_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4212_ _4211_/X _8192_/Q _4218_/S vssd1 vssd1 vccd1 vccd1 _4213_/A sky130_fd_sc_hd__mux2_1
X_7000_ _7000_/A vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__buf_1
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5192_ _8314_/Q _5187_/X _5183_/X _8306_/Q _4976_/X vssd1 vssd1 vccd1 vccd1 _5192_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4143_ _8358_/Q vssd1 vssd1 vccd1 vccd1 _4143_/X sky130_fd_sc_hd__clkbuf_2
X_4074_ _4844_/A _4843_/C vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7902_ _7902_/CLK _7902_/D vssd1 vssd1 vccd1 vccd1 _7902_/Q sky130_fd_sc_hd__dfxtp_1
X_7833_ _7833_/CLK _7833_/D vssd1 vssd1 vccd1 vccd1 _7833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7764_ _7764_/CLK _7764_/D vssd1 vssd1 vccd1 vccd1 _7764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6715_ _8399_/Q _7411_/A _7411_/B vssd1 vssd1 vccd1 vccd1 _6742_/C sky130_fd_sc_hd__nand3b_1
X_4976_ _5123_/S vssd1 vssd1 vccd1 vccd1 _4976_/X sky130_fd_sc_hd__buf_2
X_3927_ _3927_/A vssd1 vssd1 vccd1 vccd1 _8316_/D sky130_fd_sc_hd__clkbuf_1
X_7695_ _7697_/CLK _7695_/D vssd1 vssd1 vccd1 vccd1 _7695_/Q sky130_fd_sc_hd__dfxtp_1
X_3858_ _8376_/Q _3834_/X _3862_/S vssd1 vssd1 vccd1 vccd1 _3859_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3358_ clkbuf_0__3358_/X vssd1 vssd1 vccd1 vccd1 _6821__405/A sky130_fd_sc_hd__clkbuf_4
X_3789_ _8001_/Q _7996_/Q vssd1 vssd1 vccd1 vccd1 _4950_/C sky130_fd_sc_hd__xnor2_2
X_8316_ _8316_/CLK _8316_/D vssd1 vssd1 vccd1 vccd1 _8316_/Q sky130_fd_sc_hd__dfxtp_1
X_5528_ _5528_/A vssd1 vssd1 vccd1 vccd1 _7877_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8247_ _8247_/CLK _8247_/D vssd1 vssd1 vccd1 vccd1 _8247_/Q sky130_fd_sc_hd__dfxtp_1
X_5459_ _7908_/Q _5366_/X _5467_/S vssd1 vssd1 vccd1 vccd1 _5460_/A sky130_fd_sc_hd__mux2_1
X_8178_ _8178_/CLK _8178_/D vssd1 vssd1 vccd1 vccd1 _8178_/Q sky130_fd_sc_hd__dfxtp_1
X_7129_ _7129_/A _7159_/A vssd1 vssd1 vccd1 vccd1 _7130_/B sky130_fd_sc_hd__xnor2_2
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3188_ _6410_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3188_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6903__466 _6912__470/A vssd1 vssd1 vccd1 vccd1 _8061_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6984__527 _6985__528/A vssd1 vssd1 vccd1 vccd1 _8124_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6427__215 _6427__215/A vssd1 vssd1 vccd1 vccd1 _7772_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_0_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4830_ _4715_/A _4828_/X _4829_/X vssd1 vssd1 vccd1 vccd1 _4830_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7071__97 _7071__97/A vssd1 vssd1 vccd1 vccd1 _8194_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4761_ _8077_/Q _4691_/X _4687_/X _8040_/Q vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7480_ _7482_/A _7480_/B vssd1 vssd1 vccd1 vccd1 _8341_/D sky130_fd_sc_hd__nor2_1
X_4692_ _4687_/X _7816_/Q _7800_/Q _4691_/X vssd1 vssd1 vccd1 vccd1 _4692_/X sky130_fd_sc_hd__a22o_1
X_6362_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6371_/S sky130_fd_sc_hd__buf_2
XFILLER_115_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5313_ _5278_/X _7976_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5314_/A sky130_fd_sc_hd__mux2_1
X_8101_ _8101_/CLK _8101_/D vssd1 vssd1 vccd1 vccd1 _8101_/Q sky130_fd_sc_hd__dfxtp_1
X_6293_ _6221_/X _6290_/X _6291_/X _6292_/X vssd1 vssd1 vccd1 vccd1 _7718_/D sky130_fd_sc_hd__a211o_1
X_8032_ _8032_/CLK _8032_/D vssd1 vssd1 vccd1 vccd1 _8032_/Q sky130_fd_sc_hd__dfxtp_1
X_5244_ _5124_/A _5233_/X _5236_/X _5243_/X _5002_/A vssd1 vssd1 vccd1 vccd1 _5244_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_29_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5175_ _5124_/A _5164_/X _5167_/X _5002_/A _5174_/X vssd1 vssd1 vccd1 vccd1 _5175_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4126_ _8255_/Q _4125_/X _4135_/S vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4057_ _4843_/B _4731_/A _4056_/Y vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__or3b_1
XFILLER_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6779__385 _6779__385/A vssd1 vssd1 vccd1 vccd1 _7970_/CLK sky130_fd_sc_hd__inv_2
X_7816_ _7816_/CLK _7816_/D vssd1 vssd1 vccd1 vccd1 _7816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7747_ _7747_/CLK _7747_/D vssd1 vssd1 vccd1 vccd1 _7747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4959_ _7994_/Q vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__clkbuf_2
X_7678_ _7747_/CLK _7678_/D vssd1 vssd1 vccd1 vccd1 _7678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7005__545 _7005__545/A vssd1 vssd1 vccd1 vccd1 _8142_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6095__185 _6095__185/A vssd1 vssd1 vccd1 vccd1 _7654_/CLK sky130_fd_sc_hd__inv_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5931_ _5931_/A _5931_/B vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__and2_1
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5862_ _5862_/A _5866_/B vssd1 vssd1 vccd1 vccd1 _5863_/A sky130_fd_sc_hd__or2_1
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7601_ _7590_/X _7598_/Y _7599_/Y _7600_/X vssd1 vssd1 vccd1 vccd1 _8394_/D sky130_fd_sc_hd__a211oi_1
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5793_ _7653_/Q _5570_/A _5793_/S vssd1 vssd1 vccd1 vccd1 _5794_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4813_ _4696_/A _7885_/Q _7829_/Q _4698_/A vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__a22o_1
X_7532_ _7532_/A vssd1 vssd1 vccd1 vccd1 _8358_/D sky130_fd_sc_hd__clkbuf_1
X_4744_ _4717_/X _7815_/Q _7799_/Q _4691_/X vssd1 vssd1 vccd1 vccd1 _4744_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_0__3591_ _7333_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3591_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7463_ _7470_/A _7463_/B vssd1 vssd1 vccd1 vccd1 _8334_/D sky130_fd_sc_hd__nor2_1
X_4675_ _4675_/A vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__clkbuf_2
X_7394_ _7394_/A vssd1 vssd1 vccd1 vccd1 _7394_/X sky130_fd_sc_hd__buf_1
X_6345_ _7540_/B _6345_/B vssd1 vssd1 vccd1 vccd1 _7547_/B sky130_fd_sc_hd__nor2_2
XFILLER_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6276_ _6270_/A _6273_/X _6275_/X _6246_/X vssd1 vssd1 vccd1 vccd1 _6276_/X sky130_fd_sc_hd__a31o_1
XFILLER_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8015_ _8015_/CLK _8015_/D vssd1 vssd1 vccd1 vccd1 _8015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5227_ _8123_/Q _8131_/Q _5227_/S vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _7068__95/A sky130_fd_sc_hd__clkbuf_4
X_5158_ _8125_/Q _8133_/Q _5227_/S vssd1 vssd1 vccd1 vccd1 _5158_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3342_ clkbuf_0__3342_/X vssd1 vssd1 vccd1 vccd1 _6786_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5089_ _5087_/X _5088_/X _5089_/S vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__mux2_2
X_4109_ _4109_/A vssd1 vssd1 vccd1 vccd1 _8262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7356__170 _7356__170/A vssd1 vssd1 vccd1 vccd1 _8297_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6207__194 _6208__195/A vssd1 vssd1 vccd1 vccd1 _7706_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _3828_/X _8095_/Q _4462_/S vssd1 vssd1 vccd1 vccd1 _4461_/A sky130_fd_sc_hd__mux2_1
X_4391_ _4391_/A vssd1 vssd1 vccd1 vccd1 _8122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6130_ _6128_/X _7847_/Q _6126_/X _6129_/X _7671_/Q vssd1 vssd1 vccd1 vccd1 _7671_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7299__124 _7300__125/A vssd1 vssd1 vccd1 vccd1 _8251_/CLK sky130_fd_sc_hd__inv_2
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6061_ _6079_/D vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__buf_2
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5243_/A vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6963_ _6975_/A vssd1 vssd1 vccd1 vccd1 _6963_/X sky130_fd_sc_hd__buf_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7017__53 _7019__55/A vssd1 vssd1 vccd1 vccd1 _8150_/CLK sky130_fd_sc_hd__inv_2
X_5914_ _5914_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__and2_1
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5845_ _5845_/A vssd1 vssd1 vccd1 vccd1 _5845_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5776_ _5776_/A vssd1 vssd1 vccd1 vccd1 _7705_/D sky130_fd_sc_hd__clkbuf_1
X_7515_ _8350_/Q _7511_/X _7514_/X _7448_/X vssd1 vssd1 vccd1 vccd1 _8350_/D sky130_fd_sc_hd__o211a_1
X_4727_ _8110_/Q _4724_/X _4725_/X _8086_/Q _4726_/X vssd1 vssd1 vccd1 vccd1 _4727_/X
+ sky130_fd_sc_hd__o221a_1
X_7446_ _7489_/A _7513_/A _7439_/C vssd1 vssd1 vccd1 vccd1 _7446_/Y sky130_fd_sc_hd__o21ai_4
X_4658_ _4867_/B _4655_/X _4657_/X vssd1 vssd1 vccd1 vccd1 _4658_/X sky130_fd_sc_hd__a21o_1
Xinput90 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _6349_/C sky130_fd_sc_hd__buf_8
X_4589_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4589_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6328_ _8393_/Q vssd1 vssd1 vccd1 vccd1 _7596_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6259_ _8405_/Q vssd1 vssd1 vccd1 vccd1 _7422_/A sky130_fd_sc_hd__buf_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3256_ clkbuf_0__3256_/X vssd1 vssd1 vccd1 vccd1 _6661__359/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3187_ clkbuf_0__3187_/X vssd1 vssd1 vccd1 vccd1 _6434_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7574__46 _7574__46/A vssd1 vssd1 vccd1 vccd1 _8385_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ _8306_/Q _3959_/X _3964_/S vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _3890_/X _8366_/Q _3891_/S vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3391_ clkbuf_0__3391_/X vssd1 vssd1 vccd1 vccd1 _6968__515/A sky130_fd_sc_hd__clkbuf_4
X_5630_ _5630_/A vssd1 vssd1 vccd1 vccd1 _7815_/D sky130_fd_sc_hd__clkbuf_1
X_5561_ _5561_/A vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4512_ _8073_/Q _4511_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4513_/A sky130_fd_sc_hd__mux2_1
X_8280_ _8280_/CLK _8280_/D vssd1 vssd1 vccd1 vccd1 _8280_/Q sky130_fd_sc_hd__dfxtp_1
X_5492_ _5492_/A vssd1 vssd1 vccd1 vccd1 _7893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7231_ _7220_/X _7230_/Y _7222_/X _7223_/X _7125_/A vssd1 vssd1 vccd1 vccd1 _7232_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4443_ _4443_/A vssd1 vssd1 vccd1 vccd1 _8103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7162_ _7226_/A _7226_/B _7621_/A vssd1 vssd1 vccd1 vccd1 _7162_/Y sky130_fd_sc_hd__a21oi_1
X_4374_ _4211_/X _8128_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7093_ _8217_/Q vssd1 vssd1 vccd1 vccd1 _7129_/A sky130_fd_sc_hd__clkbuf_2
X_6113_ _6104_/X _7694_/Q _6107_/X _6111_/X _7662_/Q vssd1 vssd1 vccd1 vccd1 _7662_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6044_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6044_/X sky130_fd_sc_hd__and2_1
XFILLER_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8442__217 vssd1 vssd1 vccd1 vccd1 _8442__217/HI manufacturerID[9] sky130_fd_sc_hd__conb_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7995_ _7995_/CLK _7995_/D vssd1 vssd1 vccd1 vccd1 _7995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6858__430 _6858__430/A vssd1 vssd1 vccd1 vccd1 _8025_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6819__403 _6820__404/A vssd1 vssd1 vccd1 vccd1 _7996_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6877_ _6877_/A vssd1 vssd1 vccd1 vccd1 _6877_/X sky130_fd_sc_hd__buf_1
XFILLER_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5828_ _5955_/A vssd1 vssd1 vccd1 vccd1 _5944_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0__3589_ clkbuf_0__3589_/X vssd1 vssd1 vccd1 vccd1 _7329__148/A sky130_fd_sc_hd__clkbuf_4
X_5759_ _7757_/Q _5570_/A _5759_/S vssd1 vssd1 vccd1 vccd1 _5760_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7429_ _7429_/A _7429_/B vssd1 vssd1 vccd1 vccd1 _7429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3239_ clkbuf_0__3239_/X vssd1 vssd1 vccd1 vccd1 _6577__292/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _7988_/Q vssd1 vssd1 vccd1 vccd1 _4090_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _6800_/A vssd1 vssd1 vccd1 vccd1 _7986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7780_ _7780_/CLK _7780_/D vssd1 vssd1 vccd1 vccd1 _7780_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3512_ clkbuf_0__3512_/X vssd1 vssd1 vccd1 vccd1 _7186__110/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4992_ _5237_/S vssd1 vssd1 vccd1 vccd1 _5171_/S sky130_fd_sc_hd__buf_2
X_6731_ _7421_/A _7425_/A vssd1 vssd1 vccd1 vccd1 _6731_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3943_ _4211_/A vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__clkbuf_2
X_6662_ _6164_/A _6249_/X _6666_/S vssd1 vssd1 vccd1 vccd1 _6663_/A sky130_fd_sc_hd__mux2_1
X_3874_ _3874_/A vssd1 vssd1 vccd1 vccd1 _8372_/D sky130_fd_sc_hd__clkbuf_1
X_8401_ _8407_/CLK _8401_/D vssd1 vssd1 vccd1 vccd1 _8401_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3374_ clkbuf_0__3374_/X vssd1 vssd1 vccd1 vccd1 _6889__455/A sky130_fd_sc_hd__clkbuf_4
X_5613_ _5567_/X _7822_/Q _5615_/S vssd1 vssd1 vccd1 vccd1 _5614_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8332_ _8332_/CLK _8332_/D vssd1 vssd1 vccd1 vccd1 _8332_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3411_ _7063_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3411_/X sky130_fd_sc_hd__clkbuf_16
X_5544_ _5544_/A vssd1 vssd1 vccd1 vccd1 _7870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3342_ _6767_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3342_/X sky130_fd_sc_hd__clkbuf_16
X_5475_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5491_/S sky130_fd_sc_hd__nor2_2
X_8263_ _8263_/CLK _8263_/D vssd1 vssd1 vccd1 vccd1 _8263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7214_ _6198_/X _7130_/B _7198_/X _7194_/X _7098_/B vssd1 vssd1 vccd1 vccd1 _7215_/B
+ sky130_fd_sc_hd__o32a_1
X_8194_ _8194_/CLK _8194_/D vssd1 vssd1 vccd1 vccd1 _8194_/Q sky130_fd_sc_hd__dfxtp_1
X_4426_ _8110_/Q _4401_/X _4426_/S vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7145_ _7127_/Y _7128_/X _7130_/X _7135_/X _7144_/X vssd1 vssd1 vccd1 vccd1 _7146_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4357_ _4357_/A vssd1 vssd1 vccd1 vccd1 _8136_/D sky130_fd_sc_hd__clkbuf_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3590_ clkbuf_0__3590_/X vssd1 vssd1 vccd1 vccd1 _7339_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4303_/S vssd1 vssd1 vccd1 vccd1 _4297_/S sky130_fd_sc_hd__clkbuf_4
X_7076_ _7187_/A vssd1 vssd1 vccd1 vccd1 _7076_/X sky130_fd_sc_hd__buf_1
X_6027_ _7677_/Q _6025_/X _7608_/A vssd1 vssd1 vccd1 vccd1 _6028_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7978_ _7978_/CLK _7978_/D vssd1 vssd1 vccd1 vccd1 _7978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6685__374 _6686__375/A vssd1 vssd1 vccd1 vccd1 _7958_/CLK sky130_fd_sc_hd__inv_2
X_6646__347 _6647__348/A vssd1 vssd1 vccd1 vccd1 _7928_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _5260_/A vssd1 vssd1 vccd1 vccd1 _7999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4211_ _4211_/A vssd1 vssd1 vccd1 vccd1 _4211_/X sky130_fd_sc_hd__clkbuf_4
X_5191_ _5191_/A _5191_/B vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__or2_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4142_ _4142_/A vssd1 vssd1 vccd1 vccd1 _8250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4073_ _8065_/Q _6253_/A vssd1 vssd1 vccd1 vccd1 _4843_/C sky130_fd_sc_hd__and2_1
XFILLER_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7901_ _7901_/CLK _7901_/D vssd1 vssd1 vccd1 vccd1 _7901_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8359_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7832_ _7832_/CLK _7832_/D vssd1 vssd1 vccd1 vccd1 _7832_/Q sky130_fd_sc_hd__dfxtp_1
X_7763_ _7763_/CLK _7763_/D vssd1 vssd1 vccd1 vccd1 _7763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4975_ _4987_/A vssd1 vssd1 vccd1 vccd1 _5123_/S sky130_fd_sc_hd__clkbuf_4
X_7350__165 _7350__165/A vssd1 vssd1 vccd1 vccd1 _8292_/CLK sky130_fd_sc_hd__inv_2
X_6714_ _7621_/A _6714_/B vssd1 vssd1 vccd1 vccd1 _6742_/B sky130_fd_sc_hd__nand2_1
X_3926_ _3881_/X _8316_/Q _3926_/S vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__mux2_1
X_7694_ _7697_/CLK _7694_/D vssd1 vssd1 vccd1 vccd1 _7694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3857_ _3857_/A vssd1 vssd1 vccd1 vccd1 _8377_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3357_ clkbuf_0__3357_/X vssd1 vssd1 vccd1 vccd1 _6834_/A sky130_fd_sc_hd__clkbuf_4
X_3788_ _8000_/Q _7995_/Q vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__xor2_1
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8315_ _8315_/CLK _8315_/D vssd1 vssd1 vccd1 vccd1 _8315_/Q sky130_fd_sc_hd__dfxtp_1
X_5527_ _7877_/Q _4226_/A _5527_/S vssd1 vssd1 vccd1 vccd1 _5528_/A sky130_fd_sc_hd__mux2_1
X_8448__223 vssd1 vssd1 vccd1 vccd1 _8448__223/HI partID[9] sky130_fd_sc_hd__conb_1
X_8246_ _8246_/CLK _8246_/D vssd1 vssd1 vccd1 vccd1 _8246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _5473_/S vssd1 vssd1 vccd1 vccd1 _5467_/S sky130_fd_sc_hd__clkbuf_4
X_4409_ _4409_/A vssd1 vssd1 vccd1 vccd1 _8116_/D sky130_fd_sc_hd__clkbuf_1
X_5389_ _7939_/Q _4511_/X _5395_/S vssd1 vssd1 vccd1 vccd1 _5390_/A sky130_fd_sc_hd__mux2_1
X_8177_ _8177_/CLK _8177_/D vssd1 vssd1 vccd1 vccd1 _8177_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3256_ _6657_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3256_/X sky130_fd_sc_hd__clkbuf_16
X_7128_ _8399_/Q _7230_/A _7230_/B vssd1 vssd1 vccd1 vccd1 _7128_/X sky130_fd_sc_hd__and3_1
Xclkbuf_0__3187_ _6409_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3187_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6942__494 _6943__495/A vssd1 vssd1 vccd1 vccd1 _8091_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6652__351 _6656__355/A vssd1 vssd1 vccd1 vccd1 _7932_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7293__119 _7294__120/A vssd1 vssd1 vccd1 vccd1 _8246_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4715_/X _4758_/X _4759_/X vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4691_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4691_/X sky130_fd_sc_hd__clkbuf_4
X_6361_ _6361_/A vssd1 vssd1 vccd1 vccd1 _7736_/D sky130_fd_sc_hd__clkbuf_1
X_5312_ _5327_/S vssd1 vssd1 vccd1 vccd1 _5321_/S sky130_fd_sc_hd__clkbuf_4
X_8100_ _8100_/CLK _8100_/D vssd1 vssd1 vccd1 vccd1 _8100_/Q sky130_fd_sc_hd__dfxtp_1
X_6292_ _7600_/A vssd1 vssd1 vccd1 vccd1 _6292_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8031_ _8031_/CLK _8031_/D vssd1 vssd1 vccd1 vccd1 _8031_/Q sky130_fd_sc_hd__dfxtp_1
X_5243_ _5243_/A _5243_/B _5243_/C vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__or3_1
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5174_ _5243_/A _5174_/B _5174_/C vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__or3_1
XFILLER_96_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _8364_/Q vssd1 vssd1 vccd1 vccd1 _4125_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4056_ _8052_/Q _8047_/Q vssd1 vssd1 vccd1 vccd1 _4056_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_52_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7815_ _7815_/CLK _7815_/D vssd1 vssd1 vccd1 vccd1 _7815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7746_ _7854_/CLK _7746_/D vssd1 vssd1 vccd1 vccd1 _7746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _7995_/Q _7994_/Q _7993_/Q vssd1 vssd1 vccd1 vccd1 _4982_/B sky130_fd_sc_hd__and3_1
X_7677_ _7747_/CLK _7677_/D vssd1 vssd1 vccd1 vccd1 _7677_/Q sky130_fd_sc_hd__dfxtp_1
X_3909_ _3887_/X _8322_/Q _3911_/S vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__mux2_1
X_4889_ _8039_/Q _4407_/X _4891_/S vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__mux2_1
X_7380__14 _7381__15/A vssd1 vssd1 vccd1 vccd1 _8316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3409_ clkbuf_0__3409_/X vssd1 vssd1 vccd1 vccd1 _7055__84/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6559_ _6559_/A vssd1 vssd1 vccd1 vccd1 _7862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8229_ _8235_/CLK _8229_/D vssd1 vssd1 vccd1 vccd1 _8229_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3239_ _6575_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3239_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6489__265 _6489__265/A vssd1 vssd1 vccd1 vccd1 _7822_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6990__532 _6991__533/A vssd1 vssd1 vccd1 vccd1 _8129_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6433__220 _6433__220/A vssd1 vssd1 vccd1 vccd1 _7777_/CLK sky130_fd_sc_hd__inv_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7078__102 _7080__104/A vssd1 vssd1 vccd1 vccd1 _8199_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5930_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5930_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6583__297 _6583__297/A vssd1 vssd1 vccd1 vccd1 _7878_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5861_ _5861_/A vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__clkbuf_1
X_7600_ _7600_/A vssd1 vssd1 vccd1 vccd1 _7600_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6659__357 _6661__359/A vssd1 vssd1 vccd1 vccd1 _7938_/CLK sky130_fd_sc_hd__inv_2
X_5792_ _5792_/A vssd1 vssd1 vccd1 vccd1 _7654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4812_ _4807_/X _4808_/X _4865_/B _4811_/X vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__a211o_1
X_7531_ _7533_/A _7547_/B _7531_/C vssd1 vssd1 vccd1 vccd1 _7532_/A sky130_fd_sc_hd__and3_1
X_4743_ _7783_/Q _4573_/B _4676_/X vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_0__3590_ _7332_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3590_/X sky130_fd_sc_hd__clkbuf_16
X_7462_ _8334_/Q _7458_/X _7461_/X _7426_/B vssd1 vssd1 vccd1 vccd1 _7463_/B sky130_fd_sc_hd__o2bb2a_1
X_4674_ _4674_/A vssd1 vssd1 vccd1 vccd1 _4863_/B sky130_fd_sc_hd__clkbuf_2
X_6344_ _6909_/A _6909_/B _6344_/C _6909_/D vssd1 vssd1 vccd1 vccd1 _6345_/B sky130_fd_sc_hd__or4_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6275_ _6340_/B _6254_/Y _6274_/X _6243_/X vssd1 vssd1 vccd1 vccd1 _6275_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5226_ _5148_/X _5224_/X _5225_/X vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__o21a_1
X_8014_ _8014_/CLK _8014_/D vssd1 vssd1 vccd1 vccd1 _8014_/Q sky130_fd_sc_hd__dfxtp_1
X_6785__390 _6785__390/A vssd1 vssd1 vccd1 vccd1 _7975_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3410_ clkbuf_0__3410_/X vssd1 vssd1 vccd1 vccd1 _7061__89/A sky130_fd_sc_hd__clkbuf_4
X_5157_ _5103_/X _5155_/X _5156_/X vssd1 vssd1 vccd1 vccd1 _5161_/B sky130_fd_sc_hd__o21a_1
X_5088_ _8151_/Q _8135_/Q _8127_/Q _8159_/Q _5043_/A _5037_/X vssd1 vssd1 vccd1 vccd1
+ _5088_/X sky130_fd_sc_hd__mux4_2
X_4108_ _8262_/Q _3943_/X _4112_/S vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4039_ _4039_/A vssd1 vssd1 vccd1 vccd1 _8275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6603__312 _6606__315/A vssd1 vssd1 vccd1 vccd1 _7893_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7729_ _7747_/CLK _7729_/D vssd1 vssd1 vccd1 vccd1 _7729_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7011__550 _7011__550/A vssd1 vssd1 vccd1 vccd1 _8147_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6504__276 _6508__280/A vssd1 vssd1 vccd1 vccd1 _7833_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4390_ _8122_/Q _4386_/X _4402_/S vssd1 vssd1 vccd1 vccd1 _4391_/A sky130_fd_sc_hd__mux2_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _7687_/Q _6048_/X _6051_/X _6059_/X vssd1 vssd1 vccd1 vccd1 _6060_/X sky130_fd_sc_hd__o22a_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5011_ _8312_/Q _8304_/Q _8296_/Q _8320_/Q _5149_/S _5010_/X vssd1 vssd1 vccd1 vccd1
+ _5011_/X sky130_fd_sc_hd__mux4_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6997__538 _6998__539/A vssd1 vssd1 vccd1 vccd1 _8135_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5913_ _5913_/A vssd1 vssd1 vccd1 vccd1 _5913_/X sky130_fd_sc_hd__clkbuf_1
X_5844_ _7629_/A _5844_/B vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__or2_1
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7514_ _8351_/Q _7523_/B _7513_/X vssd1 vssd1 vccd1 vccd1 _7514_/X sky130_fd_sc_hd__or3b_1
X_5775_ _5567_/X _7705_/Q _5777_/S vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4726_ _4726_/A vssd1 vssd1 vccd1 vccd1 _4726_/X sky130_fd_sc_hd__buf_2
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7445_ _7496_/B vssd1 vssd1 vccd1 vccd1 _7513_/A sky130_fd_sc_hd__clkbuf_2
X_4657_ _4594_/X _4656_/X _4819_/A vssd1 vssd1 vccd1 vccd1 _4657_/X sky130_fd_sc_hd__a21o_1
X_7376_ _7382_/A vssd1 vssd1 vccd1 vccd1 _7376_/X sky130_fd_sc_hd__buf_1
Xinput91 wbs_we_i vssd1 vssd1 vccd1 vccd1 _6185_/C sky130_fd_sc_hd__buf_8
Xinput80 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _7629_/A sky130_fd_sc_hd__buf_6
X_6327_ _7725_/Q _6320_/X _6324_/X _6326_/X vssd1 vssd1 vccd1 vccd1 _7725_/D sky130_fd_sc_hd__a211o_1
X_4588_ _4714_/A vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6258_ _7713_/Q _6216_/X _6257_/X vssd1 vssd1 vccd1 vccd1 _7713_/D sky130_fd_sc_hd__a21o_1
X_6189_ _6188_/X _6189_/B vssd1 vssd1 vccd1 vccd1 _6190_/A sky130_fd_sc_hd__and2b_1
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5209_ _5191_/A _5207_/X _5208_/X vssd1 vssd1 vccd1 vccd1 _5210_/C sky130_fd_sc_hd__o21a_1
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3255_ clkbuf_0__3255_/X vssd1 vssd1 vccd1 vccd1 _6656__355/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3890_ _8358_/Q vssd1 vssd1 vccd1 vccd1 _3890_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0__3390_ clkbuf_0__3390_/X vssd1 vssd1 vccd1 vccd1 _6961__509/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5560_/A vssd1 vssd1 vccd1 vccd1 _7841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4511_ _8364_/Q vssd1 vssd1 vccd1 vccd1 _4511_/X sky130_fd_sc_hd__clkbuf_2
X_5491_ _7893_/Q _4226_/A _5491_/S vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__mux2_1
X_7230_ _7230_/A _7230_/B vssd1 vssd1 vccd1 vccd1 _7230_/Y sky130_fd_sc_hd__nand2_1
X_4442_ _4214_/X _8103_/Q _4444_/S vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7161_ _7430_/A _7226_/A _7226_/B vssd1 vssd1 vccd1 vccd1 _7161_/X sky130_fd_sc_hd__and3_1
X_4373_ _4373_/A vssd1 vssd1 vccd1 vccd1 _8129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7092_ _7092_/A _7098_/A _7098_/B _7134_/A vssd1 vssd1 vccd1 vccd1 _7221_/A sky130_fd_sc_hd__or4_1
X_6112_ _6104_/X _7693_/Q _6107_/X _6111_/X _7661_/Q vssd1 vssd1 vccd1 vccd1 _7661_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6043_ _7680_/Q _6032_/X _6039_/X _6042_/X vssd1 vssd1 vccd1 vccd1 _6043_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6446__230 _6446__230/A vssd1 vssd1 vccd1 vccd1 _7787_/CLK sky130_fd_sc_hd__inv_2
X_7994_ _7994_/CLK _7994_/D vssd1 vssd1 vccd1 vccd1 _7994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_5827_ _5827_/A vssd1 vssd1 vccd1 vccd1 _5827_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3588_ clkbuf_0__3588_/X vssd1 vssd1 vccd1 vccd1 _7325__145/A sky130_fd_sc_hd__clkbuf_4
X_5758_ _5758_/A vssd1 vssd1 vccd1 vccd1 _7758_/D sky130_fd_sc_hd__clkbuf_1
X_4709_ _8025_/Q _7980_/Q _7840_/Q _8208_/Q _4596_/X _4580_/X vssd1 vssd1 vccd1 vccd1
+ _4709_/X sky130_fd_sc_hd__mux4_1
X_7428_ _7615_/A _6714_/B _7425_/X _7426_/X _7427_/X vssd1 vssd1 vccd1 vccd1 _7435_/B
+ sky130_fd_sc_hd__o2111a_1
X_5689_ _5743_/A _5689_/B vssd1 vssd1 vccd1 vccd1 _5705_/S sky130_fd_sc_hd__nor2_2
XFILLER_116_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6730_ _8406_/Q _8331_/Q vssd1 vssd1 vccd1 vccd1 _7425_/A sky130_fd_sc_hd__xor2_1
X_4991_ _5100_/B vssd1 vssd1 vccd1 vccd1 _5237_/S sky130_fd_sc_hd__buf_2
X_3942_ _8363_/Q vssd1 vssd1 vccd1 vccd1 _4211_/A sky130_fd_sc_hd__clkbuf_4
X_3873_ _3872_/X _8372_/Q _3882_/S vssd1 vssd1 vccd1 vccd1 _3874_/A sky130_fd_sc_hd__mux2_1
X_8400_ _8407_/CLK _8400_/D vssd1 vssd1 vccd1 vccd1 _8400_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3373_ clkbuf_0__3373_/X vssd1 vssd1 vccd1 vccd1 _6913_/A sky130_fd_sc_hd__clkbuf_4
X_5612_ _5612_/A vssd1 vssd1 vccd1 vccd1 _7823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8331_ _8399_/CLK _8331_/D vssd1 vssd1 vccd1 vccd1 _8331_/Q sky130_fd_sc_hd__dfxtp_1
X_5543_ _5304_/X _7870_/Q _5545_/S vssd1 vssd1 vccd1 vccd1 _5544_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3410_ _7057_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3410_/X sky130_fd_sc_hd__clkbuf_16
X_8262_ _8262_/CLK _8262_/D vssd1 vssd1 vccd1 vccd1 _8262_/Q sky130_fd_sc_hd__dfxtp_1
X_5474_ _5474_/A vssd1 vssd1 vccd1 vccd1 _7901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4425_ _4425_/A vssd1 vssd1 vccd1 vccd1 _8111_/D sky130_fd_sc_hd__clkbuf_1
X_7213_ _7218_/A _7213_/B vssd1 vssd1 vccd1 vccd1 _8216_/D sky130_fd_sc_hd__nor2_1
X_8193_ _8193_/CLK _8193_/D vssd1 vssd1 vccd1 vccd1 _8193_/Q sky130_fd_sc_hd__dfxtp_1
X_7144_ _7138_/X _7139_/Y _7141_/Y _7142_/Y _7143_/X vssd1 vssd1 vccd1 vccd1 _7144_/X
+ sky130_fd_sc_hd__o2111a_1
X_4356_ _8136_/Q _4128_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4287_ _5348_/A _4368_/B vssd1 vssd1 vccd1 vccd1 _4303_/S sky130_fd_sc_hd__or2_4
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7075_/A vssd1 vssd1 vccd1 vccd1 _7075_/X sky130_fd_sc_hd__buf_1
XFILLER_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6026_ _7546_/A vssd1 vssd1 vccd1 vccd1 _7608_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7977_ _7977_/CLK _7977_/D vssd1 vssd1 vccd1 vccd1 _7977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6859_ _6871_/A vssd1 vssd1 vccd1 vccd1 _6859_/X sky130_fd_sc_hd__buf_1
XFILLER_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6954__503 _6955__504/A vssd1 vssd1 vccd1 vccd1 _8100_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4210_ _4210_/A vssd1 vssd1 vccd1 vccd1 _8193_/D sky130_fd_sc_hd__clkbuf_1
X_5190_ _8290_/Q _8298_/Q _5207_/S vssd1 vssd1 vccd1 vccd1 _5191_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4141_ _8250_/Q _4140_/X _4144_/S vssd1 vssd1 vccd1 vccd1 _4142_/A sky130_fd_sc_hd__mux2_1
X_4072_ _4057_/X _4060_/X _4068_/X _4071_/Y vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__a211o_2
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7900_ _7900_/CLK _7900_/D vssd1 vssd1 vccd1 vccd1 _7900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7831_ _7831_/CLK _7831_/D vssd1 vssd1 vccd1 vccd1 _7831_/Q sky130_fd_sc_hd__dfxtp_1
X_7762_ _7762_/CLK _7762_/D vssd1 vssd1 vccd1 vccd1 _7762_/Q sky130_fd_sc_hd__dfxtp_1
X_4974_ _5008_/A vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__clkbuf_2
X_6713_ _6713_/A vssd1 vssd1 vccd1 vccd1 _6714_/B sky130_fd_sc_hd__clkbuf_2
X_7693_ _8365_/CLK _7693_/D vssd1 vssd1 vccd1 vccd1 _7693_/Q sky130_fd_sc_hd__dfxtp_1
X_3925_ _3925_/A vssd1 vssd1 vccd1 vccd1 _8317_/D sky130_fd_sc_hd__clkbuf_1
X_6644_ _6644_/A vssd1 vssd1 vccd1 vccd1 _6644_/X sky130_fd_sc_hd__buf_1
X_3856_ _8377_/Q _3831_/X _3856_/S vssd1 vssd1 vccd1 vccd1 _3857_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3787_ _7999_/Q _7998_/Q vssd1 vssd1 vccd1 vccd1 _3893_/A sky130_fd_sc_hd__nand2_1
X_6575_ _6575_/A vssd1 vssd1 vccd1 vccd1 _6575_/X sky130_fd_sc_hd__buf_1
XFILLER_118_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8314_ _8314_/CLK _8314_/D vssd1 vssd1 vccd1 vccd1 _8314_/Q sky130_fd_sc_hd__dfxtp_1
X_5526_ _5526_/A vssd1 vssd1 vccd1 vccd1 _7878_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8245_ _8245_/CLK _8245_/D vssd1 vssd1 vccd1 vccd1 _8245_/Q sky130_fd_sc_hd__dfxtp_1
X_5457_ _5475_/A _5457_/B vssd1 vssd1 vccd1 vccd1 _5473_/S sky130_fd_sc_hd__nor2_2
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4408_ _8116_/Q _4407_/X _4411_/S vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__mux2_1
X_5388_ _5388_/A vssd1 vssd1 vccd1 vccd1 _7940_/D sky130_fd_sc_hd__clkbuf_1
X_8176_ _8176_/CLK _8176_/D vssd1 vssd1 vccd1 vccd1 _8176_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3255_ _6651_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3255_/X sky130_fd_sc_hd__clkbuf_16
X_7127_ _7230_/A _7230_/B _7615_/A vssd1 vssd1 vccd1 vccd1 _7127_/Y sky130_fd_sc_hd__a21oi_1
X_4339_ _4338_/X _8142_/Q _4339_/S vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__mux2_1
X_6009_ _6400_/A vssd1 vssd1 vccd1 vccd1 _6023_/S sky130_fd_sc_hd__buf_2
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7327__146 _7329__148/A vssd1 vssd1 vccd1 vccd1 _8273_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7056__85 _7056__85/A vssd1 vssd1 vccd1 vccd1 _8182_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _4696_/A vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__buf_2
X_6360_ _5918_/A _7736_/Q _6360_/S vssd1 vssd1 vccd1 vccd1 _6361_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5311_ _5795_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _5327_/S sky130_fd_sc_hd__or2_2
XFILLER_114_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6291_ _7718_/Q _6320_/A vssd1 vssd1 vccd1 vccd1 _6291_/X sky130_fd_sc_hd__and2_1
X_8030_ _8030_/CLK _8030_/D vssd1 vssd1 vccd1 vccd1 _8030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5242_ _5148_/A _5240_/X _5241_/X vssd1 vssd1 vccd1 vccd1 _5243_/C sky130_fd_sc_hd__o21a_1
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8408__230 vssd1 vssd1 vccd1 vccd1 core1Index[0] _8408__230/LO sky130_fd_sc_hd__conb_1
X_5173_ _5130_/A _5171_/X _5172_/X vssd1 vssd1 vccd1 vccd1 _5174_/C sky130_fd_sc_hd__o21a_1
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4124_ _4124_/A vssd1 vssd1 vccd1 vccd1 _8256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
X_4055_ _4059_/B vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7814_ _7814_/CLK _7814_/D vssd1 vssd1 vccd1 vccd1 _7814_/Q sky130_fd_sc_hd__dfxtp_1
X_7745_ _7854_/CLK _7745_/D vssd1 vssd1 vccd1 vccd1 _7745_/Q sky130_fd_sc_hd__dfxtp_1
X_4957_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7676_ _7854_/CLK _7676_/D vssd1 vssd1 vccd1 vccd1 _7676_/Q sky130_fd_sc_hd__dfxtp_1
X_4888_ _4888_/A vssd1 vssd1 vccd1 vccd1 _8040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3908_ _3908_/A vssd1 vssd1 vccd1 vccd1 _8323_/D sky130_fd_sc_hd__clkbuf_1
X_3839_ _3839_/A vssd1 vssd1 vccd1 vccd1 _8383_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3408_ clkbuf_0__3408_/X vssd1 vssd1 vccd1 vccd1 _7048__78/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6558_ _7862_/Q _5891_/A _6564_/S vssd1 vssd1 vccd1 vccd1 _6559_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5509_ _5308_/X _7885_/Q _5509_/S vssd1 vssd1 vccd1 vccd1 _5510_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8228_ _8364_/CLK _8228_/D vssd1 vssd1 vccd1 vccd1 _8228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8159_ _8159_/CLK _8159_/D vssd1 vssd1 vccd1 vccd1 _8159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7029__63 _7029__63/A vssd1 vssd1 vccd1 vccd1 _8160_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _7605_/B _5866_/B vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__or2_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4869_/B _4809_/X _4810_/X vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5791_ _7654_/Q _5567_/A _5793_/S vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7530_ _8357_/Q _7529_/B _7529_/Y _7493_/A vssd1 vssd1 vccd1 vccd1 _8357_/D sky130_fd_sc_hd__o211a_1
X_4742_ _4338_/X _4538_/X _4741_/X _4609_/X vssd1 vssd1 vccd1 vccd1 _8060_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7461_ _7474_/A vssd1 vssd1 vccd1 vccd1 _7461_/X sky130_fd_sc_hd__clkbuf_2
X_4673_ _4335_/X _4538_/X _4672_/X _4609_/X vssd1 vssd1 vccd1 vccd1 _8061_/D sky130_fd_sc_hd__o211a_1
X_6343_ _7734_/Q _6343_/B vssd1 vssd1 vccd1 vccd1 _6909_/D sky130_fd_sc_hd__nand2_1
XFILLER_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6274_ _8061_/Q _6231_/A _6201_/X _6235_/X vssd1 vssd1 vccd1 vccd1 _6274_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8013_ _8364_/CLK _8013_/D vssd1 vssd1 vccd1 vccd1 _8013_/Q sky130_fd_sc_hd__dfxtp_1
X_5225_ _8091_/Q _5150_/X _5125_/A _8249_/Q _5003_/A vssd1 vssd1 vccd1 vccd1 _5225_/X
+ sky130_fd_sc_hd__o221a_1
X_5156_ _8093_/Q _5150_/X _5125_/A _8251_/Q _5003_/A vssd1 vssd1 vccd1 vccd1 _5156_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4107_ _4107_/A vssd1 vssd1 vccd1 vccd1 _8263_/D sky130_fd_sc_hd__clkbuf_1
X_5087_ _8253_/Q _8167_/Q _7905_/Q _8095_/Q _5037_/A _5220_/S vssd1 vssd1 vccd1 vccd1
+ _5087_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4038_ _8275_/Q _3955_/X _4042_/S vssd1 vssd1 vccd1 vccd1 _4039_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5989_ _7666_/Q _5988_/X _5989_/S vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__mux2_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7728_ _7747_/CLK _7728_/D vssd1 vssd1 vccd1 vccd1 _7728_/Q sky130_fd_sc_hd__dfxtp_1
X_7659_ _7659_/CLK _7659_/D vssd1 vssd1 vccd1 vccd1 _7659_/Q sky130_fd_sc_hd__dfxtp_1
X_6495__270 _6495__270/A vssd1 vssd1 vccd1 vccd1 _7827_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput190 _5998_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__buf_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5912_ _5912_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__and2_1
X_5843_ _5843_/A vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7513_ _7513_/A vssd1 vssd1 vccd1 vccd1 _7513_/X sky130_fd_sc_hd__clkbuf_1
X_5774_ _5774_/A vssd1 vssd1 vccd1 vccd1 _7706_/D sky130_fd_sc_hd__clkbuf_1
X_4725_ _4725_/A vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__clkbuf_2
X_7444_ _7529_/A _7447_/B _7442_/Y _7450_/A _7493_/A vssd1 vssd1 vccd1 vccd1 _8330_/D
+ sky130_fd_sc_hd__o221a_1
X_4656_ _8087_/Q _8079_/Q _8042_/Q _8111_/Q _4582_/X _4571_/X vssd1 vssd1 vccd1 vccd1
+ _4656_/X sky130_fd_sc_hd__mux4_1
X_4587_ _4567_/X _4581_/X _4586_/X vssd1 vssd1 vccd1 vccd1 _4587_/X sky130_fd_sc_hd__a21o_1
Xinput81 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _7626_/A sky130_fd_sc_hd__buf_6
Xinput70 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__buf_4
X_6326_ _7599_/A _6326_/B _6332_/C _6326_/D vssd1 vssd1 vccd1 vccd1 _6326_/X sky130_fd_sc_hd__and4_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _6221_/X _6252_/X _6256_/X _6246_/X vssd1 vssd1 vccd1 vccd1 _6257_/X sky130_fd_sc_hd__a31o_1
X_6188_ _6188_/A _6188_/B _6188_/C vssd1 vssd1 vccd1 vccd1 _6188_/X sky130_fd_sc_hd__and3_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _5114_/X _7910_/Q _5125_/X _8180_/Q _5123_/S vssd1 vssd1 vccd1 vccd1 _5208_/X
+ sky130_fd_sc_hd__o221a_1
X_5139_ _5130_/A _5137_/X _5138_/X vssd1 vssd1 vccd1 vccd1 _5140_/C sky130_fd_sc_hd__o21a_1
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i _7717_/CLK vssd1 vssd1 vccd1 vccd1 _7854_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7559__34 _7559__34/A vssd1 vssd1 vccd1 vccd1 _8373_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3254_ clkbuf_0__3254_/X vssd1 vssd1 vccd1 vccd1 _6681_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7023__58 _7025__60/A vssd1 vssd1 vccd1 vccd1 _8155_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6510__281 _6511__282/A vssd1 vssd1 vccd1 vccd1 _7838_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5490_ _5490_/A vssd1 vssd1 vccd1 vccd1 _7894_/D sky130_fd_sc_hd__clkbuf_1
X_4510_ _4510_/A vssd1 vssd1 vccd1 vccd1 _8074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4441_ _4441_/A vssd1 vssd1 vccd1 vccd1 _8104_/D sky130_fd_sc_hd__clkbuf_1
X_7160_ _8219_/Q _7110_/C _7129_/A _7119_/A _8220_/Q vssd1 vssd1 vccd1 vccd1 _7226_/B
+ sky130_fd_sc_hd__a41o_1
X_6111_ _6129_/A vssd1 vssd1 vccd1 vccd1 _6111_/X sky130_fd_sc_hd__buf_4
X_4372_ _4208_/X _8129_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _8216_/Q _7208_/A _8214_/Q _7140_/B vssd1 vssd1 vccd1 vccd1 _7134_/A sky130_fd_sc_hd__nand4_4
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6042_ _6042_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6042_/X sky130_fd_sc_hd__and2_1
XFILLER_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7993_ _7993_/CLK _7993_/D vssd1 vssd1 vccd1 vccd1 _7993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6944_ _6944_/A vssd1 vssd1 vccd1 vccd1 _6944_/X sky130_fd_sc_hd__buf_1
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5826_ _6518_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5827_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3587_ clkbuf_0__3587_/X vssd1 vssd1 vccd1 vccd1 _7316__137/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5757_ _7758_/Q _5567_/A _5759_/S vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__mux2_1
X_4708_ _4677_/X _4693_/X _4865_/B _4707_/X vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__a211o_1
XFILLER_108_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7427_ _7429_/A _7429_/B _7096_/A vssd1 vssd1 vccd1 vccd1 _7427_/X sky130_fd_sc_hd__a21o_1
X_5688_ _5688_/A vssd1 vssd1 vccd1 vccd1 _7789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4639_ _4594_/X _4638_/X _4575_/X vssd1 vssd1 vccd1 vccd1 _4639_/X sky130_fd_sc_hd__a21o_1
X_6309_ _6309_/A vssd1 vssd1 vccd1 vccd1 _6337_/B sky130_fd_sc_hd__clkbuf_1
X_6826__409 _6826__409/A vssd1 vssd1 vccd1 vccd1 _8002_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7289_ _7295_/A vssd1 vssd1 vccd1 vccd1 _7289_/X sky130_fd_sc_hd__buf_1
XFILLER_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6616__323 _6618__325/A vssd1 vssd1 vccd1 vccd1 _7904_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4990_ _5003_/A vssd1 vssd1 vccd1 vccd1 _4990_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3941_ _3941_/A vssd1 vssd1 vccd1 vccd1 _8311_/D sky130_fd_sc_hd__clkbuf_1
X_3872_ _8364_/Q vssd1 vssd1 vccd1 vccd1 _3872_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3372_ clkbuf_0__3372_/X vssd1 vssd1 vccd1 vccd1 _6882__450/A sky130_fd_sc_hd__clkbuf_4
X_7553__29 _7553__29/A vssd1 vssd1 vccd1 vccd1 _8368_/CLK sky130_fd_sc_hd__inv_2
X_5611_ _5564_/X _7823_/Q _5615_/S vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__mux2_1
X_8330_ _8332_/CLK _8330_/D vssd1 vssd1 vccd1 vccd1 _8330_/Q sky130_fd_sc_hd__dfxtp_1
X_5542_ _5542_/A vssd1 vssd1 vccd1 vccd1 _7871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8261_ _8261_/CLK _8261_/D vssd1 vssd1 vccd1 vccd1 _8261_/Q sky130_fd_sc_hd__dfxtp_1
X_5473_ _7901_/Q _4226_/A _5473_/S vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6517__287 _6517__287/A vssd1 vssd1 vccd1 vccd1 _7844_/CLK sky130_fd_sc_hd__inv_2
X_4424_ _8111_/Q _4398_/X _4426_/S vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__mux2_1
X_7212_ _6198_/X _7135_/B _7198_/X _7194_/X _7211_/Y vssd1 vssd1 vccd1 vccd1 _7213_/B
+ sky130_fd_sc_hd__o32a_1
X_8192_ _8192_/CLK _8192_/D vssd1 vssd1 vccd1 vccd1 _8192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7143_ _7143_/A _7199_/A vssd1 vssd1 vccd1 vccd1 _7143_/X sky130_fd_sc_hd__or2_1
X_4355_ _4355_/A vssd1 vssd1 vccd1 vccd1 _8137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4286_ _4286_/A _4286_/B _4120_/C vssd1 vssd1 vccd1 vccd1 _4368_/B sky130_fd_sc_hd__or3b_4
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _7728_/Q input10/X _6025_/S vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7976_ _7976_/CLK _7976_/D vssd1 vssd1 vccd1 vccd1 _7976_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5809_ _4096_/X _7646_/Q _5811_/S vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6912__470 _6912__470/A vssd1 vssd1 vccd1 vccd1 _8067_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_50 _5914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8432__207 vssd1 vssd1 vccd1 vccd1 _8432__207/HI core1Index[7] sky130_fd_sc_hd__conb_1
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4140_ _8359_/Q vssd1 vssd1 vccd1 vccd1 _4140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4071_ _4536_/D _4070_/X _4853_/A vssd1 vssd1 vccd1 vccd1 _4071_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7830_ _7830_/CLK _7830_/D vssd1 vssd1 vccd1 vccd1 _7830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7761_ _7761_/CLK _7761_/D vssd1 vssd1 vccd1 vccd1 _7761_/Q sky130_fd_sc_hd__dfxtp_1
X_4973_ _4982_/B _5126_/A vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7692_ _8342_/CLK _7692_/D vssd1 vssd1 vccd1 vccd1 _7692_/Q sky130_fd_sc_hd__dfxtp_1
X_6712_ _6702_/B _6702_/C _6716_/A _6711_/Y vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__a22o_1
X_3924_ _3878_/X _8317_/Q _3926_/S vssd1 vssd1 vccd1 vccd1 _3925_/A sky130_fd_sc_hd__mux2_1
X_7392__24 _7393__25/A vssd1 vssd1 vccd1 vccd1 _8326_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3855_ _3855_/A vssd1 vssd1 vccd1 vccd1 _8378_/D sky130_fd_sc_hd__clkbuf_1
X_3786_ _8001_/Q _3783_/Y _4950_/B _5249_/B vssd1 vssd1 vccd1 vccd1 _3793_/B sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8341_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_8313_ _8313_/CLK _8313_/D vssd1 vssd1 vccd1 vccd1 _8313_/Q sky130_fd_sc_hd__dfxtp_1
X_5525_ _7878_/Q _4223_/A _5527_/S vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5456_ _5456_/A vssd1 vssd1 vccd1 vccd1 _7909_/D sky130_fd_sc_hd__clkbuf_1
X_8244_ _8244_/CLK _8244_/D vssd1 vssd1 vccd1 vccd1 _8244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3254_ _6650_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3254_/X sky130_fd_sc_hd__clkbuf_16
X_4407_ _7986_/Q vssd1 vssd1 vccd1 vccd1 _4407_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5387_ _7940_/Q _5366_/X _5395_/S vssd1 vssd1 vccd1 vccd1 _5388_/A sky130_fd_sc_hd__mux2_1
X_8175_ _8175_/CLK _8175_/D vssd1 vssd1 vccd1 vccd1 _8175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7126_ _7119_/A _7159_/B _8221_/Q vssd1 vssd1 vccd1 vccd1 _7230_/B sky130_fd_sc_hd__a21o_1
X_4338_ _7988_/Q vssd1 vssd1 vccd1 vccd1 _4338_/X sky130_fd_sc_hd__buf_2
XFILLER_101_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7057_/X sky130_fd_sc_hd__buf_1
X_4269_ _4284_/S vssd1 vssd1 vccd1 vccd1 _4278_/S sky130_fd_sc_hd__clkbuf_2
X_6008_ _7723_/Q input5/X _6008_/S vssd1 vssd1 vccd1 vccd1 _6008_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7959_/CLK _7959_/D vssd1 vssd1 vccd1 vccd1 _7959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6878__446 _6879__447/A vssd1 vssd1 vccd1 vccd1 _8041_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6290_ _6719_/A _6839_/C _6337_/D _6288_/X _6289_/X vssd1 vssd1 vccd1 vccd1 _6290_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5310_ _5310_/A vssd1 vssd1 vccd1 vccd1 _7977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5241_ _5113_/A _7909_/Q _5151_/A _8179_/Q _5008_/A vssd1 vssd1 vccd1 vccd1 _5241_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6668__360 _6668__360/A vssd1 vssd1 vccd1 vccd1 _7944_/CLK sky130_fd_sc_hd__inv_2
X_5172_ _5113_/A _7911_/Q _5151_/A _8181_/Q _4987_/A vssd1 vssd1 vccd1 vccd1 _5172_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6629__333 _6631__335/A vssd1 vssd1 vccd1 vccd1 _7914_/CLK sky130_fd_sc_hd__inv_2
X_4123_ _8256_/Q _3966_/X _4135_/S vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__mux2_1
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4054_ _8046_/Q vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__inv_2
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7813_ _7813_/CLK _7813_/D vssd1 vssd1 vccd1 vccd1 _7813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7744_ _7854_/CLK _7744_/D vssd1 vssd1 vccd1 vccd1 _7744_/Q sky130_fd_sc_hd__dfxtp_1
X_4956_ _4956_/A _7265_/A vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__nor2_1
X_7675_ _7854_/CLK _7675_/D vssd1 vssd1 vccd1 vccd1 _7675_/Q sky130_fd_sc_hd__dfxtp_1
X_4887_ _8040_/Q _4404_/X _4891_/S vssd1 vssd1 vccd1 vccd1 _4888_/A sky130_fd_sc_hd__mux2_1
X_3907_ _3884_/X _8323_/Q _3911_/S vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__mux2_1
X_3838_ _8383_/Q _3837_/X _3841_/S vssd1 vssd1 vccd1 vccd1 _3839_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3407_ clkbuf_0__3407_/X vssd1 vssd1 vccd1 vccd1 _7063_/A sky130_fd_sc_hd__clkbuf_4
X_6626_ _6632_/A vssd1 vssd1 vccd1 vccd1 _6626_/X sky130_fd_sc_hd__buf_1
X_6557_ _6557_/A vssd1 vssd1 vccd1 vccd1 _7861_/D sky130_fd_sc_hd__clkbuf_1
X_5508_ _5508_/A vssd1 vssd1 vccd1 vccd1 _7886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8227_ _8364_/CLK _8227_/D vssd1 vssd1 vccd1 vccd1 _8227_/Q sky130_fd_sc_hd__dfxtp_1
X_5439_ _5439_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5455_/S sky130_fd_sc_hd__or2_2
X_8158_ _8158_/CLK _8158_/D vssd1 vssd1 vccd1 vccd1 _8158_/Q sky130_fd_sc_hd__dfxtp_1
X_7109_ _8223_/Q vssd1 vssd1 vccd1 vccd1 _7237_/A sky130_fd_sc_hd__inv_2
X_8089_ _8089_/CLK _8089_/D vssd1 vssd1 vccd1 vccd1 _8089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925__480 _6925__480/A vssd1 vssd1 vccd1 vccd1 _8077_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8438__213 vssd1 vssd1 vccd1 vccd1 _8438__213/HI manufacturerID[5] sky130_fd_sc_hd__conb_1
X_4810_ _4703_/X _7805_/Q _7645_/Q _4725_/X _4726_/X vssd1 vssd1 vccd1 vccd1 _4810_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5790_ _5790_/A vssd1 vssd1 vccd1 vccd1 _7655_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4540_/X _8060_/Q _4632_/X _4740_/X _4605_/X vssd1 vssd1 vccd1 vccd1 _4741_/X
+ sky130_fd_sc_hd__a221o_1
X_7460_ _7470_/A _7460_/B vssd1 vssd1 vccd1 vccd1 _8333_/D sky130_fd_sc_hd__nor2_1
X_4672_ _4540_/X _8061_/Q _4632_/X _4671_/X _4605_/X vssd1 vssd1 vccd1 vccd1 _4672_/X
+ sky130_fd_sc_hd__a221o_1
X_6967__514 _6968__515/A vssd1 vssd1 vccd1 vccd1 _8111_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6342_ _6342_/A _6342_/B _7732_/Q vssd1 vssd1 vccd1 vccd1 _6344_/C sky130_fd_sc_hd__or3b_1
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6273_ _8403_/Q _6249_/X _6251_/X _6228_/X vssd1 vssd1 vccd1 vccd1 _6273_/X sky130_fd_sc_hd__a31o_1
X_8012_ _8065_/CLK _8012_/D vssd1 vssd1 vccd1 vccd1 _8012_/Q sky130_fd_sc_hd__dfxtp_1
X_5224_ _8163_/Q _7901_/Q _5224_/S vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5155_ _8165_/Q _7903_/Q _5224_/S vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4106_ _8263_/Q _3939_/X _4112_/S vssd1 vssd1 vccd1 vccd1 _4107_/A sky130_fd_sc_hd__mux2_1
X_5086_ _5009_/X _5085_/X _5119_/A vssd1 vssd1 vccd1 vccd1 _5086_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _4037_/A vssd1 vssd1 vccd1 vccd1 _8276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _7717_/Q input30/X _5991_/S vssd1 vssd1 vccd1 vccd1 _5988_/X sky130_fd_sc_hd__mux2_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7727_ _7747_/CLK _7727_/D vssd1 vssd1 vccd1 vccd1 _7727_/Q sky130_fd_sc_hd__dfxtp_1
X_4939_ _4335_/X _8018_/Q _4941_/S vssd1 vssd1 vccd1 vccd1 _4940_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7658_ _7658_/CLK _7658_/D vssd1 vssd1 vccd1 vccd1 _7658_/Q sky130_fd_sc_hd__dfxtp_1
X_6417__206 _6418__207/A vssd1 vssd1 vccd1 vccd1 _7763_/CLK sky130_fd_sc_hd__inv_2
X_7589_ _7602_/A vssd1 vssd1 vccd1 vccd1 _7615_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_opt_1_0_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
X_6610__318 _6611__319/A vssd1 vssd1 vccd1 vccd1 _7899_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput191 _6001_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__buf_2
Xoutput180 _6063_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__buf_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3399_ clkbuf_0__3399_/X vssd1 vssd1 vccd1 vccd1 _7011__550/A sky130_fd_sc_hd__clkbuf_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6769__376 _6772__379/A vssd1 vssd1 vccd1 vccd1 _7961_/CLK sky130_fd_sc_hd__inv_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5920_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5842_ _7538_/B _5844_/B vssd1 vssd1 vccd1 vccd1 _5843_/A sky130_fd_sc_hd__or2_1
XFILLER_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5773_ _5564_/X _7706_/Q _5777_/S vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__mux2_1
X_7512_ _7527_/B vssd1 vssd1 vccd1 vccd1 _7523_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4724_ _4724_/A vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__clkbuf_2
X_7443_ _7519_/A vssd1 vssd1 vccd1 vccd1 _7493_/A sky130_fd_sc_hd__clkbuf_2
X_4655_ _8245_/Q _8143_/Q _7825_/Q _8269_/Q _4579_/X _4562_/X vssd1 vssd1 vccd1 vccd1
+ _4655_/X sky130_fd_sc_hd__mux4_1
X_4586_ _4557_/A _4583_/X _4819_/A vssd1 vssd1 vccd1 vccd1 _4586_/X sky130_fd_sc_hd__a21o_1
Xinput82 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _7546_/B sky130_fd_sc_hd__buf_6
Xinput60 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _7591_/B sky130_fd_sc_hd__buf_4
Xinput71 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__buf_4
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6325_ _8394_/Q vssd1 vssd1 vccd1 vccd1 _7599_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3037_ clkbuf_0__3037_/X vssd1 vssd1 vccd1 vccd1 _6213__199/A sky130_fd_sc_hd__clkbuf_4
X_6256_ _6253_/Y _6254_/Y _6255_/X _6243_/X vssd1 vssd1 vccd1 vccd1 _6256_/X sky130_fd_sc_hd__a22o_1
X_6187_ _6187_/A vssd1 vssd1 vccd1 vccd1 _7701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5207_ _8172_/Q _7894_/Q _5207_/S vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5138_ _5113_/A _7912_/Q _5151_/A _8182_/Q _4987_/A vssd1 vssd1 vccd1 vccd1 _5138_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5069_ _8152_/Q _8136_/Q _8128_/Q _8160_/Q _5043_/A _5037_/X vssd1 vssd1 vccd1 vccd1
+ _5069_/X sky130_fd_sc_hd__mux4_2
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3253_ clkbuf_0__3253_/X vssd1 vssd1 vccd1 vccd1 _6649__350/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6085__176 _6087__178/A vssd1 vssd1 vccd1 vccd1 _7645_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4211_/X _8104_/Q _4444_/S vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__mux2_1
X_7346__161 _7350__165/A vssd1 vssd1 vccd1 vccd1 _8288_/CLK sky130_fd_sc_hd__inv_2
X_6110_ _6154_/A vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__buf_4
X_4371_ _4371_/A vssd1 vssd1 vccd1 vccd1 _8130_/D sky130_fd_sc_hd__clkbuf_1
X_7090_ _8213_/Q vssd1 vssd1 vccd1 vccd1 _7140_/B sky130_fd_sc_hd__clkbuf_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6052_/A vssd1 vssd1 vccd1 vccd1 _6049_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7992_ _7992_/CLK _7992_/D vssd1 vssd1 vccd1 vccd1 _7992_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3724_ clkbuf_0__3724_/X vssd1 vssd1 vccd1 vccd1 _7574__46/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5825_ _5825_/A vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3586_ clkbuf_0__3586_/X vssd1 vssd1 vccd1 vccd1 _7311__133/A sky130_fd_sc_hd__clkbuf_4
X_5756_ _5756_/A vssd1 vssd1 vccd1 vccd1 _7759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4707_ _4869_/B _4700_/X _4706_/X vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__o21a_1
X_5687_ _7789_/Q _5596_/X _5687_/S vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__mux2_1
X_7426_ _8403_/Q _7426_/B vssd1 vssd1 vccd1 vccd1 _7426_/X sky130_fd_sc_hd__xor2_1
X_4638_ _8019_/Q _7874_/Q _7778_/Q _7762_/Q _4582_/X _4580_/A vssd1 vssd1 vccd1 vccd1
+ _4638_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4569_ _4596_/A vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__buf_2
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7357_ _7357_/A vssd1 vssd1 vccd1 vccd1 _7357_/X sky130_fd_sc_hd__buf_1
XFILLER_89_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6308_ _8398_/Q vssd1 vssd1 vccd1 vccd1 _7612_/A sky130_fd_sc_hd__buf_4
X_6239_ _6350_/C _6285_/A _6226_/B _6909_/C _6238_/Y vssd1 vssd1 vccd1 vccd1 _6254_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6623__328 _6625__330/A vssd1 vssd1 vccd1 vccd1 _7909_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3940_ _8311_/Q _3939_/X _3952_/S vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3871_ _3871_/A vssd1 vssd1 vccd1 vccd1 _8373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3371_ clkbuf_0__3371_/X vssd1 vssd1 vccd1 vccd1 _6873__442/A sky130_fd_sc_hd__clkbuf_4
X_5610_ _5610_/A vssd1 vssd1 vccd1 vccd1 _7824_/D sky130_fd_sc_hd__clkbuf_1
X_5541_ _5300_/X _7871_/Q _5545_/S vssd1 vssd1 vccd1 vccd1 _5542_/A sky130_fd_sc_hd__mux2_1
X_8260_ _8260_/CLK _8260_/D vssd1 vssd1 vccd1 vccd1 _8260_/Q sky130_fd_sc_hd__dfxtp_1
X_7211_ _8216_/Q vssd1 vssd1 vccd1 vccd1 _7211_/Y sky130_fd_sc_hd__inv_2
X_5472_ _5472_/A vssd1 vssd1 vccd1 vccd1 _7902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4423_ _4423_/A vssd1 vssd1 vccd1 vccd1 _8112_/D sky130_fd_sc_hd__clkbuf_1
X_8191_ _8191_/CLK _8191_/D vssd1 vssd1 vccd1 vccd1 _8191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7142_ _7143_/A _7199_/A vssd1 vssd1 vccd1 vccd1 _7142_/Y sky130_fd_sc_hd__nand2_1
X_4354_ _8137_/Q _4125_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _6024_/A vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__clkbuf_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _4285_/A vssd1 vssd1 vccd1 vccd1 _8163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7975_ _7975_/CLK _7975_/D vssd1 vssd1 vccd1 vccd1 _7975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6938_/A vssd1 vssd1 vccd1 vccd1 _6926_/X sky130_fd_sc_hd__buf_1
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5808_ _5808_/A vssd1 vssd1 vccd1 vccd1 _7647_/D sky130_fd_sc_hd__clkbuf_1
X_6832__414 _6833__415/A vssd1 vssd1 vccd1 vccd1 _8007_/CLK sky130_fd_sc_hd__inv_2
X_5739_ _7766_/Q _5567_/A _5741_/S vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7409_ _7409_/A _7409_/B _7409_/C _7409_/D vssd1 vssd1 vccd1 vccd1 _7410_/D sky130_fd_sc_hd__and4_1
XFILLER_2_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8389_ _8389_/CLK _8389_/D vssd1 vssd1 vccd1 vccd1 _8389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3399_ _7006_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3399_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_40 _7629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_51 _5916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7068__95 _7068__95/A vssd1 vssd1 vccd1 vccd1 _8192_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6961__509 _6961__509/A vssd1 vssd1 vccd1 vccd1 _8106_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _8052_/Q _8051_/Q _4536_/B vssd1 vssd1 vccd1 vccd1 _4070_/X sky130_fd_sc_hd__a21o_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7377__11 _7379__13/A vssd1 vssd1 vccd1 vccd1 _8313_/CLK sky130_fd_sc_hd__inv_2
X_4972_ _7940_/Q _7932_/Q _7924_/Q _7959_/Q _5198_/S _4971_/X vssd1 vssd1 vccd1 vccd1
+ _4972_/X sky130_fd_sc_hd__mux4_1
X_7760_ _7760_/CLK _7760_/D vssd1 vssd1 vccd1 vccd1 _7760_/Q sky130_fd_sc_hd__dfxtp_1
X_7691_ _8342_/CLK _7691_/D vssd1 vssd1 vccd1 vccd1 _7691_/Q sky130_fd_sc_hd__dfxtp_1
X_6711_ _8338_/Q vssd1 vssd1 vccd1 vccd1 _6711_/Y sky130_fd_sc_hd__inv_2
X_3923_ _3923_/A vssd1 vssd1 vccd1 vccd1 _8318_/D sky130_fd_sc_hd__clkbuf_1
X_3854_ _8378_/Q _3828_/X _3856_/S vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3785_ _8000_/Q _7999_/Q _7998_/Q vssd1 vssd1 vccd1 vccd1 _5249_/B sky130_fd_sc_hd__and3_1
X_8312_ _8312_/CLK _8312_/D vssd1 vssd1 vccd1 vccd1 _8312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5524_ _5524_/A vssd1 vssd1 vccd1 vccd1 _7879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5455_ _3840_/X _7909_/Q _5455_/S vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__mux2_1
X_8243_ _8243_/CLK _8243_/D vssd1 vssd1 vccd1 vccd1 _8243_/Q sky130_fd_sc_hd__dfxtp_1
X_4406_ _4406_/A vssd1 vssd1 vccd1 vccd1 _8117_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3253_ _6644_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3253_/X sky130_fd_sc_hd__clkbuf_16
X_8174_ _8174_/CLK _8174_/D vssd1 vssd1 vccd1 vccd1 _8174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7125_ _7125_/A _7134_/A _7125_/C vssd1 vssd1 vccd1 vccd1 _7230_/A sky130_fd_sc_hd__or3_1
X_5386_ _5401_/S vssd1 vssd1 vccd1 vccd1 _5395_/S sky130_fd_sc_hd__buf_2
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _4337_/A vssd1 vssd1 vccd1 vccd1 _8143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4268_ _5511_/B _5457_/B vssd1 vssd1 vccd1 vccd1 _4284_/S sky130_fd_sc_hd__nor2_4
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6007_ _6007_/A vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4199_ _4199_/A vssd1 vssd1 vccd1 vccd1 _8197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7958_ _7958_/CLK _7958_/D vssd1 vssd1 vccd1 vccd1 _7958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7889_ _7889_/CLK _7889_/D vssd1 vssd1 vccd1 vccd1 _7889_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6909_/A _6909_/B _6909_/C _6909_/D vssd1 vssd1 vccd1 vccd1 _6910_/B sky130_fd_sc_hd__nor4_1
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6466__246 _6467__247/A vssd1 vssd1 vccd1 vccd1 _7803_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _8171_/Q _7893_/Q _5240_/S vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ _8173_/Q _7895_/Q _5171_/S vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4144_/S vssd1 vssd1 vccd1 vccd1 _4135_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4053_ _7941_/Q _3814_/A _4052_/X _6350_/B vssd1 vssd1 vccd1 vccd1 _4844_/A sky130_fd_sc_hd__a31oi_4
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7812_ _7812_/CLK _7812_/D vssd1 vssd1 vccd1 vccd1 _7812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7743_ _7854_/CLK _7743_/D vssd1 vssd1 vccd1 vccd1 _7743_/Q sky130_fd_sc_hd__dfxtp_1
X_4955_ _4956_/A vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3906_ _3906_/A vssd1 vssd1 vccd1 vccd1 _8324_/D sky130_fd_sc_hd__clkbuf_1
X_7674_ _7991_/CLK _7674_/D vssd1 vssd1 vccd1 vccd1 _7674_/Q sky130_fd_sc_hd__dfxtp_1
X_4886_ _4886_/A vssd1 vssd1 vccd1 vccd1 _8041_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3406_ clkbuf_0__3406_/X vssd1 vssd1 vccd1 vccd1 _7043__75/A sky130_fd_sc_hd__clkbuf_4
X_3837_ _8359_/Q vssd1 vssd1 vccd1 vccd1 _3837_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6556_ _7861_/Q _5888_/A _6564_/S vssd1 vssd1 vccd1 vccd1 _6557_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5507_ _5304_/X _7886_/Q _5509_/S vssd1 vssd1 vccd1 vccd1 _5508_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8226_ _8364_/CLK _8226_/D vssd1 vssd1 vccd1 vccd1 _8226_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3199_ clkbuf_0__3199_/X vssd1 vssd1 vccd1 vccd1 _6496_/A sky130_fd_sc_hd__clkbuf_4
X_5438_ _5438_/A vssd1 vssd1 vccd1 vccd1 _7917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5369_ _7951_/Q _5366_/X _5377_/S vssd1 vssd1 vccd1 vccd1 _5370_/A sky130_fd_sc_hd__mux2_1
X_8157_ _8157_/CLK _8157_/D vssd1 vssd1 vccd1 vccd1 _8157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8088_ _8088_/CLK _8088_/D vssd1 vssd1 vccd1 vccd1 _8088_/Q sky130_fd_sc_hd__dfxtp_1
X_7108_ _8224_/Q _8223_/Q _8222_/Q _8221_/Q vssd1 vssd1 vccd1 vccd1 _7150_/D sky130_fd_sc_hd__and4_1
XFILLER_101_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7340__156 _7341__157/A vssd1 vssd1 vccd1 vccd1 _8283_/CLK sky130_fd_sc_hd__inv_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4863_/B _4708_/X _4713_/X _4739_/X vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__a31o_1
X_4671_ _4549_/X _4658_/X _4662_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4671_/X sky130_fd_sc_hd__a31o_1
X_6410_ _6422_/A vssd1 vssd1 vccd1 vccd1 _6410_/X sky130_fd_sc_hd__buf_1
X_6341_ _6341_/A _6341_/B _6341_/C _6341_/D vssd1 vssd1 vccd1 vccd1 _6909_/B sky130_fd_sc_hd__or4_4
X_6272_ _7715_/Q _6265_/X _6270_/X _7610_/A vssd1 vssd1 vccd1 vccd1 _7715_/D sky130_fd_sc_hd__a211o_1
XFILLER_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8011_ _8011_/CLK _8011_/D vssd1 vssd1 vccd1 vccd1 _8011_/Q sky130_fd_sc_hd__dfxtp_1
X_5223_ _5218_/X _5219_/X _5267_/A _5222_/X vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__a211o_1
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ _5154_/A _5154_/B _5154_/C vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__or3_1
XFILLER_110_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ _4105_/A vssd1 vssd1 vccd1 vccd1 _8264_/D sky130_fd_sc_hd__clkbuf_1
X_5085_ _8309_/Q _8301_/Q _8293_/Q _8317_/Q _5204_/S _4971_/A vssd1 vssd1 vccd1 vccd1
+ _5085_/X sky130_fd_sc_hd__mux4_2
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _8276_/Q _3951_/X _4036_/S vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7035__68 _7035__68/A vssd1 vssd1 vccd1 vccd1 _8165_/CLK sky130_fd_sc_hd__inv_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _5987_/A vssd1 vssd1 vccd1 vccd1 _5987_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7726_ _8391_/CLK _7726_/D vssd1 vssd1 vccd1 vccd1 _7726_/Q sky130_fd_sc_hd__dfxtp_1
X_4938_ _4938_/A vssd1 vssd1 vccd1 vccd1 _8019_/D sky130_fd_sc_hd__clkbuf_1
X_7657_ _7657_/CLK _7657_/D vssd1 vssd1 vccd1 vccd1 _7657_/Q sky130_fd_sc_hd__dfxtp_1
X_4869_ _4869_/A _4869_/B vssd1 vssd1 vccd1 vccd1 _4869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7588_ _7942_/Q _7618_/B vssd1 vssd1 vccd1 vccd1 _7602_/A sky130_fd_sc_hd__and2_1
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6539_ _6539_/A vssd1 vssd1 vccd1 vccd1 _7853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8209_ _8209_/CLK _8209_/D vssd1 vssd1 vccd1 vccd1 _8209_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput170 _6040_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput181 _6065_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput192 _6004_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3398_ clkbuf_0__3398_/X vssd1 vssd1 vccd1 vccd1 _7004__544/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7188__111 _7190__113/A vssd1 vssd1 vccd1 vccd1 _8210_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5910_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5910_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6890_ _6896_/A vssd1 vssd1 vccd1 vccd1 _6890_/X sky130_fd_sc_hd__buf_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5841_ _5841_/A vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5772_ _5772_/A vssd1 vssd1 vccd1 vccd1 _7707_/D sky130_fd_sc_hd__clkbuf_1
X_7511_ _7529_/B vssd1 vssd1 vccd1 vccd1 _7511_/X sky130_fd_sc_hd__clkbuf_2
X_6479__256 _6482__259/A vssd1 vssd1 vccd1 vccd1 _7813_/CLK sky130_fd_sc_hd__inv_2
X_4723_ _8078_/Q _4691_/X _4687_/X _8041_/Q vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__a22o_1
X_7442_ _7442_/A vssd1 vssd1 vccd1 vccd1 _7442_/Y sky130_fd_sc_hd__inv_2
X_4654_ _4332_/X _4538_/X _4653_/X _4609_/X vssd1 vssd1 vccd1 vccd1 _8062_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4585_ _4714_/A vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__buf_2
Xinput50 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__clkbuf_8
Xinput61 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _7584_/B sky130_fd_sc_hd__buf_4
Xinput72 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__buf_4
X_6324_ _6324_/A vssd1 vssd1 vccd1 vccd1 _6324_/X sky130_fd_sc_hd__clkbuf_2
Xinput83 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _7617_/A sky130_fd_sc_hd__buf_6
XFILLER_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6255_ _8058_/Q _6231_/X _6201_/X _6235_/X vssd1 vssd1 vccd1 vccd1 _6255_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5206_ _7934_/Q _5125_/X _4965_/A _5205_/X vssd1 vssd1 vccd1 vccd1 _5210_/B sky130_fd_sc_hd__o211a_1
X_6186_ _6189_/B _6186_/B _6188_/C vssd1 vssd1 vccd1 vccd1 _6187_/A sky130_fd_sc_hd__and3_1
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5137_ _8174_/Q _7896_/Q _5171_/S vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ _8254_/Q _8168_/Q _7906_/Q _8096_/Q _5042_/X _5220_/S vssd1 vssd1 vccd1 vccd1
+ _5068_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4019_ _4019_/A vssd1 vssd1 vccd1 vccd1 _8284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6423__211 _6424__212/A vssd1 vssd1 vccd1 vccd1 _7768_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3252_ clkbuf_0__3252_/X vssd1 vssd1 vccd1 vccd1 _6641__343/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7709_ _7709_/CLK _7709_/D vssd1 vssd1 vccd1 vccd1 _7709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7565__39 _7566__40/A vssd1 vssd1 vccd1 vccd1 _8378_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__3396_ clkbuf_0__3396_/X vssd1 vssd1 vccd1 vccd1 _6993__535/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6775__381 _6777__383/A vssd1 vssd1 vccd1 vccd1 _7966_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4249_/X _8130_/Q _4378_/S vssd1 vssd1 vccd1 vccd1 _4371_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6040_ _7679_/Q _6032_/X _6034_/X _6039_/X vssd1 vssd1 vccd1 vccd1 _6040_/X sky130_fd_sc_hd__o22a_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7991_ _7991_/CLK _7991_/D vssd1 vssd1 vccd1 vccd1 _7991_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7001__541 _7004__544/A vssd1 vssd1 vccd1 vccd1 _8138_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3723_ clkbuf_0__3723_/X vssd1 vssd1 vccd1 vccd1 _7572__45/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6897__461 _6898__462/A vssd1 vssd1 vccd1 vccd1 _8056_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8397_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5824_ _6164_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5825_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3585_ clkbuf_0__3585_/X vssd1 vssd1 vccd1 vccd1 _7307__130/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ _7759_/Q _5564_/A _5759_/S vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4706_ _4703_/X _7808_/Q _7648_/Q _4705_/X _4669_/S vssd1 vssd1 vccd1 vccd1 _4706_/X
+ sky130_fd_sc_hd__o221a_1
X_5686_ _5686_/A vssd1 vssd1 vccd1 vccd1 _7790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4637_ _7974_/Q _7966_/Q _7770_/Q _8035_/Q _4579_/X _4580_/X vssd1 vssd1 vccd1 vccd1
+ _4637_/X sky130_fd_sc_hd__mux4_2
X_7425_ _7425_/A _7425_/B _7425_/C _7425_/D vssd1 vssd1 vccd1 vccd1 _7425_/X sky130_fd_sc_hd__and4_1
XFILLER_116_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4568_ _4682_/B vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6307_ _6324_/A vssd1 vssd1 vccd1 vccd1 _6307_/X sky130_fd_sc_hd__clkbuf_2
X_4499_ _4338_/X _8078_/Q _4499_/S vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6238_ _6909_/A vssd1 vssd1 vccd1 vccd1 _6238_/Y sky130_fd_sc_hd__inv_2
X_6091__181 _6093__183/A vssd1 vssd1 vccd1 vccd1 _7650_/CLK sky130_fd_sc_hd__inv_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6169_/A vssd1 vssd1 vccd1 vccd1 _7694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8423__198 vssd1 vssd1 vccd1 vccd1 _8423__198/HI core0Index[5] sky130_fd_sc_hd__conb_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _3865_/X _8373_/Q _3882_/S vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3370_ clkbuf_0__3370_/X vssd1 vssd1 vccd1 vccd1 _6870__440/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540_ _5540_/A vssd1 vssd1 vccd1 vccd1 _7872_/D sky130_fd_sc_hd__clkbuf_1
X_5471_ _7902_/Q _4223_/A _5473_/S vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ _8112_/Q _4395_/X _4426_/S vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__mux2_1
X_7210_ _7218_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _8215_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8190_ _8190_/CLK _8190_/D vssd1 vssd1 vccd1 vccd1 _8190_/Q sky130_fd_sc_hd__dfxtp_1
X_7141_ _8406_/Q _7141_/B vssd1 vssd1 vccd1 vccd1 _7141_/Y sky130_fd_sc_hd__xnor2_1
X_4353_ _4353_/A vssd1 vssd1 vccd1 vccd1 _8138_/D sky130_fd_sc_hd__clkbuf_1
X_4284_ _8163_/Q _4143_/X _4284_/S vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__mux2_1
X_6023_ _7676_/Q _6022_/X _6023_/S vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__mux2_4
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7974_ _7974_/CLK _7974_/D vssd1 vssd1 vccd1 vccd1 _7974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _8292_/Q _3951_/X _3999_/S vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__mux2_1
X_5807_ _4093_/X _7647_/Q _5811_/S vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5738_ _5738_/A vssd1 vssd1 vccd1 vccd1 _7767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5669_ _5570_/X _7797_/Q _5669_/S vssd1 vssd1 vccd1 vccd1 _5670_/A sky130_fd_sc_hd__mux2_1
X_7408_ _6718_/Y _6719_/X _6735_/X _6737_/X _6739_/X vssd1 vssd1 vccd1 vccd1 _7409_/D
+ sky130_fd_sc_hd__o2111a_1
X_8388_ _8388_/CLK _8388_/D vssd1 vssd1 vccd1 vccd1 _8388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3398_ _7000_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3398_/X sky130_fd_sc_hd__clkbuf_16
X_7339_ _7339_/A vssd1 vssd1 vccd1 vccd1 _7339_/X sky130_fd_sc_hd__buf_1
X_7008__547 _7010__549/A vssd1 vssd1 vccd1 vccd1 _8144_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_41 _6554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_52 _6199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_30 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6579__294 _6580__295/A vssd1 vssd1 vccd1 vccd1 _7875_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6098__187 _6098__187/A vssd1 vssd1 vccd1 vccd1 _7656_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7304__127 _7306__129/A vssd1 vssd1 vccd1 vccd1 _8254_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7717_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4971_ _4971_/A vssd1 vssd1 vccd1 vccd1 _4971_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7690_ _8342_/CLK _7690_/D vssd1 vssd1 vccd1 vccd1 _7690_/Q sky130_fd_sc_hd__dfxtp_1
X_6710_ _8337_/Q _6744_/B _6720_/B vssd1 vssd1 vccd1 vccd1 _6716_/A sky130_fd_sc_hd__nand3_1
X_3922_ _3875_/X _8318_/Q _3926_/S vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _3853_/A vssd1 vssd1 vccd1 vccd1 _8379_/D sky130_fd_sc_hd__clkbuf_1
X_3784_ _8002_/Q _7997_/Q vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__xnor2_2
X_8311_ _8311_/CLK _8311_/D vssd1 vssd1 vccd1 vccd1 _8311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5523_ _7879_/Q _4220_/A _5527_/S vssd1 vssd1 vccd1 vccd1 _5524_/A sky130_fd_sc_hd__mux2_1
X_5454_ _5454_/A vssd1 vssd1 vccd1 vccd1 _7910_/D sky130_fd_sc_hd__clkbuf_1
X_8242_ _8242_/CLK _8242_/D vssd1 vssd1 vccd1 vccd1 _8242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4405_ _8117_/Q _4404_/X _4411_/S vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__mux2_1
X_5385_ _5385_/A _5421_/B vssd1 vssd1 vccd1 vccd1 _5401_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_0__3252_ _6638_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3252_/X sky130_fd_sc_hd__clkbuf_16
X_8173_ _8173_/CLK _8173_/D vssd1 vssd1 vccd1 vccd1 _8173_/Q sky130_fd_sc_hd__dfxtp_1
X_7124_ _8221_/Q vssd1 vssd1 vccd1 vccd1 _7125_/A sky130_fd_sc_hd__inv_2
X_4336_ _4335_/X _8143_/Q _4339_/S vssd1 vssd1 vccd1 vccd1 _4337_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7359__172 _7359__172/A vssd1 vssd1 vccd1 vccd1 _8299_/CLK sky130_fd_sc_hd__inv_2
X_4267_ _4267_/A vssd1 vssd1 vccd1 vccd1 _8171_/D sky130_fd_sc_hd__clkbuf_1
X_6006_ _7671_/Q _6005_/X _6006_/S vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__mux2_4
XFILLER_86_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4198_ _8197_/Q _4093_/X _4202_/S vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7957_ _7957_/CLK _7957_/D vssd1 vssd1 vccd1 vccd1 _7957_/Q sky130_fd_sc_hd__dfxtp_1
X_6908_ _6908_/A vssd1 vssd1 vccd1 vccd1 _8065_/D sky130_fd_sc_hd__clkbuf_1
X_7888_ _7888_/CLK _7888_/D vssd1 vssd1 vccd1 vccd1 _7888_/Q sky130_fd_sc_hd__dfxtp_1
X_6839_ _6346_/B _7535_/A _6839_/C vssd1 vssd1 vccd1 vccd1 _6840_/A sky130_fd_sc_hd__and3b_1
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7182__106 _7184__108/A vssd1 vssd1 vccd1 vccd1 _8205_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3361_ clkbuf_0__3361_/X vssd1 vssd1 vccd1 vccd1 _6844__420/A sky130_fd_sc_hd__clkbuf_16
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5170_ _7935_/Q _5151_/X _5017_/A _5169_/X vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__o211a_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4121_ _4121_/A _5457_/B vssd1 vssd1 vccd1 vccd1 _4144_/S sky130_fd_sc_hd__nor2_4
XFILLER_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4052_ _4052_/A _7536_/B _6214_/A vssd1 vssd1 vccd1 vccd1 _4052_/X sky130_fd_sc_hd__and3_1
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7047__77 _7048__78/A vssd1 vssd1 vccd1 vccd1 _8174_/CLK sky130_fd_sc_hd__inv_2
X_7811_ _7811_/CLK _7811_/D vssd1 vssd1 vccd1 vccd1 _7811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7742_ _7991_/CLK _7742_/D vssd1 vssd1 vccd1 vccd1 _7742_/Q sky130_fd_sc_hd__dfxtp_1
X_4954_ _8013_/Q vssd1 vssd1 vccd1 vccd1 _4956_/A sky130_fd_sc_hd__inv_2
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3905_ _3881_/X _8324_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3906_/A sky130_fd_sc_hd__mux2_1
X_7673_ _7991_/CLK _7673_/D vssd1 vssd1 vccd1 vccd1 _7673_/Q sky130_fd_sc_hd__dfxtp_1
X_4885_ _8041_/Q _4401_/X _4885_/S vssd1 vssd1 vccd1 vccd1 _4886_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3405_ clkbuf_0__3405_/X vssd1 vssd1 vccd1 vccd1 _7035__68/A sky130_fd_sc_hd__clkbuf_4
X_8415__237 vssd1 vssd1 vccd1 vccd1 partID[11] _8415__237/LO sky130_fd_sc_hd__conb_1
X_3836_ _3836_/A vssd1 vssd1 vccd1 vccd1 _8384_/D sky130_fd_sc_hd__clkbuf_1
X_6636__339 _6637__340/A vssd1 vssd1 vccd1 vccd1 _7920_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6555_ _6570_/S vssd1 vssd1 vccd1 vccd1 _6564_/S sky130_fd_sc_hd__clkbuf_2
X_5506_ _5506_/A vssd1 vssd1 vccd1 vccd1 _7887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8225_ _8335_/CLK _8225_/D vssd1 vssd1 vccd1 vccd1 _8225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3198_ clkbuf_0__3198_/X vssd1 vssd1 vccd1 vccd1 _6467__247/A sky130_fd_sc_hd__clkbuf_4
X_5437_ _7917_/Q _4529_/X _5437_/S vssd1 vssd1 vccd1 vccd1 _5438_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8156_ _8156_/CLK _8156_/D vssd1 vssd1 vccd1 vccd1 _8156_/Q sky130_fd_sc_hd__dfxtp_1
X_5368_ _5383_/S vssd1 vssd1 vccd1 vccd1 _5377_/S sky130_fd_sc_hd__buf_2
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7107_ _7150_/C vssd1 vssd1 vccd1 vccd1 _7159_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8087_ _8087_/CLK _8087_/D vssd1 vssd1 vccd1 vccd1 _8087_/Q sky130_fd_sc_hd__dfxtp_1
X_4319_ _8148_/Q _4140_/X _4321_/S vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__mux2_1
X_5299_ _7987_/Q vssd1 vssd1 vccd1 vccd1 _5564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7038_ _7038_/A vssd1 vssd1 vccd1 vccd1 _7038_/X sky130_fd_sc_hd__buf_1
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6891__456 _6893__458/A vssd1 vssd1 vccd1 vccd1 _8051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4664_/X _4666_/X _4669_/X _4588_/X _4674_/A vssd1 vssd1 vccd1 vccd1 _4670_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6340_ _8391_/Q _6340_/B vssd1 vssd1 vccd1 vccd1 _6346_/B sky130_fd_sc_hd__and2_1
X_6271_ _7600_/A vssd1 vssd1 vccd1 vccd1 _7610_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8010_ _8010_/CLK _8010_/D vssd1 vssd1 vccd1 vccd1 _8010_/Q sky130_fd_sc_hd__dfxtp_1
X_5222_ _5218_/A _5220_/X _5221_/X _5045_/A vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__o211a_1
X_5153_ _5148_/X _5149_/X _5152_/X _5084_/A vssd1 vssd1 vccd1 vccd1 _5154_/C sky130_fd_sc_hd__o211a_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4104_ _8264_/Q _3966_/X _4112_/S vssd1 vssd1 vccd1 vccd1 _4105_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5084_ _5084_/A _5084_/B vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__and2_1
X_4035_ _4035_/A vssd1 vssd1 vccd1 vccd1 _8277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _7665_/Q _5985_/X _5989_/S vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__mux2_1
X_7725_ _7991_/CLK _7725_/D vssd1 vssd1 vccd1 vccd1 _7725_/Q sky130_fd_sc_hd__dfxtp_1
X_4937_ _4332_/X _8019_/Q _4941_/S vssd1 vssd1 vccd1 vccd1 _4938_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4868_ _4703_/X _4865_/A _4867_/Y _4836_/X vssd1 vssd1 vccd1 vccd1 _8048_/D sky130_fd_sc_hd__o211a_1
X_7656_ _7656_/CLK _7656_/D vssd1 vssd1 vccd1 vccd1 _7656_/Q sky130_fd_sc_hd__dfxtp_1
X_3819_ _3841_/S vssd1 vssd1 vccd1 vccd1 _3832_/S sky130_fd_sc_hd__clkbuf_4
X_6607_ _6613_/A vssd1 vssd1 vccd1 vccd1 _6607_/X sky130_fd_sc_hd__buf_1
X_7587_ _7610_/A _7587_/B vssd1 vssd1 vccd1 vccd1 _8391_/D sky130_fd_sc_hd__nor2_1
X_4799_ _4730_/A _7962_/Q _7766_/Q _4731_/A vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6538_ _7584_/B _7853_/Q _6546_/S vssd1 vssd1 vccd1 vccd1 _6539_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8208_ _8208_/CLK _8208_/D vssd1 vssd1 vccd1 vccd1 _8208_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput160 _6075_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput171 _6043_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput182 _6067_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__buf_2
X_8139_ _8139_/CLK _8139_/D vssd1 vssd1 vccd1 vccd1 _8139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3397_ clkbuf_0__3397_/X vssd1 vssd1 vccd1 vccd1 _6998__539/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7367__3 _7369__5/A vssd1 vssd1 vccd1 vccd1 _8305_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5840_ _7536_/B _5844_/B vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__or2_1
XFILLER_22_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5771_ _5561_/X _7707_/Q _5771_/S vssd1 vssd1 vccd1 vccd1 _5772_/A sky130_fd_sc_hd__mux2_1
X_7510_ _7510_/A vssd1 vssd1 vccd1 vccd1 _7529_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7040__72 _7041__73/A vssd1 vssd1 vccd1 vccd1 _8169_/CLK sky130_fd_sc_hd__inv_2
X_4722_ _4715_/X _4718_/X _4721_/X vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__o21a_1
X_7441_ _7441_/A vssd1 vssd1 vccd1 vccd1 _8329_/D sky130_fd_sc_hd__clkbuf_1
X_4653_ _4540_/X _8062_/Q _4632_/X _4652_/X _4605_/X vssd1 vssd1 vccd1 vccd1 _4653_/X
+ sky130_fd_sc_hd__a221o_1
Xinput40 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__buf_4
X_4584_ _4601_/B _4584_/B vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__nor2_2
Xinput51 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__clkbuf_8
Xinput62 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _7579_/B sky130_fd_sc_hd__buf_4
Xinput73 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__buf_4
XFILLER_115_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6323_ _7724_/Q _6320_/X _6307_/X _6322_/X vssd1 vssd1 vccd1 vccd1 _7724_/D sky130_fd_sc_hd__a211o_1
Xinput84 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _7614_/B sky130_fd_sc_hd__buf_6
XFILLER_107_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6254_ _6342_/A _6254_/B _6249_/A vssd1 vssd1 vccd1 vccd1 _6254_/Y sky130_fd_sc_hd__nor3b_2
X_5205_ _7953_/Q _5126_/X _5148_/X _5204_/X vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__o22a_1
X_6185_ _7702_/Q _7701_/Q _6185_/C vssd1 vssd1 vccd1 vccd1 _6188_/C sky130_fd_sc_hd__or3_1
XFILLER_97_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5136_ _7936_/Q _5108_/B _5017_/A _5135_/X vssd1 vssd1 vccd1 vccd1 _5140_/B sky130_fd_sc_hd__o211a_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5067_ _5009_/X _5066_/X _5119_/A vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3251_ clkbuf_0__3251_/X vssd1 vssd1 vccd1 vccd1 _6637__340/A sky130_fd_sc_hd__clkbuf_4
X_4018_ _3881_/X _8284_/Q _4018_/S vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5969_ _6687_/A vssd1 vssd1 vccd1 vccd1 _7546_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7708_ _7708_/CLK _7708_/D vssd1 vssd1 vccd1 vccd1 _7708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7639_ _7642_/A _7639_/B vssd1 vssd1 vccd1 vccd1 _7640_/A sky130_fd_sc_hd__or2_1
XFILLER_119_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6573__289 _6574__290/A vssd1 vssd1 vccd1 vccd1 _7870_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8428__203 vssd1 vssd1 vccd1 vccd1 _8428__203/HI core1Index[3] sky130_fd_sc_hd__conb_1
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3395_ clkbuf_0__3395_/X vssd1 vssd1 vccd1 vccd1 _6985__528/A sky130_fd_sc_hd__clkbuf_16
XFILLER_85_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6485__261 _6487__263/A vssd1 vssd1 vccd1 vccd1 _7818_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7990_ _7991_/CLK _7990_/D vssd1 vssd1 vccd1 vccd1 _7990_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3722_ clkbuf_0__3722_/X vssd1 vssd1 vccd1 vccd1 _7564__38/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7353__167 _7355__169/A vssd1 vssd1 vccd1 vccd1 _8294_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823_ _5823_/A vssd1 vssd1 vccd1 vccd1 _5823_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3584_ clkbuf_0__3584_/X vssd1 vssd1 vccd1 vccd1 _7326_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5754_ _5754_/A vssd1 vssd1 vccd1 vccd1 _7760_/D sky130_fd_sc_hd__clkbuf_1
X_5685_ _7790_/Q _5593_/X _5687_/S vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__mux2_1
X_4705_ _4705_/A vssd1 vssd1 vccd1 vccd1 _4705_/X sky130_fd_sc_hd__buf_2
X_7424_ _7423_/B _7423_/C _8404_/Q vssd1 vssd1 vccd1 vccd1 _7425_/D sky130_fd_sc_hd__a21bo_1
X_4636_ _4867_/B _4633_/X _4635_/X vssd1 vssd1 vccd1 vccd1 _4636_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6306_ _7540_/B _6289_/A _6244_/X _6289_/B _6281_/A vssd1 vssd1 vccd1 vccd1 _6324_/A
+ sky130_fd_sc_hd__a41o_1
X_4567_ _4669_/S vssd1 vssd1 vccd1 vccd1 _4567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4498_ _4498_/A vssd1 vssd1 vccd1 vccd1 _8079_/D sky130_fd_sc_hd__clkbuf_1
X_7286_ _7286_/A vssd1 vssd1 vccd1 vccd1 _8240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6237_ _6237_/A _7732_/Q _6342_/B _6309_/A vssd1 vssd1 vccd1 vccd1 _6909_/C sky130_fd_sc_hd__or4b_1
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945__496 _6945__496/A vssd1 vssd1 vccd1 vccd1 _8093_/CLK sky130_fd_sc_hd__inv_2
X_6168_ _6199_/B _7694_/Q _6174_/S vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6906__469 _6906__469/A vssd1 vssd1 vccd1 vccd1 _8064_/CLK sky130_fd_sc_hd__inv_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5119_/A vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__buf_2
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7570__43 _7572__45/A vssd1 vssd1 vccd1 vccd1 _8382_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6100__189 _6101__190/A vssd1 vssd1 vccd1 vccd1 _7658_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7389__21 _7390__22/A vssd1 vssd1 vccd1 vccd1 _8323_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5470_ _5470_/A vssd1 vssd1 vccd1 vccd1 _7903_/D sky130_fd_sc_hd__clkbuf_1
X_4421_ _4421_/A vssd1 vssd1 vccd1 vccd1 _8113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7140_ _7204_/A _7140_/B vssd1 vssd1 vccd1 vccd1 _7141_/B sky130_fd_sc_hd__xor2_1
X_4352_ _8138_/Q _4229_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4283_ _4283_/A vssd1 vssd1 vccd1 vccd1 _8164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6022_ _7727_/Q input9/X _6025_/S vssd1 vssd1 vccd1 vccd1 _6022_/X sky130_fd_sc_hd__mux2_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7973_ _7973_/CLK _7973_/D vssd1 vssd1 vccd1 vccd1 _7973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6786_ _6786_/A vssd1 vssd1 vccd1 vccd1 _6786_/X sky130_fd_sc_hd__buf_1
X_5806_ _5806_/A vssd1 vssd1 vccd1 vccd1 _7648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ _3998_/A vssd1 vssd1 vccd1 vccd1 _8293_/D sky130_fd_sc_hd__clkbuf_1
X_5737_ _7767_/Q _5564_/A _5741_/S vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7407_ _7430_/A _6713_/A _6722_/Y _6723_/X vssd1 vssd1 vccd1 vccd1 _7409_/C sky130_fd_sc_hd__o2bb2a_1
X_5668_ _5668_/A vssd1 vssd1 vccd1 vccd1 _7798_/D sky130_fd_sc_hd__clkbuf_1
X_4619_ _8121_/Q _7891_/Q _7835_/Q _7795_/Q _4559_/A _4589_/X vssd1 vssd1 vccd1 vccd1
+ _4619_/X sky130_fd_sc_hd__mux4_1
X_8387_ _8387_/CLK _8387_/D vssd1 vssd1 vccd1 vccd1 _8387_/Q sky130_fd_sc_hd__dfxtp_1
X_5599_ _5599_/A _5617_/B vssd1 vssd1 vccd1 vccd1 _5615_/S sky130_fd_sc_hd__or2_2
XFILLER_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3397_ _6994_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3397_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7269_ _7285_/S vssd1 vssd1 vccd1 vccd1 _7269_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_42 _6185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_31 _5912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_20 _5905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_53 _7629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6436__222 _6437__223/A vssd1 vssd1 vccd1 vccd1 _7779_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6848__423 _6850__425/A vssd1 vssd1 vccd1 vccd1 _8018_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _5037_/A vssd1 vssd1 vccd1 vccd1 _4971_/A sky130_fd_sc_hd__buf_4
X_3921_ _3921_/A vssd1 vssd1 vccd1 vccd1 _8319_/D sky130_fd_sc_hd__clkbuf_1
X_6855__427 _6857__429/A vssd1 vssd1 vccd1 vccd1 _8022_/CLK sky130_fd_sc_hd__inv_2
X_3852_ _8379_/Q _3825_/X _3856_/S vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6571_ _6571_/A vssd1 vssd1 vccd1 vccd1 _7868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3783_ _7996_/Q vssd1 vssd1 vccd1 vccd1 _3783_/Y sky130_fd_sc_hd__inv_2
X_8310_ _8310_/CLK _8310_/D vssd1 vssd1 vccd1 vccd1 _8310_/Q sky130_fd_sc_hd__dfxtp_1
X_5522_ _5522_/A vssd1 vssd1 vccd1 vccd1 _7880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5453_ _3837_/X _7910_/Q _5455_/S vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8241_ _8241_/CLK _8241_/D vssd1 vssd1 vccd1 vccd1 _8241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8172_ _8172_/CLK _8172_/D vssd1 vssd1 vccd1 vccd1 _8172_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3251_ _6632_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3251_/X sky130_fd_sc_hd__clkbuf_16
X_5384_ _5384_/A vssd1 vssd1 vccd1 vccd1 _7944_/D sky130_fd_sc_hd__clkbuf_1
X_4404_ _7987_/Q vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__buf_2
XFILLER_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7123_ _7117_/X _7118_/Y _7121_/X _7122_/Y vssd1 vssd1 vccd1 vccd1 _7146_/C sky130_fd_sc_hd__o211a_1
X_4335_ _7989_/Q vssd1 vssd1 vccd1 vccd1 _4335_/X sky130_fd_sc_hd__clkbuf_2
X_6788__392 _6790__394/A vssd1 vssd1 vccd1 vccd1 _7977_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4266_ _4226_/X _8171_/Q _4266_/S vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__mux2_1
X_6005_ _7722_/Q input4/X _6008_/S vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__mux2_1
X_4197_ _4197_/A vssd1 vssd1 vccd1 vccd1 _8198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _7956_/CLK _7956_/D vssd1 vssd1 vccd1 vccd1 _7956_/Q sky130_fd_sc_hd__dfxtp_1
X_6907_ _7170_/A _7960_/Q _6907_/C vssd1 vssd1 vccd1 vccd1 _6908_/A sky130_fd_sc_hd__and3_1
XFILLER_23_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7887_ _7887_/CLK _7887_/D vssd1 vssd1 vccd1 vccd1 _7887_/Q sky130_fd_sc_hd__dfxtp_1
X_6838_ _6838_/A _7547_/B vssd1 vssd1 vccd1 vccd1 _7535_/A sky130_fd_sc_hd__and2_1
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7383__16 _7385__18/A vssd1 vssd1 vccd1 vccd1 _8318_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7310__132 _7311__133/A vssd1 vssd1 vccd1 vccd1 _8259_/CLK sky130_fd_sc_hd__inv_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4120_ _4286_/A _4286_/B _4120_/C vssd1 vssd1 vccd1 vccd1 _5457_/B sky130_fd_sc_hd__or3_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _4843_/B vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_7810_ _7810_/CLK _7810_/D vssd1 vssd1 vccd1 vccd1 _7810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7741_ _8365_/CLK _7741_/D vssd1 vssd1 vccd1 vccd1 _7741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7672_ _7992_/CLK _7672_/D vssd1 vssd1 vccd1 vccd1 _7672_/Q sky130_fd_sc_hd__dfxtp_1
X_3904_ _3904_/A vssd1 vssd1 vccd1 vccd1 _8325_/D sky130_fd_sc_hd__clkbuf_1
X_4884_ _4884_/A vssd1 vssd1 vccd1 vccd1 _8042_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3404_ clkbuf_0__3404_/X vssd1 vssd1 vccd1 vccd1 _7031__65/A sky130_fd_sc_hd__clkbuf_4
X_3835_ _8384_/Q _3834_/X _3841_/S vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__mux2_1
X_6554_ _6554_/A _6554_/B vssd1 vssd1 vccd1 vccd1 _6570_/S sky130_fd_sc_hd__and2_2
X_5505_ _5300_/X _7887_/Q _5509_/S vssd1 vssd1 vccd1 vccd1 _5506_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8224_ _8335_/CLK _8224_/D vssd1 vssd1 vccd1 vccd1 _8224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5436_ _5436_/A vssd1 vssd1 vccd1 vccd1 _7918_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3197_ clkbuf_0__3197_/X vssd1 vssd1 vccd1 vccd1 _6464__245/A sky130_fd_sc_hd__clkbuf_4
X_5367_ _5511_/A _5367_/B vssd1 vssd1 vccd1 vccd1 _5383_/S sky130_fd_sc_hd__nor2_2
X_8155_ _8155_/CLK _8155_/D vssd1 vssd1 vccd1 vccd1 _8155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7106_ _8220_/Q _8219_/Q _8218_/Q _8217_/Q vssd1 vssd1 vccd1 vccd1 _7150_/C sky130_fd_sc_hd__and4_1
X_5298_ _5298_/A vssd1 vssd1 vccd1 vccd1 _7980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8086_ _8086_/CLK _8086_/D vssd1 vssd1 vccd1 vccd1 _8086_/Q sky130_fd_sc_hd__dfxtp_1
X_4318_ _4318_/A vssd1 vssd1 vccd1 vccd1 _8149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _5025_/A vssd1 vssd1 vccd1 vccd1 _4249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _7939_/CLK _7939_/D vssd1 vssd1 vccd1 vccd1 _7939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6999__540 _6999__540/A vssd1 vssd1 vccd1 vccd1 _8137_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7052__81 _7056__85/A vssd1 vssd1 vccd1 vccd1 _8178_/CLK sky130_fd_sc_hd__inv_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ _6270_/A _6270_/B _6270_/C vssd1 vssd1 vccd1 vccd1 _6270_/X sky130_fd_sc_hd__and3_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _8099_/Q _5098_/X _5183_/A _8382_/Q vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o22a_1
X_5152_ _8101_/Q _5150_/X _5151_/X _8384_/Q vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4103_ _4118_/S vssd1 vssd1 vccd1 vccd1 _4112_/S sky130_fd_sc_hd__buf_2
XFILLER_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6449__232 _6451__234/A vssd1 vssd1 vccd1 vccd1 _7789_/CLK sky130_fd_sc_hd__inv_2
X_5083_ _8386_/Q _8325_/Q _8071_/Q _8103_/Q _5042_/X _5220_/S vssd1 vssd1 vccd1 vccd1
+ _5084_/B sky130_fd_sc_hd__mux4_1
X_7317__138 _7319__140/A vssd1 vssd1 vccd1 vccd1 _8265_/CLK sky130_fd_sc_hd__inv_2
X_4034_ _8277_/Q _3947_/X _4036_/S vssd1 vssd1 vccd1 vccd1 _4035_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6642__344 _6643__345/A vssd1 vssd1 vccd1 vccd1 _7925_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7724_ _7991_/CLK _7724_/D vssd1 vssd1 vccd1 vccd1 _7724_/Q sky130_fd_sc_hd__dfxtp_1
X_5985_ _7716_/Q input29/X _5991_/S vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__mux2_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4936_ _4936_/A vssd1 vssd1 vccd1 vccd1 _8020_/D sky130_fd_sc_hd__clkbuf_1
X_4867_ _4869_/A _4867_/B vssd1 vssd1 vccd1 vccd1 _4867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7655_ _7655_/CLK _7655_/D vssd1 vssd1 vccd1 vccd1 _7655_/Q sky130_fd_sc_hd__dfxtp_1
X_7586_ _7584_/Y _7585_/Y _7586_/S vssd1 vssd1 vccd1 vccd1 _7587_/B sky130_fd_sc_hd__mux2_1
X_3818_ _4507_/A _4121_/A vssd1 vssd1 vccd1 vccd1 _3841_/S sky130_fd_sc_hd__nor2_2
X_6537_ _6552_/S vssd1 vssd1 vccd1 vccd1 _6546_/S sky130_fd_sc_hd__clkbuf_2
X_4798_ _4729_/X _4796_/X _4797_/X vssd1 vssd1 vccd1 vccd1 _4802_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3249_ clkbuf_0__3249_/X vssd1 vssd1 vccd1 vccd1 _6625__330/A sky130_fd_sc_hd__clkbuf_4
Xoutput150 _5850_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__buf_2
X_6399_ _6399_/A vssd1 vssd1 vccd1 vccd1 _7753_/D sky130_fd_sc_hd__clkbuf_1
Xoutput161 _5972_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__buf_2
X_8207_ _8207_/CLK _8207_/D vssd1 vssd1 vccd1 vccd1 _8207_/Q sky130_fd_sc_hd__dfxtp_1
X_5419_ _7925_/Q _4529_/X _5419_/S vssd1 vssd1 vccd1 vccd1 _5420_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput183 _5981_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput172 _5977_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__buf_2
X_8138_ _8138_/CLK _8138_/D vssd1 vssd1 vccd1 vccd1 _8138_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3603_ clkbuf_0__3603_/X vssd1 vssd1 vccd1 vccd1 _7554__30/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8069_ _8069_/CLK _8069_/D vssd1 vssd1 vccd1 vccd1 _8069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7577__49 _7578__50/A vssd1 vssd1 vccd1 vccd1 _8388_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _5770_/A vssd1 vssd1 vccd1 vccd1 _7708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _8268_/Q _4719_/Y _4720_/X _8244_/Q _4556_/A vssd1 vssd1 vccd1 vccd1 _4721_/X
+ sky130_fd_sc_hd__o221a_1
X_7440_ _7519_/A _7440_/B _7442_/A vssd1 vssd1 vccd1 vccd1 _7441_/A sky130_fd_sc_hd__and3_1
X_4652_ _4549_/X _4636_/X _4640_/X _4651_/X vssd1 vssd1 vccd1 vccd1 _4652_/X sky130_fd_sc_hd__a31o_1
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
X_4583_ _8248_/Q _8146_/Q _7828_/Q _8272_/Q _4582_/X _4571_/X vssd1 vssd1 vccd1 vccd1
+ _4583_/X sky130_fd_sc_hd__mux4_1
Xinput41 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _5934_/A sky130_fd_sc_hd__buf_4
Xinput63 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _5875_/A sky130_fd_sc_hd__buf_4
Xinput52 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__buf_4
X_6322_ _7167_/A _6326_/B _6322_/C _6326_/D vssd1 vssd1 vccd1 vccd1 _6322_/X sky130_fd_sc_hd__and4_1
Xinput85 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _7611_/B sky130_fd_sc_hd__buf_6
Xinput74 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__buf_4
XFILLER_103_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6253_ _6253_/A vssd1 vssd1 vccd1 vccd1 _6253_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6980__525 _6980__525/A vssd1 vssd1 vccd1 vccd1 _8122_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5204_ _7918_/Q _7926_/Q _5204_/S vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__mux2_1
X_6184_ _7702_/Q _7701_/Q vssd1 vssd1 vccd1 vccd1 _6186_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5135_ _7955_/Q _5126_/X _5148_/A _5134_/X vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5066_ _8310_/Q _8302_/Q _8294_/Q _8318_/Q _5149_/S _4971_/A vssd1 vssd1 vccd1 vccd1
+ _5066_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3250_ clkbuf_0__3250_/X vssd1 vssd1 vccd1 vccd1 _6631__335/A sky130_fd_sc_hd__clkbuf_4
X_4017_ _4017_/A vssd1 vssd1 vccd1 vccd1 _8285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5968_ _7712_/Q input3/X _6052_/A vssd1 vssd1 vccd1 vccd1 _5968_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919_ _4919_/A vssd1 vssd1 vccd1 vccd1 _8027_/D sky130_fd_sc_hd__clkbuf_1
X_7707_ _7707_/CLK _7707_/D vssd1 vssd1 vccd1 vccd1 _7707_/Q sky130_fd_sc_hd__dfxtp_1
X_5899_ _5899_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5900_/A sky130_fd_sc_hd__or2_1
X_7638_ _8406_/Q _7533_/B _7641_/S vssd1 vssd1 vccd1 vccd1 _7639_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6430__217 _6432__219/A vssd1 vssd1 vccd1 vccd1 _7774_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6591__302 _6592__303/A vssd1 vssd1 vccd1 vccd1 _7883_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6782__387 _6782__387/A vssd1 vssd1 vccd1 vccd1 _7972_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3721_ clkbuf_0__3721_/X vssd1 vssd1 vccd1 vccd1 _7560__35/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6871_ _6871_/A vssd1 vssd1 vccd1 vccd1 _6871_/X sky130_fd_sc_hd__buf_1
X_5822_ _6185_/C _5826_/B vssd1 vssd1 vccd1 vccd1 _5823_/A sky130_fd_sc_hd__and2_1
XFILLER_50_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5753_ _7760_/Q _5561_/A _5753_/S vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__mux2_1
X_4704_ _4704_/A vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__clkbuf_2
X_5684_ _5684_/A vssd1 vssd1 vccd1 vccd1 _7791_/D sky130_fd_sc_hd__clkbuf_1
X_7423_ _7135_/A _7423_/B _7423_/C vssd1 vssd1 vccd1 vccd1 _7425_/C sky130_fd_sc_hd__nand3b_1
X_4635_ _4594_/X _4634_/X _4819_/A vssd1 vssd1 vccd1 vccd1 _4635_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8231_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4566_ _4726_/A vssd1 vssd1 vccd1 vccd1 _4669_/S sky130_fd_sc_hd__clkbuf_4
X_6305_ _6221_/X _6303_/X _6304_/X _6292_/X vssd1 vssd1 vccd1 vccd1 _7720_/D sky130_fd_sc_hd__a211o_1
X_4497_ _4335_/X _8079_/Q _4499_/S vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__mux2_1
X_7285_ _8240_/Q _7265_/B _7285_/S vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__mux2_1
X_6236_ _6236_/A vssd1 vssd1 vccd1 vccd1 _6350_/C sky130_fd_sc_hd__clkbuf_2
X_6167_ _6167_/A vssd1 vssd1 vccd1 vccd1 _7693_/D sky130_fd_sc_hd__clkbuf_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5191_/A _5112_/X _5117_/X vssd1 vssd1 vccd1 vccd1 _5118_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _8255_/Q _8169_/Q _7907_/Q _8097_/Q _5042_/X _5220_/S vssd1 vssd1 vccd1 vccd1
+ _5049_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6655__354 _6655__354/A vssd1 vssd1 vccd1 vccd1 _7935_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4420_ _8113_/Q _4392_/X _4426_/S vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4351_ _4366_/S vssd1 vssd1 vccd1 vccd1 _4360_/S sky130_fd_sc_hd__clkbuf_4
X_4282_ _8164_/Q _4140_/X _4284_/S vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6021_ _6021_/A vssd1 vssd1 vccd1 vccd1 _6021_/X sky130_fd_sc_hd__clkbuf_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7972_ _7972_/CLK _7972_/D vssd1 vssd1 vccd1 vccd1 _7972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6598__308 _6600__310/A vssd1 vssd1 vccd1 vccd1 _7889_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5805_ _4090_/X _7648_/Q _5805_/S vssd1 vssd1 vccd1 vccd1 _5806_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3997_ _8293_/Q _3947_/X _3999_/S vssd1 vssd1 vccd1 vccd1 _3998_/A sky130_fd_sc_hd__mux2_1
X_5736_ _5736_/A vssd1 vssd1 vccd1 vccd1 _7768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3603_ _7395_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3603_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5667_ _5567_/X _7798_/Q _5669_/S vssd1 vssd1 vccd1 vccd1 _5668_/A sky130_fd_sc_hd__mux2_1
X_7406_ _8394_/Q _7420_/B vssd1 vssd1 vccd1 vccd1 _7409_/B sky130_fd_sc_hd__xor2_1
X_4618_ _4567_/X _4615_/X _4617_/X vssd1 vssd1 vccd1 vccd1 _4618_/X sky130_fd_sc_hd__a21o_1
X_5598_ _5598_/A vssd1 vssd1 vccd1 vccd1 _7829_/D sky130_fd_sc_hd__clkbuf_1
X_8386_ _8386_/CLK _8386_/D vssd1 vssd1 vccd1 vccd1 _8386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _4549_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3396_ _6988_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3396_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_89_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7268_ _8232_/Q _7277_/B vssd1 vssd1 vccd1 vccd1 _7268_/X sky130_fd_sc_hd__or2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6219_ _6309_/A _6237_/A vssd1 vssd1 vccd1 vccd1 _7540_/B sky130_fd_sc_hd__nand2b_4
XFILLER_58_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_10 _8351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7199_ _7199_/A vssd1 vssd1 vccd1 vccd1 _7199_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_32 _5916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_43 _4211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 _5905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_54 _7546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6210__196 _6408__200/A vssd1 vssd1 vccd1 vccd1 _7708_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6993__535 _6993__535/A vssd1 vssd1 vccd1 vccd1 _8132_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7059__87 _7061__89/A vssd1 vssd1 vccd1 vccd1 _8184_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6443__227 _6443__227/A vssd1 vssd1 vccd1 vccd1 _7784_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _3872_/X _8319_/Q _3926_/S vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3851_ _3851_/A vssd1 vssd1 vccd1 vccd1 _8380_/D sky130_fd_sc_hd__clkbuf_1
X_6570_ _7868_/Q _5903_/A _6570_/S vssd1 vssd1 vccd1 vccd1 _6571_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3782_ _4949_/B _4949_/C _3782_/S vssd1 vssd1 vccd1 vccd1 _3793_/A sky130_fd_sc_hd__mux2_1
X_5521_ _7880_/Q _4217_/A _5521_/S vssd1 vssd1 vccd1 vccd1 _5522_/A sky130_fd_sc_hd__mux2_1
X_8240_ _8364_/CLK _8240_/D vssd1 vssd1 vccd1 vccd1 _8240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5452_ _5452_/A vssd1 vssd1 vccd1 vccd1 _7911_/D sky130_fd_sc_hd__clkbuf_1
X_4403_ _4403_/A vssd1 vssd1 vccd1 vccd1 _8118_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3250_ _6626_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3250_/X sky130_fd_sc_hd__clkbuf_16
X_5383_ _7944_/Q _4529_/X _5383_/S vssd1 vssd1 vccd1 vccd1 _5384_/A sky130_fd_sc_hd__mux2_1
X_8171_ _8171_/CLK _8171_/D vssd1 vssd1 vccd1 vccd1 _8171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7122_ _7234_/A _7234_/B _7612_/A vssd1 vssd1 vccd1 vccd1 _7122_/Y sky130_fd_sc_hd__o21ai_1
X_4334_ _4334_/A vssd1 vssd1 vccd1 vccd1 _8144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4265_ _4265_/A vssd1 vssd1 vccd1 vccd1 _8172_/D sky130_fd_sc_hd__clkbuf_1
X_6004_ _6004_/A vssd1 vssd1 vccd1 vccd1 _6004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4196_ _8198_/Q _4090_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6606__315 _6606__315/A vssd1 vssd1 vccd1 vccd1 _7896_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7955_ _7955_/CLK _7955_/D vssd1 vssd1 vccd1 vccd1 _7955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7886_ _7886_/CLK _7886_/D vssd1 vssd1 vccd1 vccd1 _7886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6498__272 _6500__274/A vssd1 vssd1 vccd1 vccd1 _7829_/CLK sky130_fd_sc_hd__inv_2
X_6768_ _6786_/A vssd1 vssd1 vccd1 vccd1 _6768_/X sky130_fd_sc_hd__buf_1
X_6699_ _8396_/Q _6699_/B vssd1 vssd1 vccd1 vccd1 _7410_/A sky130_fd_sc_hd__xor2_1
X_5719_ _7775_/Q _5590_/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__mux2_1
X_8369_ _8369_/CLK _8369_/D vssd1 vssd1 vccd1 vccd1 _8369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6507__279 _6507__279/A vssd1 vssd1 vccd1 vccd1 _7836_/CLK sky130_fd_sc_hd__inv_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6861__432 _6863__434/A vssd1 vssd1 vccd1 vccd1 _8027_/CLK sky130_fd_sc_hd__inv_2
X_4050_ _8051_/Q vssd1 vssd1 vccd1 vccd1 _4843_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _8012_/Q _7265_/A vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__and2_1
X_7740_ _8065_/CLK _7740_/D vssd1 vssd1 vccd1 vccd1 _7740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7671_ _7992_/CLK _7671_/D vssd1 vssd1 vccd1 vccd1 _7671_/Q sky130_fd_sc_hd__dfxtp_1
X_4883_ _8042_/Q _4398_/X _4885_/S vssd1 vssd1 vccd1 vccd1 _4884_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3903_ _3878_/X _8325_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3834_ _8360_/Q vssd1 vssd1 vccd1 vccd1 _3834_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6553_ _6553_/A vssd1 vssd1 vccd1 vccd1 _7860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5504_ _5504_/A vssd1 vssd1 vccd1 vccd1 _7888_/D sky130_fd_sc_hd__clkbuf_1
X_6484_ _6496_/A vssd1 vssd1 vccd1 vccd1 _6484_/X sky130_fd_sc_hd__buf_1
XFILLER_106_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8223_ _8223_/CLK _8223_/D vssd1 vssd1 vccd1 vccd1 _8223_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3196_ clkbuf_0__3196_/X vssd1 vssd1 vccd1 vccd1 _6457__239/A sky130_fd_sc_hd__clkbuf_4
X_5435_ _7918_/Q _4526_/X _5437_/S vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__mux2_1
X_8154_ _8154_/CLK _8154_/D vssd1 vssd1 vccd1 vccd1 _8154_/Q sky130_fd_sc_hd__dfxtp_1
X_5366_ _8365_/Q vssd1 vssd1 vccd1 vccd1 _5366_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7105_ _7150_/B vssd1 vssd1 vccd1 vccd1 _7159_/A sky130_fd_sc_hd__clkbuf_2
X_5297_ _5296_/X _7980_/Q _5297_/S vssd1 vssd1 vccd1 vccd1 _5298_/A sky130_fd_sc_hd__mux2_1
X_8085_ _8085_/CLK _8085_/D vssd1 vssd1 vccd1 vccd1 _8085_/Q sky130_fd_sc_hd__dfxtp_1
X_4317_ _8149_/Q _4137_/X _4321_/S vssd1 vssd1 vccd1 vccd1 _4318_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4248_ _4248_/A vssd1 vssd1 vccd1 vccd1 _8179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4179_ _8207_/Q _4093_/X _4183_/S vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7938_ _7938_/CLK _7938_/D vssd1 vssd1 vccd1 vccd1 _7938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7869_ _7869_/CLK _7869_/D vssd1 vssd1 vccd1 vccd1 _7869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _8321_/Q _8067_/Q _5220_/S vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _5151_/A vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _5367_/B _4204_/B vssd1 vssd1 vccd1 vccd1 _4118_/S sky130_fd_sc_hd__nor2_2
X_5082_ _4990_/X _5079_/X _5081_/X vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__a21o_1
X_4033_ _4033_/A vssd1 vssd1 vccd1 vccd1 _8278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7723_ _7991_/CLK _7723_/D vssd1 vssd1 vccd1 vccd1 _7723_/Q sky130_fd_sc_hd__dfxtp_1
X_5984_ _5984_/A vssd1 vssd1 vccd1 vccd1 _5984_/X sky130_fd_sc_hd__clkbuf_1
X_4935_ _4329_/X _8020_/Q _4941_/S vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4866_ _8049_/Q _4865_/A _4865_/Y _4774_/X vssd1 vssd1 vccd1 vccd1 _8049_/D sky130_fd_sc_hd__o211a_1
X_7654_ _7654_/CLK _7654_/D vssd1 vssd1 vccd1 vccd1 _7654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7585_ _8391_/Q vssd1 vssd1 vccd1 vccd1 _7585_/Y sky130_fd_sc_hd__clkinv_2
X_3817_ _5385_/A vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__clkbuf_4
X_4797_ _4724_/A _7758_/Q _4704_/A _8015_/Q _4621_/A vssd1 vssd1 vccd1 vccd1 _4797_/X
+ sky130_fd_sc_hd__o221a_1
X_8419__194 vssd1 vssd1 vccd1 vccd1 _8419__194/HI core0Index[1] sky130_fd_sc_hd__conb_1
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6536_ _6536_/A _6554_/B vssd1 vssd1 vccd1 vccd1 _6552_/S sky130_fd_sc_hd__nand2_2
XFILLER_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3248_ clkbuf_0__3248_/X vssd1 vssd1 vccd1 vccd1 _6644_/A sky130_fd_sc_hd__clkbuf_4
X_6868__438 _6868__438/A vssd1 vssd1 vccd1 vccd1 _8033_/CLK sky130_fd_sc_hd__inv_2
Xoutput140 _5894_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput151 _5852_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__buf_2
X_6398_ _7860_/Q _7753_/Q _6666_/S vssd1 vssd1 vccd1 vccd1 _6399_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8206_ _8206_/CLK _8206_/D vssd1 vssd1 vccd1 vccd1 _8206_/Q sky130_fd_sc_hd__dfxtp_1
X_5418_ _5418_/A vssd1 vssd1 vccd1 vccd1 _7926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5349_ _5364_/S vssd1 vssd1 vccd1 vccd1 _5358_/S sky130_fd_sc_hd__clkbuf_4
Xoutput184 _6069_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__buf_2
Xoutput162 _6007_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__buf_2
X_8137_ _8137_/CLK _8137_/D vssd1 vssd1 vccd1 vccd1 _8137_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput173 _6045_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3602_ clkbuf_0__3602_/X vssd1 vssd1 vccd1 vccd1 _7573_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8068_ _8068_/CLK _8068_/D vssd1 vssd1 vccd1 vccd1 _8068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7025__60 _7025__60/A vssd1 vssd1 vccd1 vccd1 _8157_/CLK sky130_fd_sc_hd__inv_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4720_ _4725_/A vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4651_ _4644_/X _4647_/X _4650_/X _4588_/X _4674_/A vssd1 vssd1 vccd1 vccd1 _4651_/X
+ sky130_fd_sc_hd__o221a_1
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__clkbuf_1
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
X_4582_ _4596_/A vssd1 vssd1 vccd1 vccd1 _4582_/X sky130_fd_sc_hd__buf_2
Xinput53 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _6349_/A sky130_fd_sc_hd__buf_8
Xinput42 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__buf_4
Xinput64 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__buf_4
X_7370_ _7388_/A vssd1 vssd1 vccd1 vccd1 _7370_/X sky130_fd_sc_hd__buf_1
X_6321_ _8395_/Q vssd1 vssd1 vccd1 vccd1 _7167_/A sky130_fd_sc_hd__clkbuf_4
Xinput75 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _5899_/A sky130_fd_sc_hd__buf_4
Xinput86 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _6164_/A sky130_fd_sc_hd__buf_8
XFILLER_107_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6252_ _8406_/Q _6249_/X _6251_/X _6228_/X vssd1 vssd1 vccd1 vccd1 _6252_/X sky130_fd_sc_hd__a31o_1
X_7323__143 _7325__145/A vssd1 vssd1 vccd1 vccd1 _8270_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6183_ _7702_/Q _6182_/X _6281_/A vssd1 vssd1 vccd1 vccd1 _6189_/B sky130_fd_sc_hd__o21ba_1
XFILLER_88_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5203_ _5271_/A _5201_/X _5202_/X vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _7920_/Q _7928_/Q _5237_/S vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _5084_/A _5065_/B vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__and2_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4016_ _3878_/X _8285_/Q _4018_/S vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5967_ _6029_/S vssd1 vssd1 vccd1 vccd1 _6052_/A sky130_fd_sc_hd__clkbuf_4
X_4918_ _8027_/Q _4395_/X _4922_/S vssd1 vssd1 vccd1 vccd1 _4919_/A sky130_fd_sc_hd__mux2_1
X_7706_ _7706_/CLK _7706_/D vssd1 vssd1 vccd1 vccd1 _7706_/Q sky130_fd_sc_hd__dfxtp_1
X_5898_ _5898_/A vssd1 vssd1 vccd1 vccd1 _5898_/X sky130_fd_sc_hd__clkbuf_1
X_7637_ _7637_/A vssd1 vssd1 vccd1 vccd1 _8405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4849_ _6801_/A vssd1 vssd1 vccd1 vccd1 _6907_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6915__472 _6918__475/A vssd1 vssd1 vccd1 vccd1 _8069_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6519_ _6534_/S vssd1 vssd1 vccd1 vccd1 _6528_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7499_ _7498_/Y _7450_/A _7402_/B _7510_/A _7490_/Y vssd1 vssd1 vccd1 vccd1 _7499_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5821_ _5821_/A vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3582_ clkbuf_0__3582_/X vssd1 vssd1 vccd1 vccd1 _7294__120/A sky130_fd_sc_hd__clkbuf_4
X_5752_ _5752_/A vssd1 vssd1 vccd1 vccd1 _7761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4703_ _4703_/A vssd1 vssd1 vccd1 vccd1 _4703_/X sky130_fd_sc_hd__clkbuf_4
X_5683_ _7791_/Q _5590_/X _5687_/S vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__mux2_1
X_7422_ _7422_/A _7422_/B vssd1 vssd1 vccd1 vccd1 _7425_/B sky130_fd_sc_hd__xnor2_1
X_4634_ _8088_/Q _8080_/Q _8043_/Q _8112_/Q _4569_/X _4571_/X vssd1 vssd1 vccd1 vccd1
+ _4634_/X sky130_fd_sc_hd__mux4_1
X_4565_ _4621_/A vssd1 vssd1 vccd1 vccd1 _4726_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6492__267 _6492__267/A vssd1 vssd1 vccd1 vccd1 _7824_/CLK sky130_fd_sc_hd__inv_2
X_6304_ _7720_/Q _7546_/C vssd1 vssd1 vccd1 vccd1 _6304_/X sky130_fd_sc_hd__and2_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4496_ _4496_/A vssd1 vssd1 vccd1 vccd1 _8080_/D sky130_fd_sc_hd__clkbuf_1
X_7284_ _8011_/Q _7266_/A _7283_/X _7178_/X vssd1 vssd1 vccd1 vccd1 _8239_/D sky130_fd_sc_hd__o211a_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6235_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6166_ _6687_/B _7693_/Q _6174_/S vssd1 vssd1 vccd1 vccd1 _6167_/A sky130_fd_sc_hd__mux2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _8316_/Q _5114_/X _5183_/A _8308_/Q _5123_/S vssd1 vssd1 vccd1 vccd1 _5117_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5048_ _5171_/S vssd1 vssd1 vccd1 vccd1 _5220_/S sky130_fd_sc_hd__buf_4
X_7074__100 _7073__99/A vssd1 vssd1 vccd1 vccd1 _8197_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4350_ _5367_/B _4368_/B vssd1 vssd1 vccd1 vccd1 _4366_/S sky130_fd_sc_hd__nor2_4
XFILLER_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4281_ _4281_/A vssd1 vssd1 vccd1 vccd1 _8165_/D sky130_fd_sc_hd__clkbuf_1
X_6020_ _7675_/Q _6019_/X _6023_/S vssd1 vssd1 vccd1 vccd1 _6021_/A sky130_fd_sc_hd__mux2_4
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7971_ _7971_/CLK _7971_/D vssd1 vssd1 vccd1 vccd1 _7971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6853_ _6877_/A vssd1 vssd1 vccd1 vccd1 _6853_/X sky130_fd_sc_hd__buf_1
X_5804_ _5804_/A vssd1 vssd1 vccd1 vccd1 _7649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3996_ _3996_/A vssd1 vssd1 vccd1 vccd1 _8294_/D sky130_fd_sc_hd__clkbuf_1
X_5735_ _7768_/Q _5561_/A _5735_/S vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__mux2_1
X_6500__274 _6500__274/A vssd1 vssd1 vccd1 vccd1 _7831_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3602_ _7394_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3602_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5666_ _5666_/A vssd1 vssd1 vccd1 vccd1 _7799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7405_ _6747_/X _6749_/Y _6754_/Y _7404_/X _6743_/B vssd1 vssd1 vccd1 vccd1 _7410_/C
+ sky130_fd_sc_hd__o2111a_1
X_4617_ _4557_/A _4616_/X _4714_/A vssd1 vssd1 vccd1 vccd1 _4617_/X sky130_fd_sc_hd__a21o_1
X_5597_ _7829_/Q _5596_/X _5597_/S vssd1 vssd1 vccd1 vccd1 _5598_/A sky130_fd_sc_hd__mux2_1
X_8385_ _8385_/CLK _8385_/D vssd1 vssd1 vccd1 vccd1 _8385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4548_ _8050_/Q _4601_/B vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__xor2_2
XFILLER_2_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3395_ _6982_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3395_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _4479_/A vssd1 vssd1 vccd1 vccd1 _8087_/D sky130_fd_sc_hd__clkbuf_1
X_7267_ _7283_/B vssd1 vssd1 vccd1 vccd1 _7277_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6218_ _7754_/Q vssd1 vssd1 vccd1 vccd1 _6237_/A sky130_fd_sc_hd__clkbuf_2
X_7198_ _7222_/A vssd1 vssd1 vccd1 vccd1 _7198_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6149_ _6145_/X _7859_/Q _6142_/X _6146_/X _7683_/Q vssd1 vssd1 vccd1 vccd1 _7683_/D
+ sky130_fd_sc_hd__o32a_1
XINSDIODE2_11 _6040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_33 _5916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_22 _5905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_55 _5914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_44 _4217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7336__153 _7336__153/A vssd1 vssd1 vccd1 vccd1 _8280_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6928__482 _6928__482/A vssd1 vssd1 vccd1 vccd1 _8079_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3850_ _8380_/Q _3822_/X _3856_/S vssd1 vssd1 vccd1 vccd1 _3851_/A sky130_fd_sc_hd__mux2_1
X_3781_ _3867_/A _7994_/Q vssd1 vssd1 vccd1 vccd1 _3782_/S sky130_fd_sc_hd__xnor2_1
X_5520_ _5520_/A vssd1 vssd1 vccd1 vccd1 _7881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5451_ _3834_/X _7911_/Q _5455_/S vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__mux2_1
X_4402_ _8118_/Q _4401_/X _4402_/S vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__mux2_1
X_5382_ _5382_/A vssd1 vssd1 vccd1 vccd1 _7945_/D sky130_fd_sc_hd__clkbuf_1
X_8170_ _8170_/CLK _8170_/D vssd1 vssd1 vccd1 vccd1 _8170_/Q sky130_fd_sc_hd__dfxtp_1
X_7121_ _8398_/Q _7234_/A _7234_/B vssd1 vssd1 vccd1 vccd1 _7121_/X sky130_fd_sc_hd__or3_1
X_4333_ _4332_/X _8144_/Q _4339_/S vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4264_ _4223_/X _8172_/Q _4266_/S vssd1 vssd1 vccd1 vccd1 _4265_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6003_ _7670_/Q _6002_/X _6006_/S vssd1 vssd1 vccd1 vccd1 _6004_/A sky130_fd_sc_hd__mux2_4
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4195_ _4195_/A vssd1 vssd1 vccd1 vccd1 _8199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7954_ _7954_/CLK _7954_/D vssd1 vssd1 vccd1 vccd1 _7954_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7885_ _7885_/CLK _7885_/D vssd1 vssd1 vccd1 vccd1 _7885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6795__398 _6796__399/A vssd1 vssd1 vccd1 vccd1 _7983_/CLK sky130_fd_sc_hd__inv_2
X_6767_ _6815_/A vssd1 vssd1 vccd1 vccd1 _6767_/X sky130_fd_sc_hd__buf_1
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5718_ _5718_/A vssd1 vssd1 vccd1 vccd1 _7776_/D sky130_fd_sc_hd__clkbuf_1
X_3979_ _3979_/A vssd1 vssd1 vccd1 vccd1 _8301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6698_ _8342_/Q _6694_/X _6705_/B vssd1 vssd1 vccd1 vccd1 _6699_/B sky130_fd_sc_hd__o21bai_2
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5649_ _7806_/Q _5593_/X _5651_/S vssd1 vssd1 vccd1 vccd1 _5650_/A sky130_fd_sc_hd__mux2_1
X_8368_ _8368_/CLK _8368_/D vssd1 vssd1 vccd1 vccd1 _8368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8299_ _8299_/CLK _8299_/D vssd1 vssd1 vccd1 vccd1 _8299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7064__91 _7066__93/A vssd1 vssd1 vccd1 vccd1 _8188_/CLK sky130_fd_sc_hd__inv_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _6841_/C vssd1 vssd1 vccd1 vccd1 _7265_/A sky130_fd_sc_hd__inv_2
X_7670_ _7992_/CLK _7670_/D vssd1 vssd1 vccd1 vccd1 _7670_/Q sky130_fd_sc_hd__dfxtp_1
X_4882_ _4882_/A vssd1 vssd1 vccd1 vccd1 _8043_/D sky130_fd_sc_hd__clkbuf_1
X_3902_ _3902_/A vssd1 vssd1 vccd1 vccd1 _8326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3833_ _3833_/A vssd1 vssd1 vccd1 vccd1 _8385_/D sky130_fd_sc_hd__clkbuf_1
X_6552_ _5886_/A _7860_/Q _6552_/S vssd1 vssd1 vccd1 vccd1 _6553_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5503_ _5296_/X _7888_/Q _5503_/S vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__mux2_1
X_8222_ _8223_/CLK _8222_/D vssd1 vssd1 vccd1 vccd1 _8222_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3195_ clkbuf_0__3195_/X vssd1 vssd1 vccd1 vccd1 _6452__235/A sky130_fd_sc_hd__clkbuf_4
X_5434_ _5434_/A vssd1 vssd1 vccd1 vccd1 _7919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8153_ _8153_/CLK _8153_/D vssd1 vssd1 vccd1 vccd1 _8153_/Q sky130_fd_sc_hd__dfxtp_1
X_6612__320 _6612__320/A vssd1 vssd1 vccd1 vccd1 _7901_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7104_ _7104_/A _7104_/B _7104_/C _7104_/D vssd1 vssd1 vccd1 vccd1 _7104_/X sky130_fd_sc_hd__or4_1
X_5365_ _5365_/A vssd1 vssd1 vccd1 vccd1 _7952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5296_ _5561_/A vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__clkbuf_2
X_4316_ _4316_/A vssd1 vssd1 vccd1 vccd1 _8150_/D sky130_fd_sc_hd__clkbuf_1
X_8084_ _8084_/CLK _8084_/D vssd1 vssd1 vccd1 vccd1 _8084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4247_ _8179_/Q _4143_/X _4247_/S vssd1 vssd1 vccd1 vccd1 _4248_/A sky130_fd_sc_hd__mux2_1
X_4178_ _4178_/A vssd1 vssd1 vccd1 vccd1 _8208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7937_ _7937_/CLK _7937_/D vssd1 vssd1 vccd1 vccd1 _7937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7868_ _8342_/CLK _7868_/D vssd1 vssd1 vccd1 vccd1 _7868_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7799_ _7799_/CLK _7799_/D vssd1 vssd1 vccd1 vccd1 _7799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6513__284 _6514__285/A vssd1 vssd1 vccd1 vccd1 _7841_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5150_ _5150_/A vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__buf_2
X_4101_ _4101_/A vssd1 vssd1 vccd1 vccd1 _8265_/D sky130_fd_sc_hd__clkbuf_1
X_5081_ _5009_/X _5080_/X _5154_/A vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _8278_/Q _3943_/X _4036_/S vssd1 vssd1 vccd1 vccd1 _4033_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5983_ _7664_/Q _5982_/X _5989_/S vssd1 vssd1 vccd1 vccd1 _5984_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7722_ _7992_/CLK _7722_/D vssd1 vssd1 vccd1 vccd1 _7722_/Q sky130_fd_sc_hd__dfxtp_1
X_4934_ _4934_/A vssd1 vssd1 vccd1 vccd1 _8021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8332_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4865_ _4865_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4865_/Y sky130_fd_sc_hd__nand2_1
X_7653_ _7653_/CLK _7653_/D vssd1 vssd1 vccd1 vccd1 _7653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7584_ _7608_/A _7584_/B vssd1 vssd1 vccd1 vccd1 _7584_/Y sky130_fd_sc_hd__nand2_1
X_3816_ _3867_/A _5262_/A _3967_/A vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__or3b_4
X_4796_ _4730_/X _7870_/Q _7774_/Q _4731_/X vssd1 vssd1 vccd1 vccd1 _4796_/X sky130_fd_sc_hd__a22o_1
X_6456__238 _6457__239/A vssd1 vssd1 vccd1 vccd1 _7795_/CLK sky130_fd_sc_hd__inv_2
X_6535_ _6535_/A vssd1 vssd1 vccd1 vccd1 _7852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3247_ clkbuf_0__3247_/X vssd1 vssd1 vccd1 vccd1 _6615__322/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8205_ _8205_/CLK _8205_/D vssd1 vssd1 vccd1 vccd1 _8205_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput141 _5896_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput130 _5874_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput152 _5854_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__buf_2
X_6397_ _6397_/A vssd1 vssd1 vccd1 vccd1 _7752_/D sky130_fd_sc_hd__clkbuf_1
X_5417_ _7926_/Q _4526_/X _5419_/S vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__mux2_1
X_5348_ _5348_/A _5421_/B vssd1 vssd1 vccd1 vccd1 _5364_/S sky130_fd_sc_hd__or2_2
Xoutput185 _6071_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput163 _6011_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__buf_2
X_8136_ _8136_/CLK _8136_/D vssd1 vssd1 vccd1 vccd1 _8136_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput174 _6047_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3601_ clkbuf_0__3601_/X vssd1 vssd1 vccd1 vccd1 _7393__25/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8067_ _8067_/CLK _8067_/D vssd1 vssd1 vccd1 vccd1 _8067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5279_ _5548_/A _5653_/B vssd1 vssd1 vccd1 vccd1 _5309_/S sky130_fd_sc_hd__or2_2
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3394_ clkbuf_0__3394_/X vssd1 vssd1 vccd1 vccd1 _7000_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8451__226 vssd1 vssd1 vccd1 vccd1 _8451__226/HI versionID[0] sky130_fd_sc_hd__conb_1
X_4650_ _4648_/X _4649_/X _4650_/S vssd1 vssd1 vccd1 vccd1 _4650_/X sky130_fd_sc_hd__mux2_1
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__clkbuf_1
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
X_6320_ _6320_/A vssd1 vssd1 vccd1 vccd1 _6320_/X sky130_fd_sc_hd__clkbuf_2
X_4581_ _8090_/Q _8082_/Q _8045_/Q _8114_/Q _4579_/X _4580_/X vssd1 vssd1 vccd1 vccd1
+ _4581_/X sky130_fd_sc_hd__mux4_2
Xinput54 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _6687_/B sky130_fd_sc_hd__clkbuf_16
Xinput43 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput87 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _6518_/A sky130_fd_sc_hd__buf_6
Xinput65 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _6199_/B sky130_fd_sc_hd__clkbuf_16
Xinput76 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _7536_/B sky130_fd_sc_hd__buf_8
X_6251_ _6301_/B vssd1 vssd1 vccd1 vccd1 _6251_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6182_ _6349_/A _7540_/A _6349_/C _7701_/Q vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__a31o_1
X_5202_ _8367_/Q _5187_/X _5183_/X _8375_/Q _4988_/X vssd1 vssd1 vccd1 vccd1 _5202_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5133_ _5218_/A _5131_/X _5132_/X vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5064_ _8387_/Q _8326_/Q _8072_/Q _8104_/Q _5042_/X _5234_/S vssd1 vssd1 vccd1 vccd1
+ _5065_/B sky130_fd_sc_hd__mux4_1
X_4015_ _4015_/A vssd1 vssd1 vccd1 vccd1 _8286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5966_/A vssd1 vssd1 vccd1 vccd1 _6029_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_80_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6874__443 _6876__445/A vssd1 vssd1 vccd1 vccd1 _8038_/CLK sky130_fd_sc_hd__inv_2
X_5897_ _5897_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__or2_1
X_4917_ _4917_/A vssd1 vssd1 vccd1 vccd1 _8028_/D sky130_fd_sc_hd__clkbuf_1
X_6835__416 _6837__418/A vssd1 vssd1 vccd1 vccd1 _8009_/CLK sky130_fd_sc_hd__inv_2
X_7705_ _7705_/CLK _7705_/D vssd1 vssd1 vccd1 vccd1 _7705_/Q sky130_fd_sc_hd__dfxtp_1
X_7636_ _7642_/A _7636_/B vssd1 vssd1 vccd1 vccd1 _7637_/A sky130_fd_sc_hd__or2_1
X_4848_ _4930_/A _4836_/X _4851_/B _5785_/S vssd1 vssd1 vccd1 vccd1 _8055_/D sky130_fd_sc_hd__a31o_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7567_ _7573_/A vssd1 vssd1 vccd1 vccd1 _7567_/X sky130_fd_sc_hd__buf_1
X_4779_ _4697_/X _7705_/Q _7654_/Q _4699_/X vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__a22o_1
X_6518_ _6518_/A _6554_/B vssd1 vssd1 vccd1 vccd1 _6534_/S sky130_fd_sc_hd__nand2_2
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7498_ _7498_/A vssd1 vssd1 vccd1 vccd1 _7498_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8119_ _8119_/CLK _8119_/D vssd1 vssd1 vccd1 vccd1 _8119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6625__330 _6625__330/A vssd1 vssd1 vccd1 vccd1 _7911_/CLK sky130_fd_sc_hd__inv_2
X_6922__477 _6922__477/A vssd1 vssd1 vccd1 vccd1 _8074_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3377_ clkbuf_0__3377_/X vssd1 vssd1 vccd1 vccd1 _6912__470/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5820_ _6349_/C _5826_/B vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__and2_1
X_5751_ _7761_/Q _5558_/A _5753_/S vssd1 vssd1 vccd1 vccd1 _5752_/A sky130_fd_sc_hd__mux2_1
X_4702_ _4724_/A vssd1 vssd1 vccd1 vccd1 _4703_/A sky130_fd_sc_hd__clkbuf_2
X_7421_ _7421_/A _7447_/A vssd1 vssd1 vccd1 vccd1 _7422_/B sky130_fd_sc_hd__xor2_1
X_5682_ _5682_/A vssd1 vssd1 vccd1 vccd1 _7792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _8246_/Q _8144_/Q _7826_/Q _8270_/Q _4872_/A _4562_/X vssd1 vssd1 vccd1 vccd1
+ _4633_/X sky130_fd_sc_hd__mux4_1
X_4564_ _4564_/A _4675_/A vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__nor2_1
X_6303_ _6289_/X _6299_/X _6301_/X _7615_/A vssd1 vssd1 vccd1 vccd1 _6303_/X sky130_fd_sc_hd__a22o_1
X_7283_ _8239_/Q _7283_/B vssd1 vssd1 vccd1 vccd1 _7283_/X sky130_fd_sc_hd__or2_1
XFILLER_104_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4495_ _4332_/X _8080_/Q _4499_/S vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__mux2_1
X_6234_ _6234_/A _6285_/B _6342_/A _6343_/B vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__or4b_1
XFILLER_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6165_ _6180_/S vssd1 vssd1 vccd1 vccd1 _6174_/S sky130_fd_sc_hd__buf_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6096_/A vssd1 vssd1 vccd1 vccd1 _6096_/X sky130_fd_sc_hd__buf_1
X_5116_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5047_ _5009_/X _5046_/X _5119_/A vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5949_ _7857_/Q _5953_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__and2_1
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7619_ _7641_/S vssd1 vssd1 vccd1 vccd1 _7635_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7081__105 _7081__105/A vssd1 vssd1 vccd1 vccd1 _8202_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6413__203 _6413__203/A vssd1 vssd1 vccd1 vccd1 _7760_/CLK sky130_fd_sc_hd__inv_2
X_4280_ _8165_/Q _4137_/X _4284_/S vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7970_ _7970_/CLK _7970_/D vssd1 vssd1 vccd1 vccd1 _7970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6852_ _6883_/A vssd1 vssd1 vccd1 vccd1 _6852_/X sky130_fd_sc_hd__buf_1
XFILLER_35_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5803_ _4087_/X _7649_/Q _5805_/S vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__mux2_1
X_3995_ _8294_/Q _3943_/X _3999_/S vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3601_ _7388_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3601_/X sky130_fd_sc_hd__clkbuf_16
X_5734_ _5734_/A vssd1 vssd1 vccd1 vccd1 _7769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5665_ _5564_/X _7799_/Q _5669_/S vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__mux2_1
X_7404_ _7430_/A _6713_/A _6742_/C _6742_/A vssd1 vssd1 vccd1 vccd1 _7404_/X sky130_fd_sc_hd__o211a_1
X_4616_ _8247_/Q _8145_/Q _7827_/Q _8271_/Q _4582_/X _4580_/A vssd1 vssd1 vccd1 vccd1
+ _4616_/X sky130_fd_sc_hd__mux4_1
X_8384_ _8384_/CLK _8384_/D vssd1 vssd1 vccd1 vccd1 _8384_/Q sky130_fd_sc_hd__dfxtp_1
X_5596_ _7985_/Q vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4547_ _4547_/A vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__buf_2
Xclkbuf_0__3394_ _6981_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3394_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4478_ _4335_/X _8087_/Q _4480_/S vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__mux2_1
X_7266_ _7266_/A vssd1 vssd1 vccd1 vccd1 _7266_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6217_ _7755_/Q vssd1 vssd1 vccd1 vccd1 _6309_/A sky130_fd_sc_hd__clkbuf_2
X_7197_ _7202_/B _7192_/Y vssd1 vssd1 vccd1 vccd1 _7222_/A sky130_fd_sc_hd__or2b_2
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6148_ _6145_/X _7858_/Q _6142_/X _6146_/X _7682_/Q vssd1 vssd1 vccd1 vccd1 _7682_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_34 _5918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_23 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_12 _6040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_56 _7546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6079_ _7600_/A _6349_/D _6349_/A _6079_/D vssd1 vssd1 vccd1 vccd1 _6080_/A sky130_fd_sc_hd__and4b_1
XINSDIODE2_45 _5227_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6887__453 _6888__454/A vssd1 vssd1 vccd1 vccd1 _8048_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3780_ _7998_/Q _7993_/Q vssd1 vssd1 vccd1 vccd1 _4949_/C sky130_fd_sc_hd__and2b_1
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5450_ _5450_/A vssd1 vssd1 vccd1 vccd1 _7912_/D sky130_fd_sc_hd__clkbuf_1
X_4401_ _7988_/Q vssd1 vssd1 vccd1 vccd1 _4401_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5381_ _7945_/Q _4526_/X _5383_/S vssd1 vssd1 vccd1 vccd1 _5382_/A sky130_fd_sc_hd__mux2_1
X_4332_ _7990_/Q vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__clkbuf_2
X_7120_ _8221_/Q _7159_/A _7159_/B _8222_/Q vssd1 vssd1 vccd1 vccd1 _7234_/B sky130_fd_sc_hd__a31oi_2
XFILLER_113_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7051_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7051_/X sky130_fd_sc_hd__buf_1
X_4263_ _4263_/A vssd1 vssd1 vccd1 vccd1 _8173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6002_ _7721_/Q input34/X _6008_/S vssd1 vssd1 vccd1 vccd1 _6002_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4194_ _8199_/Q _4087_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7953_ _7953_/CLK _7953_/D vssd1 vssd1 vccd1 vccd1 _7953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7884_ _7884_/CLK _7884_/D vssd1 vssd1 vccd1 vccd1 _7884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _6766_/A vssd1 vssd1 vccd1 vccd1 _7960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3978_ _8301_/Q _3947_/X _3980_/S vssd1 vssd1 vccd1 vccd1 _3979_/A sky130_fd_sc_hd__mux2_1
X_5717_ _7776_/Q _5587_/X _5717_/S vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6697_ _6738_/B _6744_/C _6744_/D vssd1 vssd1 vccd1 vccd1 _6705_/B sky130_fd_sc_hd__and3_1
X_5648_ _5648_/A vssd1 vssd1 vccd1 vccd1 _7807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5579_ _7835_/Q _5578_/X _5588_/S vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__mux2_1
X_8367_ _8367_/CLK _8367_/D vssd1 vssd1 vccd1 vccd1 _8367_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3377_ _6902_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3377_/X sky130_fd_sc_hd__clkbuf_16
X_8298_ _8298_/CLK _8298_/D vssd1 vssd1 vccd1 vccd1 _8298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7249_ _7251_/A _7249_/B vssd1 vssd1 vccd1 vccd1 _8227_/D sky130_fd_sc_hd__nor2_1
XFILLER_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6976__521 _6977__522/A vssd1 vssd1 vccd1 vccd1 _8118_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _4949_/X _4950_/B _4950_/C vssd1 vssd1 vccd1 vccd1 _6841_/C sky130_fd_sc_hd__nand3b_4
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4881_ _8043_/Q _4395_/X _4885_/S vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__mux2_1
X_3901_ _3875_/X _8326_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3401_ clkbuf_0__3401_/X vssd1 vssd1 vccd1 vccd1 _7038_/A sky130_fd_sc_hd__clkbuf_4
X_6620_ _6632_/A vssd1 vssd1 vccd1 vccd1 _6620_/X sky130_fd_sc_hd__buf_1
X_3832_ _8385_/Q _3831_/X _3832_/S vssd1 vssd1 vccd1 vccd1 _3833_/A sky130_fd_sc_hd__mux2_1
X_6551_ _6551_/A vssd1 vssd1 vccd1 vccd1 _7859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5502_ _5502_/A vssd1 vssd1 vccd1 vccd1 _7889_/D sky130_fd_sc_hd__clkbuf_1
X_8221_ _8335_/CLK _8221_/D vssd1 vssd1 vccd1 vccd1 _8221_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3194_ clkbuf_0__3194_/X vssd1 vssd1 vccd1 vccd1 _6446__230/A sky130_fd_sc_hd__clkbuf_4
X_5433_ _7919_/Q _4523_/X _5437_/S vssd1 vssd1 vccd1 vccd1 _5434_/A sky130_fd_sc_hd__mux2_1
X_5364_ _3840_/X _7952_/Q _5364_/S vssd1 vssd1 vccd1 vccd1 _5365_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8152_ _8152_/CLK _8152_/D vssd1 vssd1 vccd1 vccd1 _8152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7103_ _7432_/A _7216_/A _7216_/B vssd1 vssd1 vccd1 vccd1 _7104_/D sky130_fd_sc_hd__and3_1
X_4315_ _8150_/Q _4134_/X _4315_/S vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5295_ _7988_/Q vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__clkbuf_4
X_8083_ _8083_/CLK _8083_/D vssd1 vssd1 vccd1 vccd1 _8083_/Q sky130_fd_sc_hd__dfxtp_1
X_4246_ _4246_/A vssd1 vssd1 vccd1 vccd1 _8180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _8208_/Q _4090_/X _4177_/S vssd1 vssd1 vccd1 vccd1 _4178_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2978_ clkbuf_0__2978_/X vssd1 vssd1 vccd1 vccd1 _6103__191/A sky130_fd_sc_hd__clkbuf_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088__179 _6089__180/A vssd1 vssd1 vccd1 vccd1 _7648_/CLK sky130_fd_sc_hd__inv_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7936_ _7936_/CLK _7936_/D vssd1 vssd1 vccd1 vccd1 _7936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7867_ _8342_/CLK _7867_/D vssd1 vssd1 vccd1 vccd1 _7867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7798_ _7798_/CLK _7798_/D vssd1 vssd1 vccd1 vccd1 _7798_/Q sky130_fd_sc_hd__dfxtp_1
X_6749_ _7416_/B _7416_/C _7596_/A vssd1 vssd1 vccd1 vccd1 _6749_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7372__7 _7372__7/A vssd1 vssd1 vccd1 vccd1 _8309_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7037__70 _7037__70/A vssd1 vssd1 vccd1 vccd1 _8167_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7349__164 _7349__164/A vssd1 vssd1 vccd1 vccd1 _8291_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4100_ _8265_/Q _4099_/X _4100_/S vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__mux2_1
X_5080_ _8183_/Q _8175_/Q _7897_/Q _7913_/Q _4995_/A _5181_/A vssd1 vssd1 vccd1 vccd1
+ _5080_/X sky130_fd_sc_hd__mux4_2
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4031_ _4031_/A vssd1 vssd1 vccd1 vccd1 _8279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5982_ _7715_/Q input28/X _5991_/S vssd1 vssd1 vccd1 vccd1 _5982_/X sky130_fd_sc_hd__mux2_4
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7721_ _7991_/CLK _7721_/D vssd1 vssd1 vccd1 vccd1 _7721_/Q sky130_fd_sc_hd__dfxtp_1
X_4933_ _4323_/X _8021_/Q _4941_/S vssd1 vssd1 vccd1 vccd1 _4934_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7652_ _7652_/CLK _7652_/D vssd1 vssd1 vccd1 vccd1 _7652_/Q sky130_fd_sc_hd__dfxtp_1
X_4864_ _8050_/Q _4865_/A _4863_/Y _4774_/X vssd1 vssd1 vccd1 vccd1 _8050_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7583_ _7610_/A _7583_/B vssd1 vssd1 vccd1 vccd1 _8390_/D sky130_fd_sc_hd__nor2_1
X_3815_ _6249_/A _3799_/X _3814_/X _6350_/B vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__a31oi_4
X_4795_ _4686_/X _4793_/X _4794_/X vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6534_ _7591_/B _7852_/Q _6534_/S vssd1 vssd1 vccd1 vccd1 _6535_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6465_ _6465_/A vssd1 vssd1 vccd1 vccd1 _6465_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3246_ clkbuf_0__3246_/X vssd1 vssd1 vccd1 vccd1 _6612__320/A sky130_fd_sc_hd__clkbuf_4
X_8204_ _8231_/CLK _8204_/D vssd1 vssd1 vccd1 vccd1 _8204_/Q sky130_fd_sc_hd__dfxtp_1
X_5416_ _5416_/A vssd1 vssd1 vccd1 vccd1 _7927_/D sky130_fd_sc_hd__clkbuf_1
Xoutput142 _5898_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput120 _5926_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__buf_2
Xoutput131 _5876_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__buf_2
X_6396_ _7859_/Q _7752_/Q _6666_/S vssd1 vssd1 vccd1 vccd1 _6397_/A sky130_fd_sc_hd__mux2_1
Xoutput153 _5856_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__buf_2
X_5347_ _4120_/C _5347_/B _5347_/C vssd1 vssd1 vccd1 vccd1 _5421_/B sky130_fd_sc_hd__nand3b_2
X_8135_ _8135_/CLK _8135_/D vssd1 vssd1 vccd1 vccd1 _8135_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput175 _6050_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput186 _5984_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__buf_2
Xoutput164 _6015_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0__3600_ clkbuf_0__3600_/X vssd1 vssd1 vccd1 vccd1 _7385__18/A sky130_fd_sc_hd__clkbuf_4
X_5278_ _5547_/A vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__clkbuf_2
X_8066_ _8066_/CLK _8066_/D vssd1 vssd1 vccd1 vccd1 _8066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4229_ _8365_/Q vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__buf_2
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3393_ clkbuf_0__3393_/X vssd1 vssd1 vccd1 vccd1 _6977__522/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7919_ _7919_/CLK _7919_/D vssd1 vssd1 vccd1 vccd1 _7919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _6062_/A sky130_fd_sc_hd__clkbuf_1
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
X_4580_ _4580_/A vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__clkbuf_4
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__buf_4
Xinput55 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _7608_/B sky130_fd_sc_hd__buf_6
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput88 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _6536_/A sky130_fd_sc_hd__buf_6
Xinput66 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _5880_/A sky130_fd_sc_hd__buf_4
Xinput77 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__buf_4
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6250_ _6350_/C vssd1 vssd1 vccd1 vccd1 _6301_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6181_ _6181_/A vssd1 vssd1 vccd1 vccd1 _7700_/D sky130_fd_sc_hd__clkbuf_1
X_5201_ _7878_/Q _7945_/Q _5274_/A vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5132_ _8369_/Q _5114_/X _5183_/A _8377_/Q _5123_/S vssd1 vssd1 vccd1 vccd1 _5132_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5063_ _5269_/A _5060_/X _5062_/X vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4014_ _3875_/X _8286_/Q _4018_/S vssd1 vssd1 vccd1 vccd1 _4015_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6462__243 _6462__243/A vssd1 vssd1 vccd1 vccd1 _7800_/CLK sky130_fd_sc_hd__inv_2
X_5965_ _5965_/A vssd1 vssd1 vccd1 vccd1 _5965_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7330__149 _7331__150/A vssd1 vssd1 vccd1 vccd1 _8276_/CLK sky130_fd_sc_hd__inv_2
X_5896_ _5896_/A vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__clkbuf_1
X_4916_ _8028_/Q _4392_/X _4922_/S vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7704_ _7704_/CLK _7704_/D vssd1 vssd1 vccd1 vccd1 _7704_/Q sky130_fd_sc_hd__dfxtp_1
X_7635_ _7422_/A _4052_/X _7635_/S vssd1 vssd1 vccd1 vccd1 _7636_/B sky130_fd_sc_hd__mux2_1
X_4847_ _5793_/S vssd1 vssd1 vccd1 vccd1 _5785_/S sky130_fd_sc_hd__buf_4
X_7031__65 _7031__65/A vssd1 vssd1 vccd1 vccd1 _8162_/CLK sky130_fd_sc_hd__inv_2
X_6989__531 _6991__533/A vssd1 vssd1 vccd1 vccd1 _8128_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4778_ _8196_/Q _4681_/X _4715_/X _4777_/X vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7497_ _7402_/B _7510_/A _7490_/Y vssd1 vssd1 vccd1 vccd1 _7497_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6379_ _6379_/A vssd1 vssd1 vccd1 vccd1 _7744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8118_ _8118_/CLK _8118_/D vssd1 vssd1 vccd1 vccd1 _8118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8049_ _8049_/CLK _8049_/D vssd1 vssd1 vccd1 vccd1 _8049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3376_ clkbuf_0__3376_/X vssd1 vssd1 vccd1 vccd1 _6898__462/A sky130_fd_sc_hd__clkbuf_4
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8411__233 vssd1 vssd1 vccd1 vccd1 partID[4] _8411__233/LO sky130_fd_sc_hd__conb_1
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6671__362 _6671__362/A vssd1 vssd1 vccd1 vccd1 _7946_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5750_ _5750_/A vssd1 vssd1 vccd1 vccd1 _7762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _7792_/Q _5587_/X _5681_/S vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__mux2_1
X_4701_ _8048_/Q vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__buf_2
X_7420_ _7596_/A _7420_/B vssd1 vssd1 vccd1 vccd1 _7435_/A sky130_fd_sc_hd__xor2_1
X_4632_ _4632_/A vssd1 vssd1 vccd1 vccd1 _4632_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ _7976_/Q _7968_/Q _7772_/Q _8037_/Q _4872_/A _4562_/X vssd1 vssd1 vccd1 vccd1
+ _4563_/X sky130_fd_sc_hd__mux4_2
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7351_ _7357_/A vssd1 vssd1 vccd1 vccd1 _7351_/X sky130_fd_sc_hd__buf_1
X_4494_ _4494_/A vssd1 vssd1 vccd1 vccd1 _8081_/D sky130_fd_sc_hd__clkbuf_1
X_6302_ _8399_/Q vssd1 vssd1 vccd1 vccd1 _7615_/A sky130_fd_sc_hd__clkbuf_4
X_7282_ _8010_/Q _7266_/A _7281_/X _7178_/X vssd1 vssd1 vccd1 vccd1 _8238_/D sky130_fd_sc_hd__o211a_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6233_ _6341_/A vssd1 vssd1 vccd1 vccd1 _6342_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6164_ _6164_/A _6554_/B vssd1 vssd1 vccd1 vccd1 _6180_/S sky130_fd_sc_hd__nand2_4
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/A vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5046_ _8311_/Q _8303_/Q _8295_/Q _8319_/Q _5149_/S _5010_/X vssd1 vssd1 vccd1 vccd1
+ _5046_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5948_ _5948_/A vssd1 vssd1 vccd1 vccd1 _5948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5888_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7618_ _7618_/A _7618_/B vssd1 vssd1 vccd1 vccd1 _7641_/S sky130_fd_sc_hd__and2_1
XFILLER_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7549_ _7617_/A _7549_/B _7549_/C vssd1 vssd1 vccd1 vccd1 _7550_/A sky130_fd_sc_hd__and3_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6469__249 _6470__250/A vssd1 vssd1 vccd1 vccd1 _7806_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3359_ clkbuf_0__3359_/X vssd1 vssd1 vccd1 vccd1 _6826__409/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6970__516 _6971__517/A vssd1 vssd1 vccd1 vccd1 _8113_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6920_ _6944_/A vssd1 vssd1 vccd1 vccd1 _6920_/X sky130_fd_sc_hd__buf_1
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6851_ _6851_/A vssd1 vssd1 vccd1 vccd1 _6851_/X sky130_fd_sc_hd__buf_1
X_5802_ _5802_/A vssd1 vssd1 vccd1 vccd1 _7650_/D sky130_fd_sc_hd__clkbuf_1
X_6678__368 _6680__370/A vssd1 vssd1 vccd1 vccd1 _7952_/CLK sky130_fd_sc_hd__inv_2
X_3994_ _3994_/A vssd1 vssd1 vccd1 vccd1 _8295_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3600_ _7382_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3600_/X sky130_fd_sc_hd__clkbuf_16
X_5733_ _7769_/Q _5558_/A _5735_/S vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5664_ _5664_/A vssd1 vssd1 vccd1 vccd1 _7800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7403_ _7399_/A input1/X _7447_/B _7400_/X _7506_/A vssd1 vssd1 vccd1 vccd1 _7439_/B
+ sky130_fd_sc_hd__o311a_1
X_4615_ _8089_/Q _8081_/Q _8044_/Q _8113_/Q _4579_/X _4580_/X vssd1 vssd1 vccd1 vccd1
+ _4615_/X sky130_fd_sc_hd__mux4_1
X_8383_ _8383_/CLK _8383_/D vssd1 vssd1 vccd1 vccd1 _8383_/Q sky130_fd_sc_hd__dfxtp_1
X_5595_ _5595_/A vssd1 vssd1 vccd1 vccd1 _7830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4546_ _8049_/Q _4564_/A vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__and2_1
Xclkbuf_0__3393_ _6975_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3393_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4477_ _4477_/A vssd1 vssd1 vccd1 vccd1 _8088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7265_ _7265_/A _7265_/B vssd1 vssd1 vccd1 vccd1 _7266_/A sky130_fd_sc_hd__or2_1
X_6216_ _6320_/A vssd1 vssd1 vccd1 vccd1 _6216_/X sky130_fd_sc_hd__clkbuf_2
X_7196_ _7199_/A _7202_/A vssd1 vssd1 vccd1 vccd1 _7196_/X sky130_fd_sc_hd__or2_1
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6147_ _6145_/X _7857_/Q _6142_/X _6146_/X _7681_/Q vssd1 vssd1 vccd1 vccd1 _7681_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_13 _6054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6118_/A vssd1 vssd1 vccd1 vccd1 _7600_/A sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_35 _5918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_46 _5181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _5029_/A vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6475__253 _6477__255/A vssd1 vssd1 vccd1 vccd1 _7810_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7343__159 _7344__160/A vssd1 vssd1 vccd1 vccd1 _8286_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6935__488 _6936__489/A vssd1 vssd1 vccd1 vccd1 _8085_/CLK sky130_fd_sc_hd__inv_2
X_4400_ _4400_/A vssd1 vssd1 vccd1 vccd1 _8119_/D sky130_fd_sc_hd__clkbuf_1
X_5380_ _5380_/A vssd1 vssd1 vccd1 vccd1 _7946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4331_ _4331_/A vssd1 vssd1 vccd1 vccd1 _8145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4262_ _4220_/X _8173_/Q _4266_/S vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6001_ _6001_/A vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__clkbuf_1
X_4193_ _4193_/A vssd1 vssd1 vccd1 vccd1 _8200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7952_ _7952_/CLK _7952_/D vssd1 vssd1 vccd1 vccd1 _7952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7883_ _7883_/CLK _7883_/D vssd1 vssd1 vccd1 vccd1 _7883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6834_ _6834_/A vssd1 vssd1 vccd1 vccd1 _6834_/X sky130_fd_sc_hd__buf_1
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6765_ _7519_/A _6765_/B _7402_/B vssd1 vssd1 vccd1 vccd1 _6766_/A sky130_fd_sc_hd__and3_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3977_ _3977_/A vssd1 vssd1 vccd1 vccd1 _8302_/D sky130_fd_sc_hd__clkbuf_1
X_5716_ _5716_/A vssd1 vssd1 vccd1 vccd1 _7777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6696_ _8342_/Q _8341_/Q _8340_/Q _8339_/Q vssd1 vssd1 vccd1 vccd1 _6744_/D sky130_fd_sc_hd__and4_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5647_ _7807_/Q _5590_/X _5651_/S vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5578_ _7991_/Q vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__clkbuf_4
X_8366_ _8366_/CLK _8366_/D vssd1 vssd1 vccd1 vccd1 _8366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3376_ _6896_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3376_/X sky130_fd_sc_hd__clkbuf_16
X_4529_ _8358_/Q vssd1 vssd1 vccd1 vccd1 _4529_/X sky130_fd_sc_hd__clkbuf_4
X_8297_ _8297_/CLK _8297_/D vssd1 vssd1 vccd1 vccd1 _8297_/Q sky130_fd_sc_hd__dfxtp_1
X_7248_ _7202_/A _7247_/Y _7222_/A _7233_/A _7151_/A vssd1 vssd1 vccd1 vccd1 _7249_/B
+ sky130_fd_sc_hd__o32a_1
X_7179_ _7262_/B _7174_/C _7178_/X vssd1 vssd1 vccd1 vccd1 _7179_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4880_ _4880_/A vssd1 vssd1 vccd1 vccd1 _8044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3900_ _3900_/A vssd1 vssd1 vccd1 vccd1 _8327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7070__96 _7071__97/A vssd1 vssd1 vccd1 vccd1 _8193_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3400_ clkbuf_0__3400_/X vssd1 vssd1 vccd1 vccd1 _7332_/A sky130_fd_sc_hd__clkbuf_4
X_3831_ _8361_/Q vssd1 vssd1 vccd1 vccd1 _3831_/X sky130_fd_sc_hd__clkbuf_4
X_6550_ _5884_/A _7859_/Q _6552_/S vssd1 vssd1 vccd1 vccd1 _6551_/A sky130_fd_sc_hd__mux2_1
X_5501_ _5292_/X _7889_/Q _5503_/S vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3262_ clkbuf_0__3262_/X vssd1 vssd1 vccd1 vccd1 _6683__372/A sky130_fd_sc_hd__clkbuf_4
X_8220_ _8335_/CLK _8220_/D vssd1 vssd1 vccd1 vccd1 _8220_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3193_ clkbuf_0__3193_/X vssd1 vssd1 vccd1 vccd1 _6465_/A sky130_fd_sc_hd__clkbuf_4
X_5432_ _5432_/A vssd1 vssd1 vccd1 vccd1 _7920_/D sky130_fd_sc_hd__clkbuf_1
X_5363_ _5363_/A vssd1 vssd1 vccd1 vccd1 _7953_/D sky130_fd_sc_hd__clkbuf_1
X_8151_ _8151_/CLK _8151_/D vssd1 vssd1 vccd1 vccd1 _8151_/Q sky130_fd_sc_hd__dfxtp_1
X_6983__526 _6985__528/A vssd1 vssd1 vccd1 vccd1 _8123_/CLK sky130_fd_sc_hd__inv_2
X_7102_ _7216_/A _7216_/B _7432_/A vssd1 vssd1 vccd1 vccd1 _7104_/C sky130_fd_sc_hd__a21oi_1
X_4314_ _4314_/A vssd1 vssd1 vccd1 vccd1 _8151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8082_ _8082_/CLK _8082_/D vssd1 vssd1 vccd1 vccd1 _8082_/Q sky130_fd_sc_hd__dfxtp_1
X_5294_ _5294_/A vssd1 vssd1 vccd1 vccd1 _7981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4245_ _8180_/Q _4140_/X _4247_/S vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__mux2_1
X_4176_ _4176_/A vssd1 vssd1 vccd1 vccd1 _8209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6426__214 _6427__215/A vssd1 vssd1 vccd1 vccd1 _7771_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__2977_ clkbuf_0__2977_/X vssd1 vssd1 vccd1 vccd1 _6101__190/A sky130_fd_sc_hd__clkbuf_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7935_ _7935_/CLK _7935_/D vssd1 vssd1 vccd1 vccd1 _7935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7866_ _8342_/CLK _7866_/D vssd1 vssd1 vccd1 vccd1 _7866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7797_ _7797_/CLK _7797_/D vssd1 vssd1 vccd1 vccd1 _7797_/Q sky130_fd_sc_hd__dfxtp_1
X_6748_ _6748_/A vssd1 vssd1 vccd1 vccd1 _7416_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_117_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8349_ _8349_/CLK _8349_/D vssd1 vssd1 vccd1 vccd1 _8349_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3359_ _6822_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3359_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6778__384 _6779__385/A vssd1 vssd1 vccd1 vccd1 _7969_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4030_ _8279_/Q _3939_/X _4036_/S vssd1 vssd1 vccd1 vccd1 _4031_/A sky130_fd_sc_hd__mux2_1
X_7004__544 _7004__544/A vssd1 vssd1 vccd1 vccd1 _8141_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5981_ _5981_/A vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__clkbuf_1
X_7720_ _8391_/CLK _7720_/D vssd1 vssd1 vccd1 vccd1 _7720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4932_ _4947_/S vssd1 vssd1 vccd1 vccd1 _4941_/S sky130_fd_sc_hd__clkbuf_4
X_7651_ _7651_/CLK _7651_/D vssd1 vssd1 vccd1 vccd1 _7651_/Q sky130_fd_sc_hd__dfxtp_1
X_4863_ _4869_/A _4863_/B vssd1 vssd1 vccd1 vccd1 _4863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7582_ _7579_/Y _7399_/A _7586_/S vssd1 vssd1 vccd1 vccd1 _7583_/B sky130_fd_sc_hd__mux2_1
X_3814_ _3814_/A vssd1 vssd1 vccd1 vccd1 _3814_/X sky130_fd_sc_hd__buf_2
XFILLER_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4794_ _8108_/Q _4724_/X _4725_/X _8084_/Q _4726_/X vssd1 vssd1 vccd1 vccd1 _4794_/X
+ sky130_fd_sc_hd__o221a_1
X_6533_ _6533_/A vssd1 vssd1 vccd1 vccd1 _7851_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3245_ clkbuf_0__3245_/X vssd1 vssd1 vccd1 vccd1 _6602__311/A sky130_fd_sc_hd__clkbuf_4
Xoutput110 _5961_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__buf_2
XFILLER_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8203_ _8231_/CLK _8203_/D vssd1 vssd1 vccd1 vccd1 _8203_/Q sky130_fd_sc_hd__dfxtp_1
X_5415_ _7927_/Q _4523_/X _5419_/S vssd1 vssd1 vccd1 vccd1 _5416_/A sky130_fd_sc_hd__mux2_1
Xoutput143 _5900_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput132 _5878_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput121 _5826_/B vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__buf_2
X_6395_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6666_/S sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8364_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput154 _5825_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _5346_/A vssd1 vssd1 vccd1 vccd1 _7961_/D sky130_fd_sc_hd__clkbuf_1
X_8134_ _8134_/CLK _8134_/D vssd1 vssd1 vccd1 vccd1 _8134_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput165 _6018_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput176 _6054_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _7992_/Q vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__clkbuf_2
X_8065_ _8065_/CLK _8065_/D vssd1 vssd1 vccd1 vccd1 _8065_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput187 _5987_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__buf_2
X_6094__184 _6095__185/A vssd1 vssd1 vccd1 vccd1 _7653_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4228_ _4228_/A vssd1 vssd1 vccd1 vccd1 _8187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3392_ clkbuf_0__3392_/X vssd1 vssd1 vccd1 vccd1 _6974__520/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4159_ _4159_/A vssd1 vssd1 vccd1 vccd1 _8244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _7918_/CLK _7918_/D vssd1 vssd1 vccd1 vccd1 _7918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7849_ _7991_/CLK _7849_/D vssd1 vssd1 vccd1 vccd1 _7849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 _6034_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _6064_/A sky130_fd_sc_hd__clkbuf_1
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__buf_8
XFILLER_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput78 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__buf_4
Xinput89 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _6554_/A sky130_fd_sc_hd__clkbuf_8
Xinput67 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _5882_/A sky130_fd_sc_hd__buf_4
Xinput56 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _7605_/B sky130_fd_sc_hd__buf_6
XFILLER_115_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6180_ _7617_/A _7700_/Q _6180_/S vssd1 vssd1 vccd1 vccd1 _6181_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5200_ _5271_/A _5198_/X _5199_/X _5269_/A vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5131_ _7880_/Q _7947_/Q _5234_/S vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5062_ _4976_/X _5061_/X _5154_/A vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__a21o_1
X_4013_ _4013_/A vssd1 vssd1 vccd1 vccd1 _8287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7016__52 _7016__52/A vssd1 vssd1 vccd1 vccd1 _8149_/CLK sky130_fd_sc_hd__inv_2
X_5964_ _7864_/Q _5964_/B vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__and2_1
X_7703_ _8335_/CLK _7703_/D vssd1 vssd1 vccd1 vccd1 _7703_/Q sky130_fd_sc_hd__dfxtp_1
X_5895_ _5895_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5896_/A sky130_fd_sc_hd__or2_1
X_4915_ _4915_/A vssd1 vssd1 vccd1 vccd1 _8029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7634_ _7634_/A vssd1 vssd1 vccd1 vccd1 _8404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4846_ _5795_/B _5725_/A vssd1 vssd1 vccd1 vccd1 _5793_/S sky130_fd_sc_hd__nor2_4
XFILLER_119_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6206__193 _6208__195/A vssd1 vssd1 vccd1 vccd1 _7705_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _4717_/X _7814_/Q _7798_/Q _4691_/X vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__a22o_1
X_7496_ _7496_/A _7496_/B vssd1 vssd1 vccd1 vccd1 _7510_/A sky130_fd_sc_hd__and2_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6447_ _6453_/A vssd1 vssd1 vccd1 vccd1 _6447_/X sky130_fd_sc_hd__buf_1
X_6378_ _5936_/A _7744_/Q _6382_/S vssd1 vssd1 vccd1 vccd1 _6379_/A sky130_fd_sc_hd__mux2_1
X_7298__123 _7298__123/A vssd1 vssd1 vccd1 vccd1 _8250_/CLK sky130_fd_sc_hd__inv_2
X_8117_ _8117_/CLK _8117_/D vssd1 vssd1 vccd1 vccd1 _8117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5329_ _5761_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _5345_/S sky130_fd_sc_hd__or2_2
XFILLER_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6881__449 _6882__450/A vssd1 vssd1 vccd1 vccd1 _8044_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3513_ clkbuf_0__3513_/X vssd1 vssd1 vccd1 vccd1 _7288__115/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8048_ _8048_/CLK _8048_/D vssd1 vssd1 vccd1 vccd1 _8048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3375_ clkbuf_0__3375_/X vssd1 vssd1 vccd1 vccd1 _6895__460/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5680_ _5680_/A vssd1 vssd1 vccd1 vccd1 _7793_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4700_ _4697_/X _7707_/Q _7656_/Q _4699_/X vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__a22o_1
X_4631_ _4329_/X _4538_/X _4630_/X _4609_/X vssd1 vssd1 vccd1 vccd1 _8063_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4562_ _4580_/A vssd1 vssd1 vccd1 vccd1 _4562_/X sky130_fd_sc_hd__clkbuf_4
X_4493_ _4329_/X _8081_/Q _4499_/S vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__mux2_1
X_6301_ _6332_/C _6301_/B _6312_/A vssd1 vssd1 vccd1 vccd1 _6301_/X sky130_fd_sc_hd__and3_1
X_7281_ _8238_/Q _7283_/B vssd1 vssd1 vccd1 vccd1 _7281_/X sky130_fd_sc_hd__or2_1
X_6232_ _8057_/Q vssd1 vssd1 vccd1 vccd1 _6232_/Y sky130_fd_sc_hd__inv_2
X_6163_ _6350_/B _6188_/B vssd1 vssd1 vccd1 vccd1 _6554_/B sky130_fd_sc_hd__nor2_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A _5045_/B vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__and2_1
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5947_ _7856_/Q _5953_/B vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__and2_1
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5878_ _5878_/A vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__clkbuf_1
X_7617_ _7617_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7617_/Y sky130_fd_sc_hd__nand2_1
X_7185__109 _7186__110/A vssd1 vssd1 vccd1 vccd1 _8208_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4829_ _4703_/A _7757_/Q _4705_/A _8014_/Q _4726_/A vssd1 vssd1 vccd1 vccd1 _4829_/X
+ sky130_fd_sc_hd__o221a_1
X_7548_ _7548_/A vssd1 vssd1 vccd1 vccd1 _8364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7479_ _8341_/Q _7466_/X _7474_/X _7418_/B vssd1 vssd1 vccd1 vccd1 _7480_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8441__216 vssd1 vssd1 vccd1 vccd1 _8441__216/HI manufacturerID[8] sky130_fd_sc_hd__conb_1
XFILLER_29_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3358_ clkbuf_0__3358_/X vssd1 vssd1 vccd1 vccd1 _6820__404/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6818__402 _6820__404/A vssd1 vssd1 vccd1 vccd1 _7995_/CLK sky130_fd_sc_hd__inv_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _4084_/X _7650_/Q _5805_/S vssd1 vssd1 vccd1 vccd1 _5802_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5732_ _5732_/A vssd1 vssd1 vccd1 vccd1 _7770_/D sky130_fd_sc_hd__clkbuf_1
X_3993_ _8295_/Q _3939_/X _3999_/S vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__mux2_1
X_6420__209 _6421__210/A vssd1 vssd1 vccd1 vccd1 _7766_/CLK sky130_fd_sc_hd__inv_2
X_5663_ _5561_/X _7800_/Q _5663_/S vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__mux2_1
X_7402_ _7489_/A _7402_/B vssd1 vssd1 vccd1 vccd1 _7506_/A sky130_fd_sc_hd__or2_1
X_4614_ _4867_/B _4611_/X _4613_/X vssd1 vssd1 vccd1 vccd1 _4614_/X sky130_fd_sc_hd__a21o_1
X_8382_ _8382_/CLK _8382_/D vssd1 vssd1 vccd1 vccd1 _8382_/Q sky130_fd_sc_hd__dfxtp_1
X_5594_ _7830_/Q _5593_/X _5597_/S vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__mux2_1
X_4545_ _8048_/Q _8047_/Q _8046_/Q vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__and3_1
X_7333_ _7339_/A vssd1 vssd1 vccd1 vccd1 _7333_/X sky130_fd_sc_hd__buf_1
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3392_ _6969_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3392_/X sky130_fd_sc_hd__clkbuf_16
X_4476_ _4332_/X _8088_/Q _4480_/S vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__mux2_1
X_7264_ _7178_/X _7254_/B _7263_/Y _7260_/Y _8231_/Q vssd1 vssd1 vccd1 vccd1 _8231_/D
+ sky130_fd_sc_hd__a32o_1
X_6215_ _7546_/C vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7195_ _7220_/A vssd1 vssd1 vccd1 vccd1 _7202_/A sky130_fd_sc_hd__clkbuf_2
X_6146_ _6154_/A vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__clkbuf_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_14 _6054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_36 _5920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6077_ _6144_/A vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_47 _5972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5028_ _4953_/X _5023_/X _5025_/X _5027_/X vssd1 vssd1 vccd1 vccd1 _8011_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6772__379 _6772__379/A vssd1 vssd1 vccd1 vccd1 _7964_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6894__459 _6895__460/A vssd1 vssd1 vccd1 vccd1 _8054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4329_/X _8145_/Q _4339_/S vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__mux2_1
X_4261_ _4261_/A vssd1 vssd1 vccd1 vccd1 _8174_/D sky130_fd_sc_hd__clkbuf_1
X_6000_ _7669_/Q _5999_/X _6006_/S vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__mux2_4
XFILLER_86_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4192_ _8200_/Q _4084_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__mux2_1
X_6684__373 _6686__375/A vssd1 vssd1 vccd1 vccd1 _7957_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6645__346 _6647__348/A vssd1 vssd1 vccd1 vccd1 _7927_/CLK sky130_fd_sc_hd__inv_2
X_7951_ _7951_/CLK _7951_/D vssd1 vssd1 vccd1 vccd1 _7951_/Q sky130_fd_sc_hd__dfxtp_1
X_6902_ _6913_/A vssd1 vssd1 vccd1 vccd1 _6902_/X sky130_fd_sc_hd__buf_1
X_7882_ _7882_/CLK _7882_/D vssd1 vssd1 vccd1 vccd1 _7882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6764_ _8349_/Q _8348_/Q _8347_/Q vssd1 vssd1 vccd1 vccd1 _7402_/B sky130_fd_sc_hd__and3_1
X_3976_ _8302_/Q _3943_/X _3980_/S vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6695_ _6744_/B vssd1 vssd1 vccd1 vccd1 _6738_/B sky130_fd_sc_hd__clkbuf_2
X_5715_ _7777_/Q _5584_/X _5717_/S vssd1 vssd1 vccd1 vccd1 _5716_/A sky130_fd_sc_hd__mux2_1
X_5646_ _5646_/A vssd1 vssd1 vccd1 vccd1 _7808_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3513_ _7187_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3513_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5577_ _5577_/A vssd1 vssd1 vccd1 vccd1 _7836_/D sky130_fd_sc_hd__clkbuf_1
X_8365_ _8365_/CLK _8365_/D vssd1 vssd1 vccd1 vccd1 _8365_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4528_ _4528_/A vssd1 vssd1 vccd1 vccd1 _8068_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3375_ _6890_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3375_/X sky130_fd_sc_hd__clkbuf_16
X_8296_ _8296_/CLK _8296_/D vssd1 vssd1 vccd1 vccd1 _8296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7247_ _7247_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7247_/Y sky130_fd_sc_hd__nand2_1
X_4459_ _4459_/A vssd1 vssd1 vccd1 vccd1 _8096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7178_ _7285_/S vssd1 vssd1 vccd1 vccd1 _7178_/X sky130_fd_sc_hd__clkbuf_2
X_6129_ _6129_/A vssd1 vssd1 vccd1 vccd1 _6129_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8447__222 vssd1 vssd1 vccd1 vccd1 _8447__222/HI partID[7] sky130_fd_sc_hd__conb_1
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6941__493 _6941__493/A vssd1 vssd1 vccd1 vccd1 _8090_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7319__140 _7319__140/A vssd1 vssd1 vccd1 vccd1 _8267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _3830_/A vssd1 vssd1 vccd1 vccd1 _8386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5500_ _5500_/A vssd1 vssd1 vccd1 vccd1 _7890_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3261_ clkbuf_0__3261_/X vssd1 vssd1 vccd1 vccd1 _6680__370/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3192_ clkbuf_0__3192_/X vssd1 vssd1 vccd1 vccd1 _6437__223/A sky130_fd_sc_hd__clkbuf_4
X_5431_ _7920_/Q _4520_/X _5431_/S vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__mux2_1
X_5362_ _3837_/X _7953_/Q _5364_/S vssd1 vssd1 vccd1 vccd1 _5363_/A sky130_fd_sc_hd__mux2_1
X_8150_ _8150_/CLK _8150_/D vssd1 vssd1 vccd1 vccd1 _8150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8081_ _8081_/CLK _8081_/D vssd1 vssd1 vccd1 vccd1 _8081_/Q sky130_fd_sc_hd__dfxtp_1
X_7101_ _8402_/Q vssd1 vssd1 vccd1 vccd1 _7432_/A sky130_fd_sc_hd__inv_2
X_4313_ _8151_/Q _4131_/X _4315_/S vssd1 vssd1 vccd1 vccd1 _4314_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5293_ _5292_/X _7981_/Q _5297_/S vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__mux2_1
X_7032_ _7038_/A vssd1 vssd1 vccd1 vccd1 _7032_/X sky130_fd_sc_hd__buf_1
XFILLER_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4244_ _4244_/A vssd1 vssd1 vccd1 vccd1 _8181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4175_ _8209_/Q _4087_/X _4177_/S vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__mux2_1
X_7292__118 _7294__120/A vssd1 vssd1 vccd1 vccd1 _8245_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__2976_ clkbuf_0__2976_/X vssd1 vssd1 vccd1 vccd1 _6093__183/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7934_ _7934_/CLK _7934_/D vssd1 vssd1 vccd1 vccd1 _7934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7865_ _8342_/CLK _7865_/D vssd1 vssd1 vccd1 vccd1 _7865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7796_ _7796_/CLK _7796_/D vssd1 vssd1 vccd1 vccd1 _7796_/Q sky130_fd_sc_hd__dfxtp_1
X_6816_ _6834_/A vssd1 vssd1 vccd1 vccd1 _6816_/X sky130_fd_sc_hd__buf_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6747_ _8393_/Q _7416_/B _6748_/A vssd1 vssd1 vccd1 vccd1 _6747_/X sky130_fd_sc_hd__and3_1
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _4223_/A vssd1 vssd1 vccd1 vccd1 _3959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5629_ _5564_/X _7815_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__mux2_1
X_8348_ _8348_/CLK _8348_/D vssd1 vssd1 vccd1 vccd1 _8348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3358_ _6816_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3358_/X sky130_fd_sc_hd__clkbuf_16
X_8279_ _8279_/CLK _8279_/D vssd1 vssd1 vccd1 vccd1 _8279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6488__264 _6489__265/A vssd1 vssd1 vccd1 vccd1 _7821_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5980_ _7663_/Q _5979_/X _5989_/S vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4931_ _5795_/A _5743_/B vssd1 vssd1 vccd1 vccd1 _4947_/S sky130_fd_sc_hd__or2_2
X_7650_ _7650_/CLK _7650_/D vssd1 vssd1 vccd1 vccd1 _7650_/Q sky130_fd_sc_hd__dfxtp_1
X_4862_ _4872_/B vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7043__75 _7043__75/A vssd1 vssd1 vccd1 vccd1 _8172_/CLK sky130_fd_sc_hd__inv_2
X_3813_ _6236_/A _6285_/A _6241_/D vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__a21boi_2
X_6601_ _6601_/A vssd1 vssd1 vccd1 vccd1 _6601_/X sky130_fd_sc_hd__buf_1
X_7581_ _7943_/Q _7618_/B vssd1 vssd1 vccd1 vccd1 _7586_/S sky130_fd_sc_hd__nand2_1
X_4793_ _8076_/Q _4716_/X _4687_/X _8039_/Q vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6532_ _7595_/B _7851_/Q _6534_/S vssd1 vssd1 vccd1 vccd1 _6533_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3244_ clkbuf_0__3244_/X vssd1 vssd1 vccd1 vccd1 _6600__310/A sky130_fd_sc_hd__clkbuf_4
Xoutput100 _5941_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__buf_2
X_8202_ _8202_/CLK _8202_/D vssd1 vssd1 vccd1 vccd1 _8202_/Q sky130_fd_sc_hd__dfxtp_1
X_5414_ _5414_/A vssd1 vssd1 vccd1 vccd1 _7928_/D sky130_fd_sc_hd__clkbuf_1
Xoutput111 _5963_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput133 _5839_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput122 _5837_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__buf_2
X_6394_ _6394_/A vssd1 vssd1 vccd1 vccd1 _7751_/D sky130_fd_sc_hd__clkbuf_1
X_8133_ _8133_/CLK _8133_/D vssd1 vssd1 vccd1 vccd1 _8133_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput144 _5841_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput155 _5827_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5345_ _5308_/X _7961_/Q _5345_/S vssd1 vssd1 vccd1 vccd1 _5346_/A sky130_fd_sc_hd__mux2_1
X_6948__499 _6949__500/A vssd1 vssd1 vccd1 vccd1 _8096_/CLK sky130_fd_sc_hd__inv_2
Xoutput166 _6021_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput177 _6056_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8064_ _8064_/CLK _8064_/D vssd1 vssd1 vccd1 vccd1 _8064_/Q sky130_fd_sc_hd__dfxtp_1
X_5276_ _5276_/A vssd1 vssd1 vccd1 vccd1 _7993_/D sky130_fd_sc_hd__clkbuf_1
X_6844__420 _6844__420/A vssd1 vssd1 vccd1 vccd1 _8015_/CLK sky130_fd_sc_hd__inv_2
Xoutput188 _5990_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__buf_2
X_7300__125 _7300__125/A vssd1 vssd1 vccd1 vccd1 _8252_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4227_ _4226_/X _8187_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7077__101 _7081__105/A vssd1 vssd1 vccd1 vccd1 _8198_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3391_ clkbuf_0__3391_/X vssd1 vssd1 vccd1 vccd1 _6966__513/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _8244_/Q _4090_/X _4158_/S vssd1 vssd1 vccd1 vccd1 _4159_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4089_ _4089_/A vssd1 vssd1 vccd1 vccd1 _8269_/D sky130_fd_sc_hd__clkbuf_1
X_6582__296 _6586__300/A vssd1 vssd1 vccd1 vccd1 _7877_/CLK sky130_fd_sc_hd__inv_2
X_7917_ _7917_/CLK _7917_/D vssd1 vssd1 vccd1 vccd1 _7917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7848_ _7992_/CLK _7848_/D vssd1 vssd1 vccd1 vccd1 _7848_/Q sky130_fd_sc_hd__dfxtp_1
X_6658__356 _6668__360/A vssd1 vssd1 vccd1 vccd1 _7937_/CLK sky130_fd_sc_hd__inv_2
X_7779_ _7779_/CLK _7779_/D vssd1 vssd1 vccd1 vccd1 _7779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3589_ clkbuf_0__3589_/X vssd1 vssd1 vccd1 vccd1 _7331__150/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6602__311 _6602__311/A vssd1 vssd1 vccd1 vccd1 _7892_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 _6042_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _6066_/A sky130_fd_sc_hd__clkbuf_1
Xinput35 caravel_wb_error_i vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__clkbuf_1
Xinput46 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__buf_8
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput57 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__buf_6
Xinput79 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _7538_/B sky130_fd_sc_hd__buf_8
Xinput68 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__buf_4
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A vssd1 vssd1 vccd1 vccd1 _5218_/A sky130_fd_sc_hd__clkbuf_2
X_5061_ _8184_/Q _8176_/Q _7898_/Q _7914_/Q _4995_/A _5207_/S vssd1 vssd1 vccd1 vccd1
+ _5061_/X sky130_fd_sc_hd__mux4_2
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4012_ _3872_/X _8287_/Q _4018_/S vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5963_ _5963_/A vssd1 vssd1 vccd1 vccd1 _5963_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7702_ _7747_/CLK _7702_/D vssd1 vssd1 vccd1 vccd1 _7702_/Q sky130_fd_sc_hd__dfxtp_1
X_4914_ _8029_/Q _4386_/X _4922_/S vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__mux2_1
X_5894_ _5894_/A vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7633_ _6145_/X _7633_/B vssd1 vssd1 vccd1 vccd1 _7634_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4845_ _5617_/B vssd1 vssd1 vccd1 vccd1 _5725_/A sky130_fd_sc_hd__clkbuf_4
X_4776_ _7782_/Q _4573_/B _4676_/X vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6515_ _6575_/A vssd1 vssd1 vccd1 vccd1 _6515_/X sky130_fd_sc_hd__buf_1
X_7495_ _8347_/Q vssd1 vssd1 vccd1 vccd1 _7498_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6377_ _6377_/A vssd1 vssd1 vccd1 vccd1 _7743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8116_ _8116_/CLK _8116_/D vssd1 vssd1 vccd1 vccd1 _8116_/Q sky130_fd_sc_hd__dfxtp_1
X_5328_ _5328_/A vssd1 vssd1 vccd1 vccd1 _7969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8047_ _8047_/CLK _8047_/D vssd1 vssd1 vccd1 vccd1 _8047_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0_0__3512_ clkbuf_0__3512_/X vssd1 vssd1 vccd1 vccd1 _7184__108/A sky130_fd_sc_hd__clkbuf_4
X_5259_ _3894_/B _5259_/B _7547_/A vssd1 vssd1 vccd1 vccd1 _5260_/A sky130_fd_sc_hd__and3b_1
XFILLER_57_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3374_ clkbuf_0__3374_/X vssd1 vssd1 vccd1 vccd1 _6888__454/A sky130_fd_sc_hd__clkbuf_4
X_6996__537 _6998__539/A vssd1 vssd1 vccd1 vccd1 _8134_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6439__225 _6439__225/A vssd1 vssd1 vccd1 vccd1 _7782_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4630_ _4540_/X _8063_/Q _4869_/A _4629_/X _4605_/X vssd1 vssd1 vccd1 vccd1 _4630_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6300_ _7942_/Q vssd1 vssd1 vccd1 vccd1 _6332_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4561_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4492_ _4492_/A vssd1 vssd1 vccd1 vccd1 _8082_/D sky130_fd_sc_hd__clkbuf_1
X_7280_ _8009_/Q _7266_/A _7279_/X _7178_/X vssd1 vssd1 vccd1 vccd1 _8237_/D sky130_fd_sc_hd__o211a_1
X_6231_ _6231_/A vssd1 vssd1 vccd1 vccd1 _6231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6162_ _7868_/Q _6157_/X _6116_/A _6129_/A _7692_/Q vssd1 vssd1 vccd1 vccd1 _7692_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6609__317 _6611__319/A vssd1 vssd1 vccd1 vccd1 _7898_/CLK sky130_fd_sc_hd__inv_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _8388_/Q _8327_/Q _8073_/Q _8105_/Q _5042_/X _5234_/S vssd1 vssd1 vccd1 vccd1
+ _5045_/B sky130_fd_sc_hd__mux4_1
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5946_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5877_ _5877_/A _5877_/B vssd1 vssd1 vccd1 vccd1 _5878_/A sky130_fd_sc_hd__or2_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7616_ _7599_/B _7614_/Y _7615_/Y _7600_/X vssd1 vssd1 vccd1 vccd1 _8399_/D sky130_fd_sc_hd__a211oi_2
X_4828_ _4716_/A _7869_/Q _7773_/Q _4717_/A vssd1 vssd1 vccd1 vccd1 _4828_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7547_ _7547_/A _7547_/B _7547_/C vssd1 vssd1 vccd1 vccd1 _7548_/A sky130_fd_sc_hd__and3_1
X_4759_ _8267_/Q _4719_/Y _4720_/X _8243_/Q _4556_/A vssd1 vssd1 vccd1 vccd1 _4759_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7478_ _7482_/A _7478_/B vssd1 vssd1 vccd1 vccd1 _8340_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_12_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8065_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3357_ clkbuf_0__3357_/X vssd1 vssd1 vccd1 vccd1 _6845_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7313__135 _7313__135/A vssd1 vssd1 vccd1 vccd1 _8262_/CLK sky130_fd_sc_hd__inv_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _5800_/A vssd1 vssd1 vccd1 vccd1 _7651_/D sky130_fd_sc_hd__clkbuf_1
X_6780_ _6786_/A vssd1 vssd1 vccd1 vccd1 _6780_/X sky130_fd_sc_hd__buf_1
X_3992_ _3992_/A vssd1 vssd1 vccd1 vccd1 _8296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _7770_/Q _5555_/A _5735_/S vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5662_ _5662_/A vssd1 vssd1 vccd1 vccd1 _7801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7401_ _8330_/Q _7401_/B vssd1 vssd1 vccd1 vccd1 _7489_/A sky130_fd_sc_hd__nand2_2
X_4613_ _4567_/X _4612_/X _4575_/X vssd1 vssd1 vccd1 vccd1 _4613_/X sky130_fd_sc_hd__a21o_1
X_8381_ _8381_/CLK _8381_/D vssd1 vssd1 vccd1 vccd1 _8381_/Q sky130_fd_sc_hd__dfxtp_1
X_5593_ _7986_/Q vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__clkbuf_2
X_4544_ _4872_/B vssd1 vssd1 vccd1 vccd1 _4869_/A sky130_fd_sc_hd__buf_2
Xclkbuf_0__3391_ _6963_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3391_/X sky130_fd_sc_hd__clkbuf_16
X_7332_ _7332_/A vssd1 vssd1 vccd1 vccd1 _7332_/X sky130_fd_sc_hd__buf_1
XFILLER_116_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7263_ _7263_/A vssd1 vssd1 vccd1 vccd1 _7263_/Y sky130_fd_sc_hd__inv_2
X_4475_ _4475_/A vssd1 vssd1 vccd1 vccd1 _8089_/D sky130_fd_sc_hd__clkbuf_1
X_6214_ _6214_/A vssd1 vssd1 vccd1 vccd1 _7546_/C sky130_fd_sc_hd__clkbuf_2
X_7194_ _7237_/B vssd1 vssd1 vccd1 vccd1 _7194_/X sky130_fd_sc_hd__clkbuf_2
X_6145_ _6281_/A vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__buf_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_15 _6056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6076_ _6350_/B vssd1 vssd1 vccd1 vccd1 _6144_/A sky130_fd_sc_hd__clkbuf_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_26 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_48 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_37 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5027_ _7533_/A vssd1 vssd1 vccd1 vccd1 _5027_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7386__19 _7387__20/A vssd1 vssd1 vccd1 vccd1 _8321_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5929_ _5929_/A _5931_/B vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__and2_1
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3589_ _7326_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3589_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6482__259 _6482__259/A vssd1 vssd1 vccd1 vccd1 _7816_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3409_ clkbuf_0__3409_/X vssd1 vssd1 vccd1 vccd1 _7056__85/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4260_ _4217_/X _8174_/Q _4260_/S vssd1 vssd1 vccd1 vccd1 _4261_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4191_/A vssd1 vssd1 vccd1 vccd1 _8201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7950_ _7950_/CLK _7950_/D vssd1 vssd1 vccd1 vccd1 _7950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7881_ _7881_/CLK _7881_/D vssd1 vssd1 vccd1 vccd1 _7881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6953__502 _6955__504/A vssd1 vssd1 vccd1 vccd1 _8099_/CLK sky130_fd_sc_hd__inv_2
X_6763_ _6763_/A _6763_/B _7410_/B _7496_/A vssd1 vssd1 vccd1 vccd1 _6765_/B sky130_fd_sc_hd__and4_1
X_3975_ _3975_/A vssd1 vssd1 vccd1 vccd1 _8303_/D sky130_fd_sc_hd__clkbuf_1
X_6694_ _8341_/Q _6702_/A _6702_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _6694_/X sky130_fd_sc_hd__and4_1
X_5714_ _5714_/A vssd1 vssd1 vccd1 vccd1 _7778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5645_ _7808_/Q _5587_/X _5645_/S vssd1 vssd1 vccd1 vccd1 _5646_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3512_ _7181_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3512_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5576_ _7836_/Q _5573_/X _5588_/S vssd1 vssd1 vccd1 vccd1 _5577_/A sky130_fd_sc_hd__mux2_1
X_8364_ _8364_/CLK _8364_/D vssd1 vssd1 vccd1 vccd1 _8364_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_0__3374_ _6884_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3374_/X sky130_fd_sc_hd__clkbuf_16
X_4527_ _8068_/Q _4526_/X _4530_/S vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__mux2_1
X_8295_ _8295_/CLK _8295_/D vssd1 vssd1 vccd1 vccd1 _8295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7246_ _7251_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _8226_/D sky130_fd_sc_hd__nor2_1
X_4458_ _3825_/X _8096_/Q _4462_/S vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7177_ _7177_/A vssd1 vssd1 vccd1 vccd1 _7262_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6128_ _6157_/A vssd1 vssd1 vccd1 vccd1 _6128_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4389_ _4411_/S vssd1 vssd1 vccd1 vccd1 _4402_/S sky130_fd_sc_hd__buf_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__and2_1
XFILLER_105_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7055__84 _7055__84/A vssd1 vssd1 vccd1 vccd1 _8181_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3260_ clkbuf_0__3260_/X vssd1 vssd1 vccd1 vccd1 _6671__362/A sky130_fd_sc_hd__clkbuf_4
X_5430_ _5430_/A vssd1 vssd1 vccd1 vccd1 _7921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3191_ clkbuf_0__3191_/X vssd1 vssd1 vccd1 vccd1 _6433__220/A sky130_fd_sc_hd__clkbuf_4
X_5361_ _5361_/A vssd1 vssd1 vccd1 vccd1 _7954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _5558_/A vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__buf_2
X_8080_ _8080_/CLK _8080_/D vssd1 vssd1 vccd1 vccd1 _8080_/Q sky130_fd_sc_hd__dfxtp_1
X_7100_ _7129_/A _7119_/A _7110_/C vssd1 vssd1 vccd1 vccd1 _7216_/B sky130_fd_sc_hd__a21o_1
X_4312_ _4312_/A vssd1 vssd1 vccd1 vccd1 _8152_/D sky130_fd_sc_hd__clkbuf_1
X_4243_ _8181_/Q _4137_/X _4247_/S vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4174_ _4174_/A vssd1 vssd1 vccd1 vccd1 _8210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2975_ clkbuf_0__2975_/X vssd1 vssd1 vccd1 vccd1 _6089__180/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7933_ _7933_/CLK _7933_/D vssd1 vssd1 vccd1 vccd1 _7933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7864_ _8345_/CLK _7864_/D vssd1 vssd1 vccd1 vccd1 _7864_/Q sky130_fd_sc_hd__dfxtp_1
X_7795_ _7795_/CLK _7795_/D vssd1 vssd1 vccd1 vccd1 _7795_/Q sky130_fd_sc_hd__dfxtp_1
X_6815_ _6815_/A vssd1 vssd1 vccd1 vccd1 _6815_/X sky130_fd_sc_hd__buf_1
X_6746_ _8345_/Q _8344_/Q _6757_/D vssd1 vssd1 vccd1 vccd1 _6748_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3958_ _8359_/Q vssd1 vssd1 vccd1 vccd1 _4223_/A sky130_fd_sc_hd__buf_2
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3889_ _3889_/A vssd1 vssd1 vccd1 vccd1 _8367_/D sky130_fd_sc_hd__clkbuf_1
X_5628_ _5628_/A vssd1 vssd1 vccd1 vccd1 _7816_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3389_ clkbuf_0__3389_/X vssd1 vssd1 vccd1 vccd1 _6955__504/A sky130_fd_sc_hd__clkbuf_4
X_8347_ _8349_/CLK _8347_/D vssd1 vssd1 vccd1 vccd1 _8347_/Q sky130_fd_sc_hd__dfxtp_1
X_5559_ _5558_/X _7841_/Q _5562_/S vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3357_ _6815_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3357_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8278_ _8278_/CLK _8278_/D vssd1 vssd1 vccd1 vccd1 _8278_/Q sky130_fd_sc_hd__dfxtp_1
X_7229_ _7244_/A _7229_/B vssd1 vssd1 vccd1 vccd1 _8220_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6594__305 _6594__305/A vssd1 vssd1 vccd1 vccd1 _7886_/CLK sky130_fd_sc_hd__inv_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7028__62 _7029__63/A vssd1 vssd1 vccd1 vccd1 _8159_/CLK sky130_fd_sc_hd__inv_2
X_4930_ _4930_/A _4930_/B _4930_/C vssd1 vssd1 vccd1 vccd1 _5743_/B sky130_fd_sc_hd__nand3_4
XFILLER_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4861_ _4324_/A _4853_/B _4860_/Y vssd1 vssd1 vccd1 vccd1 _8051_/D sky130_fd_sc_hd__a21oi_1
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3812_ _3812_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6241_/D sky130_fd_sc_hd__nor2_1
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7580_ _6350_/C _6226_/C _6285_/A _7540_/B _6226_/B vssd1 vssd1 vccd1 vccd1 _7618_/B
+ sky130_fd_sc_hd__a2111oi_4
X_4792_ _4715_/X _4790_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _4792_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6531_ _6531_/A vssd1 vssd1 vccd1 vccd1 _7850_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3243_ clkbuf_0__3243_/X vssd1 vssd1 vccd1 vccd1 _6592__303/A sky130_fd_sc_hd__clkbuf_4
Xoutput101 _5943_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__buf_2
X_6393_ _7858_/Q _7751_/Q _6393_/S vssd1 vssd1 vccd1 vccd1 _6394_/A sky130_fd_sc_hd__mux2_1
X_8201_ _8201_/CLK _8201_/D vssd1 vssd1 vccd1 vccd1 _8201_/Q sky130_fd_sc_hd__dfxtp_1
X_5413_ _7928_/Q _4520_/X _5413_/S vssd1 vssd1 vccd1 vccd1 _5414_/A sky130_fd_sc_hd__mux2_1
Xoutput112 _5965_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput134 _5881_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput123 _5859_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__buf_2
X_5344_ _5344_/A vssd1 vssd1 vccd1 vccd1 _7962_/D sky130_fd_sc_hd__clkbuf_1
X_8132_ _8132_/CLK _8132_/D vssd1 vssd1 vccd1 vccd1 _8132_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput145 _5902_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__buf_2
Xoutput156 _5831_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__buf_2
Xoutput167 _6024_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8063_ _8063_/CLK _8063_/D vssd1 vssd1 vccd1 vccd1 _8063_/Q sky130_fd_sc_hd__dfxtp_1
X_5275_ _7533_/A _5275_/B _5275_/C vssd1 vssd1 vccd1 vccd1 _5276_/A sky130_fd_sc_hd__and3_1
Xoutput189 _5994_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__buf_2
Xoutput178 _6058_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__buf_2
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7014_ _7026_/A vssd1 vssd1 vccd1 vccd1 _7014_/X sky130_fd_sc_hd__buf_1
X_4226_ _4226_/A vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4157_ _4157_/A vssd1 vssd1 vccd1 vccd1 _8245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3390_ clkbuf_0__3390_/X vssd1 vssd1 vccd1 vccd1 _6962__510/A sky130_fd_sc_hd__clkbuf_4
X_4088_ _8269_/Q _4087_/X _4091_/S vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7916_ _7916_/CLK _7916_/D vssd1 vssd1 vccd1 vccd1 _7916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7847_ _7992_/CLK _7847_/D vssd1 vssd1 vccd1 vccd1 _7847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7778_ _7778_/CLK _7778_/D vssd1 vssd1 vccd1 vccd1 _7778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6729_ _7423_/B _7423_/C _7422_/A vssd1 vssd1 vccd1 vccd1 _6729_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3409_ _7051_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3409_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3588_ clkbuf_0__3588_/X vssd1 vssd1 vccd1 vccd1 _7322__142/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_2
Xinput36 wb_rst_i vssd1 vssd1 vccd1 vccd1 _6350_/B sky130_fd_sc_hd__clkbuf_16
Xinput47 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__buf_6
Xinput58 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _7598_/B sky130_fd_sc_hd__clkbuf_8
Xinput69 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _5886_/A sky130_fd_sc_hd__buf_4
X_7362__175 _7362__175/A vssd1 vssd1 vccd1 vccd1 _8302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5060_ _7938_/Q _7930_/Q _7922_/Q _7957_/Q _4978_/X _4995_/X vssd1 vssd1 vccd1 vccd1
+ _5060_/X sky130_fd_sc_hd__mux4_1
X_4011_ _4011_/A vssd1 vssd1 vccd1 vccd1 _8288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _7863_/Q _5964_/B vssd1 vssd1 vccd1 vccd1 _5963_/A sky130_fd_sc_hd__and2_1
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7701_ _8397_/CLK _7701_/D vssd1 vssd1 vccd1 vccd1 _7701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ _4928_/S vssd1 vssd1 vccd1 vccd1 _4922_/S sky130_fd_sc_hd__buf_4
X_5893_ _5893_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5894_/A sky130_fd_sc_hd__or2_1
X_7632_ _7135_/A _3799_/X _7635_/S vssd1 vssd1 vccd1 vccd1 _7633_/B sky130_fd_sc_hd__mux2_1
X_4844_ _4844_/A _4854_/B vssd1 vssd1 vccd1 vccd1 _5617_/B sky130_fd_sc_hd__nand2_4
XFILLER_21_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4775_ _4341_/X _4538_/A _4773_/X _4774_/X vssd1 vssd1 vccd1 vccd1 _8059_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494_ _7494_/A vssd1 vssd1 vccd1 vccd1 _8346_/D sky130_fd_sc_hd__clkbuf_1
X_6376_ _5934_/A _7743_/Q _6382_/S vssd1 vssd1 vccd1 vccd1 _6377_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8115_ _8115_/CLK _8115_/D vssd1 vssd1 vccd1 vccd1 _8115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5327_ _5308_/X _7969_/Q _5327_/S vssd1 vssd1 vccd1 vccd1 _5328_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8046_ _8046_/CLK _8046_/D vssd1 vssd1 vccd1 vccd1 _8046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _5261_/A _5261_/B _3867_/A vssd1 vssd1 vccd1 vccd1 _5259_/B sky130_fd_sc_hd__a21o_1
X_5189_ _5271_/A _5186_/X _5188_/X vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__o21a_1
X_4209_ _4208_/X _8193_/Q _4218_/S vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6213__199 _6213__199/A vssd1 vssd1 vccd1 vccd1 _7711_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3373_ clkbuf_0__3373_/X vssd1 vssd1 vccd1 vccd1 _6896_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7558__33 _7559__34/A vssd1 vssd1 vccd1 vccd1 _8372_/CLK sky130_fd_sc_hd__inv_2
X_7022__57 _7022__57/A vssd1 vssd1 vccd1 vccd1 _8154_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4682_/A vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4491_ _4323_/X _8082_/Q _4499_/S vssd1 vssd1 vccd1 vccd1 _4492_/A sky130_fd_sc_hd__mux2_1
X_6230_ _6230_/A vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6161_ _7867_/Q _6157_/X _6116_/A _6129_/A _7691_/Q vssd1 vssd1 vccd1 vccd1 _7691_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _8292_/Q _8300_/Q _5181_/A vssd1 vssd1 vccd1 vccd1 _5112_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5234_/S sky130_fd_sc_hd__buf_2
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _7000_/A vssd1 vssd1 vccd1 vccd1 _6994_/X sky130_fd_sc_hd__buf_1
X_5945_ _7855_/Q _5953_/B vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__and2_1
X_5876_ _5876_/A vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7615_ _7615_/A _7615_/B vssd1 vssd1 vccd1 vccd1 _7615_/Y sky130_fd_sc_hd__nor2_1
X_4827_ _8030_/Q _4683_/A _4720_/X _7969_/Q _4826_/X vssd1 vssd1 vccd1 vccd1 _4827_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7546_ _7546_/A _7546_/B _7546_/C vssd1 vssd1 vccd1 vccd1 _7547_/C sky130_fd_sc_hd__and3_1
X_4758_ _8141_/Q _4716_/X _4717_/X _7823_/Q vssd1 vssd1 vccd1 vccd1 _4758_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7477_ _6700_/Y _7447_/B _7461_/X _6704_/B vssd1 vssd1 vccd1 vccd1 _7478_/B sky130_fd_sc_hd__o22a_1
X_4689_ _4730_/A vssd1 vssd1 vccd1 vccd1 _4696_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6428_ _6434_/A vssd1 vssd1 vccd1 vccd1 _6428_/X sky130_fd_sc_hd__buf_1
XFILLER_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _6359_/A vssd1 vssd1 vccd1 vccd1 _7735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8029_ _8029_/CLK _8029_/D vssd1 vssd1 vccd1 vccd1 _8029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6864__435 _6864__435/A vssd1 vssd1 vccd1 vccd1 _8030_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6825__408 _6827__410/A vssd1 vssd1 vccd1 vccd1 _8001_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3991_ _8296_/Q _3966_/X _3999_/S vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _5730_/A vssd1 vssd1 vccd1 vccd1 _7771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7400_ _8330_/Q _7450_/B _7529_/A vssd1 vssd1 vccd1 vccd1 _7400_/X sky130_fd_sc_hd__or3_1
X_5661_ _5558_/X _7801_/Q _5663_/S vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__mux2_1
X_4612_ _8020_/Q _7875_/Q _7779_/Q _7763_/Q _4569_/X _4571_/X vssd1 vssd1 vccd1 vccd1
+ _4612_/X sky130_fd_sc_hd__mux4_1
X_7552__28 _7553__29/A vssd1 vssd1 vccd1 vccd1 _8367_/CLK sky130_fd_sc_hd__inv_2
X_5592_ _5592_/A vssd1 vssd1 vccd1 vccd1 _7831_/D sky130_fd_sc_hd__clkbuf_1
X_8380_ _8380_/CLK _8380_/D vssd1 vssd1 vccd1 vccd1 _8380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4543_ _4632_/A vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__3390_ _6957_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3390_/X sky130_fd_sc_hd__clkbuf_16
X_6615__322 _6615__322/A vssd1 vssd1 vccd1 vccd1 _7903_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7262_ _8231_/Q _7262_/B _7262_/C _7262_/D vssd1 vssd1 vccd1 vccd1 _7263_/A sky130_fd_sc_hd__or4_1
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4474_ _4329_/X _8089_/Q _4480_/S vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__mux2_1
X_7193_ _7177_/A _7174_/C _7192_/Y vssd1 vssd1 vccd1 vccd1 _7237_/B sky130_fd_sc_hd__o21a_1
X_6144_ _6144_/A vssd1 vssd1 vccd1 vccd1 _6281_/A sky130_fd_sc_hd__buf_2
XFILLER_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6075_ _7540_/A _7756_/Q _6072_/X _6074_/X vssd1 vssd1 vccd1 vccd1 _6075_/X sky130_fd_sc_hd__a22o_4
XFILLER_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_16 _6056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _6838_/A vssd1 vssd1 vccd1 vccd1 _7533_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_49 _5909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_38 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_27 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5928_ _5928_/A vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5859_ _5859_/A vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7529_ _7529_/A _7529_/B vssd1 vssd1 vccd1 vccd1 _7529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3588_ _7320_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3588_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6516__286 _6517__287/A vssd1 vssd1 vccd1 vccd1 _7843_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3408_ clkbuf_0__3408_/X vssd1 vssd1 vccd1 vccd1 _7050__80/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4190_ _8201_/Q _4081_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4191_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7880_ _7880_/CLK _7880_/D vssd1 vssd1 vccd1 vccd1 _7880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6762_ _7450_/A _7401_/B vssd1 vssd1 vccd1 vccd1 _7496_/A sky130_fd_sc_hd__and2_1
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _8303_/Q _3939_/X _3980_/S vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__mux2_1
X_6693_ _6744_/C vssd1 vssd1 vccd1 vccd1 _6702_/C sky130_fd_sc_hd__clkbuf_2
X_5713_ _7778_/Q _5581_/X _5717_/S vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__mux2_1
X_5644_ _5644_/A vssd1 vssd1 vccd1 vccd1 _7809_/D sky130_fd_sc_hd__clkbuf_1
X_7391__23 _7393__25/A vssd1 vssd1 vccd1 vccd1 _8325_/CLK sky130_fd_sc_hd__inv_2
X_8431__206 vssd1 vssd1 vccd1 vccd1 _8431__206/HI core1Index[6] sky130_fd_sc_hd__conb_1
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8363_ _8365_/CLK _8363_/D vssd1 vssd1 vccd1 vccd1 _8363_/Q sky130_fd_sc_hd__dfxtp_4
X_5575_ _5597_/S vssd1 vssd1 vccd1 vccd1 _5588_/S sky130_fd_sc_hd__clkbuf_4
X_7314_ _7326_/A vssd1 vssd1 vccd1 vccd1 _7314_/X sky130_fd_sc_hd__buf_1
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3373_ _6883_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3373_/X sky130_fd_sc_hd__clkbuf_16
X_4526_ _8359_/Q vssd1 vssd1 vccd1 vccd1 _4526_/X sky130_fd_sc_hd__clkbuf_2
X_8294_ _8294_/CLK _8294_/D vssd1 vssd1 vccd1 vccd1 _8294_/Q sky130_fd_sc_hd__dfxtp_1
X_7245_ _7202_/A _7164_/B _7222_/A _7233_/A _7151_/B vssd1 vssd1 vccd1 vccd1 _7246_/B
+ sky130_fd_sc_hd__o32a_1
X_4457_ _4457_/A vssd1 vssd1 vccd1 vccd1 _8097_/D sky130_fd_sc_hd__clkbuf_1
X_7176_ _8204_/Q vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__inv_2
X_6127_ _6119_/X _7846_/Q _6126_/X _6120_/X _7670_/Q vssd1 vssd1 vccd1 vccd1 _7670_/D
+ sky130_fd_sc_hd__o32a_1
X_4388_ _4912_/A _5671_/B vssd1 vssd1 vccd1 vccd1 _4411_/S sky130_fd_sc_hd__nor2_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _7686_/Q _6048_/X _6051_/X _6057_/X vssd1 vssd1 vccd1 vccd1 _6058_/X sky130_fd_sc_hd__o22a_4
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3190_ clkbuf_0__3190_/X vssd1 vssd1 vccd1 vccd1 _6427__215/A sky130_fd_sc_hd__clkbuf_4
X_6458__240 _6458__240/A vssd1 vssd1 vccd1 vccd1 _7797_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5360_ _3834_/X _7954_/Q _5364_/S vssd1 vssd1 vccd1 vccd1 _5361_/A sky130_fd_sc_hd__mux2_1
X_5291_ _7989_/Q vssd1 vssd1 vccd1 vccd1 _5558_/A sky130_fd_sc_hd__clkbuf_4
X_4311_ _8152_/Q _4128_/X _4315_/S vssd1 vssd1 vccd1 vccd1 _4312_/A sky130_fd_sc_hd__mux2_1
X_4242_ _4242_/A vssd1 vssd1 vccd1 vccd1 _8182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _8210_/Q _4084_/X _4177_/S vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2974_ clkbuf_0__2974_/X vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__clkbuf_4
X_7932_ _7932_/CLK _7932_/D vssd1 vssd1 vccd1 vccd1 _7932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7863_ _8345_/CLK _7863_/D vssd1 vssd1 vccd1 vccd1 _7863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7794_ _7794_/CLK _7794_/D vssd1 vssd1 vccd1 vccd1 _7794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6745_ _8344_/Q _6757_/D _8345_/Q vssd1 vssd1 vccd1 vccd1 _7416_/B sky130_fd_sc_hd__a21o_1
X_6918__475 _6918__475/A vssd1 vssd1 vccd1 vccd1 _8072_/CLK sky130_fd_sc_hd__inv_2
X_3957_ _3957_/A vssd1 vssd1 vccd1 vccd1 _8307_/D sky130_fd_sc_hd__clkbuf_1
X_3888_ _3887_/X _8367_/Q _3891_/S vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3388_ clkbuf_0__3388_/X vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__clkbuf_4
X_5627_ _5561_/X _7816_/Q _5627_/S vssd1 vssd1 vccd1 vccd1 _5628_/A sky130_fd_sc_hd__mux2_1
X_8346_ _8349_/CLK _8346_/D vssd1 vssd1 vccd1 vccd1 _8346_/Q sky130_fd_sc_hd__dfxtp_1
X_5558_ _5558_/A vssd1 vssd1 vccd1 vccd1 _5558_/X sky130_fd_sc_hd__buf_2
XFILLER_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4509_ _8074_/Q _4229_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__mux2_1
X_8277_ _8277_/CLK _8277_/D vssd1 vssd1 vccd1 vccd1 _8277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7228_ _7220_/X _7226_/Y _7222_/X _7223_/X _7227_/Y vssd1 vssd1 vccd1 vccd1 _7229_/B
+ sky130_fd_sc_hd__o32a_1
X_5489_ _7894_/Q _4223_/A _5491_/S vssd1 vssd1 vccd1 vccd1 _5490_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7159_ _7159_/A _7159_/B vssd1 vssd1 vccd1 vccd1 _7226_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6628__332 _6628__332/A vssd1 vssd1 vccd1 vccd1 _7913_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_7_wb_clk_i _7717_/CLK vssd1 vssd1 vccd1 vccd1 _7991_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4324_/A _4853_/B _4836_/X vssd1 vssd1 vccd1 vccd1 _4860_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3811_ _6341_/A _6341_/B _6341_/C _6341_/D vssd1 vssd1 vccd1 vccd1 _6226_/B sky130_fd_sc_hd__or4_4
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6530_ _7598_/B _7850_/Q _6534_/S vssd1 vssd1 vccd1 vccd1 _6531_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4791_ _8266_/Q _4719_/Y _4720_/X _8242_/Q _4556_/A vssd1 vssd1 vccd1 vccd1 _4791_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3396_ clkbuf_0__3396_/X vssd1 vssd1 vccd1 vccd1 _6991__533/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1_0__3242_ clkbuf_0__3242_/X vssd1 vssd1 vccd1 vccd1 _6613_/A sky130_fd_sc_hd__clkbuf_4
X_6392_ _6392_/A vssd1 vssd1 vccd1 vccd1 _7750_/D sky130_fd_sc_hd__clkbuf_1
X_8200_ _8200_/CLK _8200_/D vssd1 vssd1 vccd1 vccd1 _8200_/Q sky130_fd_sc_hd__dfxtp_1
X_5412_ _5412_/A vssd1 vssd1 vccd1 vccd1 _7929_/D sky130_fd_sc_hd__clkbuf_1
Xoutput102 _5946_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput124 _5861_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput113 _5910_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__buf_2
X_5343_ _5304_/X _7962_/Q _5345_/S vssd1 vssd1 vccd1 vccd1 _5344_/A sky130_fd_sc_hd__mux2_1
X_8131_ _8131_/CLK _8131_/D vssd1 vssd1 vccd1 vccd1 _8131_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput146 _5904_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput135 _5883_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput157 _5833_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__buf_2
Xoutput168 _6028_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8062_ _8062_/CLK _8062_/D vssd1 vssd1 vccd1 vccd1 _8062_/Q sky130_fd_sc_hd__dfxtp_1
X_5274_ _5274_/A _5274_/B vssd1 vssd1 vccd1 vccd1 _5275_/C sky130_fd_sc_hd__nand2_1
Xoutput179 _6060_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7013_ _7075_/A vssd1 vssd1 vccd1 vccd1 _7013_/X sky130_fd_sc_hd__buf_1
X_4225_ _4225_/A vssd1 vssd1 vccd1 vccd1 _8188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _8245_/Q _4087_/X _4158_/S vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _7989_/Q vssd1 vssd1 vccd1 vccd1 _4087_/X sky130_fd_sc_hd__buf_2
XFILLER_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7915_ _7915_/CLK _7915_/D vssd1 vssd1 vccd1 vccd1 _7915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7846_ _7846_/CLK _7846_/D vssd1 vssd1 vccd1 vccd1 _7846_/Q sky130_fd_sc_hd__dfxtp_1
X_8437__212 vssd1 vssd1 vccd1 vccd1 _8437__212/HI manufacturerID[4] sky130_fd_sc_hd__conb_1
X_7777_ _7777_/CLK _7777_/D vssd1 vssd1 vccd1 vccd1 _7777_/Q sky130_fd_sc_hd__dfxtp_1
X_4989_ _8381_/Q _7951_/Q _7884_/Q _8373_/Q _5198_/S _4971_/X vssd1 vssd1 vccd1 vccd1
+ _4989_/X sky130_fd_sc_hd__mux4_1
X_6728_ _6728_/A vssd1 vssd1 vccd1 vccd1 _7423_/B sky130_fd_sc_hd__clkbuf_2
X_6966__513 _6966__513/A vssd1 vssd1 vccd1 vccd1 _8110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8329_ _8399_/CLK _8329_/D vssd1 vssd1 vccd1 vccd1 _8329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3408_ _7045_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3408_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3587_ clkbuf_0__3587_/X vssd1 vssd1 vccd1 vccd1 _7319__140/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _6068_/A sky130_fd_sc_hd__clkbuf_1
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 _6044_/A sky130_fd_sc_hd__clkbuf_1
X_6791__395 _6791__395/A vssd1 vssd1 vccd1 vccd1 _7980_/CLK sky130_fd_sc_hd__inv_2
Xinput37 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__buf_4
Xinput48 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__buf_6
Xinput59 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _7595_/B sky130_fd_sc_hd__buf_4
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4010_ _3865_/X _8288_/Q _4018_/S vssd1 vssd1 vccd1 vccd1 _4011_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _5961_/A vssd1 vssd1 vccd1 vccd1 _5961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7700_ _7846_/CLK _7700_/D vssd1 vssd1 vccd1 vccd1 _7700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4912_ _4912_/A _5548_/A vssd1 vssd1 vccd1 vccd1 _4928_/S sky130_fd_sc_hd__nor2_2
X_5892_ _5892_/A vssd1 vssd1 vccd1 vccd1 _5892_/X sky130_fd_sc_hd__clkbuf_1
X_7631_ _7629_/Y _7627_/B _7630_/Y _6151_/X vssd1 vssd1 vccd1 vccd1 _8403_/D sky130_fd_sc_hd__a211oi_1
X_4843_ _4843_/A _4843_/B _4843_/C vssd1 vssd1 vccd1 vccd1 _4854_/B sky130_fd_sc_hd__and3_1
XFILLER_20_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _6910_/A vssd1 vssd1 vccd1 vccd1 _4774_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7493_ _7493_/A _7493_/B vssd1 vssd1 vccd1 vccd1 _7494_/A sky130_fd_sc_hd__and2_1
XFILLER_106_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6375_ _6375_/A vssd1 vssd1 vccd1 vccd1 _7742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8114_ _8114_/CLK _8114_/D vssd1 vssd1 vccd1 vccd1 _8114_/Q sky130_fd_sc_hd__dfxtp_1
X_5326_ _5326_/A vssd1 vssd1 vccd1 vccd1 _7970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8045_ _8045_/CLK _8045_/D vssd1 vssd1 vccd1 vccd1 _8045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5257_ _4230_/C _3894_/B _5256_/Y vssd1 vssd1 vccd1 vccd1 _8000_/D sky130_fd_sc_hd__a21oi_1
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _4208_/X sky130_fd_sc_hd__buf_2
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188_ _8156_/Q _5187_/X _5183_/X _8148_/Q _4976_/X vssd1 vssd1 vccd1 vccd1 _5188_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0_0__3372_ clkbuf_0__3372_/X vssd1 vssd1 vccd1 vccd1 _6879__447/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _4139_/A vssd1 vssd1 vccd1 vccd1 _8251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7829_ _7829_/CLK _7829_/D vssd1 vssd1 vccd1 vccd1 _7829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _4505_/S vssd1 vssd1 vccd1 vccd1 _4499_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_109_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6160_ _7866_/Q _6157_/X _6116_/A _6154_/X _7690_/Q vssd1 vssd1 vccd1 vccd1 _7690_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5130_/A vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__buf_2
XFILLER_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5100_/A vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5944_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__clkbuf_2
X_5875_ _5875_/A _5877_/B vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__or2_1
X_7614_ _7614_/A _7614_/B vssd1 vssd1 vccd1 vccd1 _7614_/Y sky130_fd_sc_hd__nand2_1
X_4826_ _4716_/A _7961_/Q _7765_/Q _4731_/X _4729_/A vssd1 vssd1 vccd1 vccd1 _4826_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7545_ _7545_/A vssd1 vssd1 vccd1 vccd1 _8363_/D sky130_fd_sc_hd__clkbuf_1
X_4757_ _4757_/A _4757_/B _4757_/C vssd1 vssd1 vccd1 vccd1 _4757_/X sky130_fd_sc_hd__or3_1
XFILLER_119_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7476_ _7482_/A _7476_/B vssd1 vssd1 vccd1 vccd1 _8339_/D sky130_fd_sc_hd__nor2_1
X_4688_ _8047_/Q vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3208_ clkbuf_0__3208_/X vssd1 vssd1 vccd1 vccd1 _6517__287/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6358_ _5916_/A _7735_/Q _6360_/S vssd1 vssd1 vccd1 vccd1 _6359_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5309_ _5308_/X _7977_/Q _5309_/S vssd1 vssd1 vccd1 vccd1 _5310_/A sky130_fd_sc_hd__mux2_1
X_6289_ _6289_/A _6289_/B vssd1 vssd1 vccd1 vccd1 _6289_/X sky130_fd_sc_hd__and2_1
X_8028_ _8028_/CLK _8028_/D vssd1 vssd1 vccd1 vccd1 _8028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8342_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6452__235 _6452__235/A vssd1 vssd1 vccd1 vccd1 _7792_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3990_ _4005_/S vssd1 vssd1 vccd1 vccd1 _3999_/S sky130_fd_sc_hd__buf_2
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _5660_/A vssd1 vssd1 vccd1 vccd1 _7802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _7975_/Q _7967_/Q _7771_/Q _8036_/Q _4872_/A _4562_/X vssd1 vssd1 vccd1 vccd1
+ _4611_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5591_ _7831_/Q _5590_/X _5597_/S vssd1 vssd1 vccd1 vccd1 _5592_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4542_ _8066_/Q _6230_/A vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__and2_1
X_4473_ _4473_/A vssd1 vssd1 vccd1 vccd1 _8090_/D sky130_fd_sc_hd__clkbuf_1
X_7261_ _8230_/Q _7254_/X _7260_/Y vssd1 vssd1 vccd1 vccd1 _8230_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7192_ _7399_/A _7220_/A vssd1 vssd1 vccd1 vccd1 _7192_/Y sky130_fd_sc_hd__nand2_2
X_6143_ _6136_/X _7856_/Q _6142_/X _6137_/X _7680_/Q vssd1 vssd1 vccd1 vccd1 _7680_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _7731_/Q _6049_/B _7614_/A vssd1 vssd1 vccd1 vccd1 _6074_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_17 _5905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5025_ _5025_/A _5029_/A vssd1 vssd1 vccd1 vccd1 _5025_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_28 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_39 _7538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6622__327 _6622__327/A vssd1 vssd1 vccd1 vccd1 _7908_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5927_ _5927_/A _5931_/B vssd1 vssd1 vccd1 vccd1 _5928_/A sky130_fd_sc_hd__and2_1
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5858_ _7608_/B _5866_/B vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__or2_1
X_4809_ _4697_/X _7704_/Q _7653_/Q _4699_/X vssd1 vssd1 vccd1 vccd1 _4809_/X sky130_fd_sc_hd__a22o_1
X_5789_ _7655_/Q _5564_/A _5793_/S vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__mux2_1
X_7528_ _8356_/Q _7529_/B _7527_/X _7519_/X vssd1 vssd1 vccd1 vccd1 _8356_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_0__3587_ _7314_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3587_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459_ _7423_/B _7423_/C _7446_/Y _7458_/X _8333_/Q vssd1 vssd1 vccd1 vccd1 _7460_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_119_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7067__94 _7068__95/A vssd1 vssd1 vccd1 vccd1 _8191_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3407_ clkbuf_0__3407_/X vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6870__440 _6870__440/A vssd1 vssd1 vccd1 vccd1 _8035_/CLK sky130_fd_sc_hd__inv_2
X_6831__413 _6833__415/A vssd1 vssd1 vccd1 vccd1 _8006_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6761_ _8329_/Q vssd1 vssd1 vccd1 vccd1 _7401_/B sky130_fd_sc_hd__clkinv_2
XFILLER_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _5712_/A vssd1 vssd1 vccd1 vccd1 _7779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _3973_/A vssd1 vssd1 vccd1 vccd1 _8304_/D sky130_fd_sc_hd__clkbuf_1
X_6692_ _8338_/Q _8337_/Q _8336_/Q _8335_/Q vssd1 vssd1 vccd1 vccd1 _6744_/C sky130_fd_sc_hd__and4_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5643_ _7809_/Q _5584_/X _5645_/S vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__mux2_1
X_8362_ _8365_/CLK _8362_/D vssd1 vssd1 vccd1 vccd1 _8362_/Q sky130_fd_sc_hd__dfxtp_4
X_5574_ _5671_/B _5725_/A vssd1 vssd1 vccd1 vccd1 _5597_/S sky130_fd_sc_hd__nor2_2
X_4525_ _4525_/A vssd1 vssd1 vccd1 vccd1 _8069_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3372_ _6877_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3372_/X sky130_fd_sc_hd__clkbuf_16
X_8293_ _8293_/CLK _8293_/D vssd1 vssd1 vccd1 vccd1 _8293_/Q sky130_fd_sc_hd__dfxtp_1
X_7244_ _7244_/A _7244_/B vssd1 vssd1 vccd1 vccd1 _8225_/D sky130_fd_sc_hd__nor2_1
X_4456_ _3822_/X _8097_/Q _4462_/S vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__mux2_1
X_7175_ _7175_/A vssd1 vssd1 vccd1 vccd1 _8203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4387_ _4414_/A _4387_/B _4413_/A vssd1 vssd1 vccd1 vccd1 _5671_/B sky130_fd_sc_hd__or3_4
X_6960__508 _6961__509/A vssd1 vssd1 vccd1 vccd1 _8105_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6126_ _6188_/A vssd1 vssd1 vccd1 vccd1 _6126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _6057_/X sky130_fd_sc_hd__and2_1
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5008_/A vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8454__229 vssd1 vssd1 vccd1 vccd1 _8454__229/HI versionID[3] sky130_fd_sc_hd__conb_1
XFILLER_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _5290_/A vssd1 vssd1 vccd1 vccd1 _7982_/D sky130_fd_sc_hd__clkbuf_1
X_4310_ _4310_/A vssd1 vssd1 vccd1 vccd1 _8153_/D sky130_fd_sc_hd__clkbuf_1
X_4241_ _8182_/Q _4134_/X _4241_/S vssd1 vssd1 vccd1 vccd1 _4242_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ _4172_/A vssd1 vssd1 vccd1 vccd1 _8211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7931_ _7931_/CLK _7931_/D vssd1 vssd1 vccd1 vccd1 _7931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _8345_/CLK _7862_/D vssd1 vssd1 vccd1 vccd1 _7862_/Q sky130_fd_sc_hd__dfxtp_1
X_7793_ _7793_/CLK _7793_/D vssd1 vssd1 vccd1 vccd1 _7793_/Q sky130_fd_sc_hd__dfxtp_1
X_6813_ _6813_/A vssd1 vssd1 vccd1 vccd1 _7992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7061__89 _7061__89/A vssd1 vssd1 vccd1 vccd1 _8186_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6744_ _8343_/Q _6744_/B _6744_/C _6744_/D vssd1 vssd1 vccd1 vccd1 _6757_/D sky130_fd_sc_hd__and4_2
XFILLER_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _8307_/Q _3955_/X _3964_/S vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__mux2_1
X_6675_ _6675_/A vssd1 vssd1 vccd1 vccd1 _6675_/X sky130_fd_sc_hd__buf_1
X_5626_ _5626_/A vssd1 vssd1 vccd1 vccd1 _7817_/D sky130_fd_sc_hd__clkbuf_1
X_3887_ _8359_/Q vssd1 vssd1 vccd1 vccd1 _3887_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8345_ _8345_/CLK _8345_/D vssd1 vssd1 vccd1 vccd1 _8345_/Q sky130_fd_sc_hd__dfxtp_1
X_5557_ _5557_/A vssd1 vssd1 vccd1 vccd1 _7842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5488_ _5488_/A vssd1 vssd1 vccd1 vccd1 _7895_/D sky130_fd_sc_hd__clkbuf_1
X_4508_ _4530_/S vssd1 vssd1 vccd1 vccd1 _4521_/S sky130_fd_sc_hd__clkbuf_4
X_8276_ _8276_/CLK _8276_/D vssd1 vssd1 vccd1 vccd1 _8276_/Q sky130_fd_sc_hd__dfxtp_1
X_7227_ _8220_/Q vssd1 vssd1 vccd1 vccd1 _7227_/Y sky130_fd_sc_hd__inv_2
X_4439_ _4439_/A vssd1 vssd1 vccd1 vccd1 _8105_/D sky130_fd_sc_hd__clkbuf_1
X_7158_ _8400_/Q vssd1 vssd1 vccd1 vccd1 _7430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6109_ _6144_/A _6188_/B vssd1 vssd1 vccd1 vccd1 _6154_/A sky130_fd_sc_hd__or2_2
X_7089_ _8215_/Q vssd1 vssd1 vccd1 vccd1 _7208_/A sky130_fd_sc_hd__clkbuf_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3037_ clkbuf_0__3037_/X vssd1 vssd1 vccd1 vccd1 _6408__200/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3810_ _7743_/Q _7744_/Q _7745_/Q _7742_/Q vssd1 vssd1 vccd1 vccd1 _6341_/D sky130_fd_sc_hd__or4b_1
X_4790_ _8140_/Q _4716_/X _4717_/X _7822_/Q vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__3395_ clkbuf_0__3395_/X vssd1 vssd1 vccd1 vccd1 _6987__530/A sky130_fd_sc_hd__clkbuf_16
X_6391_ _7857_/Q _7750_/Q _6393_/S vssd1 vssd1 vccd1 vccd1 _6392_/A sky130_fd_sc_hd__mux2_1
X_5411_ _7929_/Q _4517_/X _5413_/S vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__mux2_1
Xoutput103 _5948_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__buf_2
Xoutput114 _5913_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput125 _5863_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__buf_2
X_5342_ _5342_/A vssd1 vssd1 vccd1 vccd1 _7963_/D sky130_fd_sc_hd__clkbuf_1
X_8130_ _8130_/CLK _8130_/D vssd1 vssd1 vccd1 vccd1 _8130_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput158 _5821_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput136 _5885_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput147 _5843_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8061_ _8061_/CLK _8061_/D vssd1 vssd1 vccd1 vccd1 _8061_/Q sky130_fd_sc_hd__dfxtp_1
X_5273_ _5274_/A _5274_/B vssd1 vssd1 vccd1 vccd1 _5275_/B sky130_fd_sc_hd__or2_1
Xoutput169 _6031_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__buf_2
X_7012_ _7012_/A vssd1 vssd1 vccd1 vccd1 _7012_/X sky130_fd_sc_hd__buf_1
XFILLER_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4224_ _4223_/X _8188_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__mux2_1
X_4155_ _4155_/A vssd1 vssd1 vccd1 vccd1 _8246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _4086_/A vssd1 vssd1 vccd1 vccd1 _8270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7914_ _7914_/CLK _7914_/D vssd1 vssd1 vccd1 vccd1 _7914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7845_ _7846_/CLK _7845_/D vssd1 vssd1 vccd1 vccd1 _7845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7034__67 _7035__68/A vssd1 vssd1 vccd1 vccd1 _8164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7776_ _7776_/CLK _7776_/D vssd1 vssd1 vccd1 vccd1 _7776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4988_ _5089_/S vssd1 vssd1 vccd1 vccd1 _4988_/X sky130_fd_sc_hd__buf_2
X_6727_ _8405_/Q _6728_/A _7423_/C vssd1 vssd1 vccd1 vccd1 _6727_/X sky130_fd_sc_hd__and3_1
X_3939_ _4208_/A vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__clkbuf_2
X_7309__131 _7311__133/A vssd1 vssd1 vccd1 vccd1 _8258_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5609_ _5561_/X _7824_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5610_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8328_ _8328_/CLK _8328_/D vssd1 vssd1 vccd1 vccd1 _8328_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3407_ _7044_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3407_/X sky130_fd_sc_hd__clkbuf_16
X_6589_ _6601_/A vssd1 vssd1 vccd1 vccd1 _6589_/X sky130_fd_sc_hd__buf_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3724_ clkbuf_0__3724_/X vssd1 vssd1 vccd1 vccd1 _7578__50/A sky130_fd_sc_hd__clkbuf_4
X_8259_ _8259_/CLK _8259_/D vssd1 vssd1 vccd1 vccd1 _8259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3586_ clkbuf_0__3586_/X vssd1 vssd1 vccd1 vccd1 _7313__135/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__clkbuf_1
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _6046_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__buf_6
Xinput38 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5960_ _7862_/Q _5964_/B vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__and2_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _5891_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__or2_1
X_4911_ _4911_/A vssd1 vssd1 vccd1 vccd1 _8030_/D sky130_fd_sc_hd__clkbuf_1
X_7630_ _8403_/Q _7635_/S vssd1 vssd1 vccd1 vccd1 _7630_/Y sky130_fd_sc_hd__nor2_1
X_4842_ _4930_/A _4930_/B _4930_/C vssd1 vssd1 vccd1 vccd1 _5795_/B sky130_fd_sc_hd__nand3b_4
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _4540_/A _8059_/Q _4632_/X _4772_/X _4605_/A vssd1 vssd1 vccd1 vccd1 _4773_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7561_ _7561_/A vssd1 vssd1 vccd1 vccd1 _7561_/X sky130_fd_sc_hd__buf_1
X_7492_ _8346_/Q _7466_/A _7490_/Y _7491_/Y vssd1 vssd1 vccd1 vccd1 _7493_/B sky130_fd_sc_hd__a22o_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6374_ _5931_/A _7742_/Q _6382_/S vssd1 vssd1 vccd1 vccd1 _6375_/A sky130_fd_sc_hd__mux2_1
X_8113_ _8113_/CLK _8113_/D vssd1 vssd1 vccd1 vccd1 _8113_/Q sky130_fd_sc_hd__dfxtp_1
X_5325_ _5304_/X _7970_/Q _5327_/S vssd1 vssd1 vccd1 vccd1 _5326_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8044_ _8044_/CLK _8044_/D vssd1 vssd1 vccd1 vccd1 _8044_/Q sky130_fd_sc_hd__dfxtp_1
X_5256_ _4230_/C _3894_/B _5214_/X vssd1 vssd1 vccd1 vccd1 _5256_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4207_ _4207_/A vssd1 vssd1 vccd1 vccd1 _8194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5187_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0__3371_ clkbuf_0__3371_/X vssd1 vssd1 vccd1 vccd1 _6876__445/A sky130_fd_sc_hd__clkbuf_4
X_4138_ _8251_/Q _4137_/X _4144_/S vssd1 vssd1 vccd1 vccd1 _4139_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4069_ _4069_/A _4069_/B vssd1 vssd1 vccd1 vccd1 _4536_/D sky130_fd_sc_hd__and2_1
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7828_ _7828_/CLK _7828_/D vssd1 vssd1 vccd1 vccd1 _7828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7759_ _7759_/CLK _7759_/D vssd1 vssd1 vccd1 vccd1 _7759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7564__38 _7564__38/A vssd1 vssd1 vccd1 vccd1 _8377_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6090_ _6096_/A vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__buf_1
X_5110_ _5148_/A vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5269_/A _5036_/X _5040_/X vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5943_ _5943_/A vssd1 vssd1 vccd1 vccd1 _5943_/X sky130_fd_sc_hd__clkbuf_1
X_5874_ _5874_/A vssd1 vssd1 vccd1 vccd1 _5874_/X sky130_fd_sc_hd__clkbuf_1
X_7613_ _7599_/B _7611_/Y _7612_/Y _7600_/X vssd1 vssd1 vccd1 vccd1 _8398_/D sky130_fd_sc_hd__a211oi_1
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4825_ _4686_/X _4823_/X _4824_/X vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__o21a_1
X_7544_ _7626_/A _7629_/B _7549_/C vssd1 vssd1 vccd1 vccd1 _7545_/A sky130_fd_sc_hd__and3_1
X_4756_ _8117_/Q _4705_/X _4593_/S _4755_/X vssd1 vssd1 vccd1 vccd1 _4757_/C sky130_fd_sc_hd__o211a_1
X_7475_ _8339_/Q _7466_/X _7474_/X _7412_/B vssd1 vssd1 vccd1 vccd1 _7476_/B sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_1_1_0__3207_ clkbuf_0__3207_/X vssd1 vssd1 vccd1 vccd1 _6514__285/A sky130_fd_sc_hd__clkbuf_4
X_4687_ _4717_/A vssd1 vssd1 vccd1 vccd1 _4687_/X sky130_fd_sc_hd__buf_2
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6357_ _6357_/A vssd1 vssd1 vccd1 vccd1 _7734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5308_ _5570_/A vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__clkbuf_2
X_6288_ _8063_/Q _6231_/X _6287_/X _6244_/X vssd1 vssd1 vccd1 vccd1 _6288_/X sky130_fd_sc_hd__a31o_1
X_8027_ _8027_/CLK _8027_/D vssd1 vssd1 vccd1 vccd1 _8027_/Q sky130_fd_sc_hd__dfxtp_1
X_5239_ _7933_/Q _5151_/X _5017_/A _5238_/X vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__o211a_1
XFILLER_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3037_ _6209_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3037_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_17_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937__490 _6937__490/A vssd1 vssd1 vccd1 vccd1 _8087_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6979__524 _6980__525/A vssd1 vssd1 vccd1 vccd1 _8121_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8422__197 vssd1 vssd1 vccd1 vccd1 _8422__197/HI core0Index[4] sky130_fd_sc_hd__conb_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7288__115 _7288__115/A vssd1 vssd1 vccd1 vccd1 _8242_/CLK sky130_fd_sc_hd__inv_2
X_4610_ _4323_/X _4538_/X _4606_/X _4609_/X vssd1 vssd1 vccd1 vccd1 _8064_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5590_ _7987_/Q vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__clkbuf_2
X_4541_ _4604_/B _4604_/C vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__nand2_1
X_4472_ _4323_/X _8090_/Q _4480_/S vssd1 vssd1 vccd1 vccd1 _4473_/A sky130_fd_sc_hd__mux2_1
X_7260_ _7254_/B _7259_/X _7219_/A vssd1 vssd1 vccd1 vccd1 _7260_/Y sky130_fd_sc_hd__a21oi_1
X_7191_ _8390_/Q vssd1 vssd1 vccd1 vccd1 _7399_/A sky130_fd_sc_hd__clkinv_2
X_6142_ _6188_/A vssd1 vssd1 vccd1 vccd1 _6142_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _7546_/A vssd1 vssd1 vccd1 vccd1 _7614_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_18 _5905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5024_ _8012_/Q _7265_/A vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__nand2_1
XINSDIODE2_29 _5907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6429__216 _6432__219/A vssd1 vssd1 vccd1 vccd1 _7773_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6975_ _6975_/A vssd1 vssd1 vccd1 vccd1 _6975_/X sky130_fd_sc_hd__buf_1
XFILLER_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5926_ _5926_/A vssd1 vssd1 vccd1 vccd1 _5926_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3724_ _7573_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3724_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _5903_/B vssd1 vssd1 vccd1 vccd1 _5866_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5788_ _5788_/A vssd1 vssd1 vccd1 vccd1 _7656_/D sky130_fd_sc_hd__clkbuf_1
X_4808_ _7781_/Q _4683_/A _4681_/X _8195_/Q _4664_/A vssd1 vssd1 vccd1 vccd1 _4808_/X
+ sky130_fd_sc_hd__o221a_1
X_7527_ _8357_/Q _7527_/B _7513_/A vssd1 vssd1 vccd1 vccd1 _7527_/X sky130_fd_sc_hd__or3b_1
X_4739_ _4757_/A _4722_/X _4728_/X _4738_/X _4549_/X vssd1 vssd1 vccd1 vccd1 _4739_/X
+ sky130_fd_sc_hd__o311a_1
Xclkbuf_0__3586_ _7308_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3586_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7458_ _7466_/A vssd1 vssd1 vccd1 vccd1 _7458_/X sky130_fd_sc_hd__buf_2
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6409_ _6502_/A vssd1 vssd1 vccd1 vccd1 _6409_/X sky130_fd_sc_hd__buf_1
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3406_ clkbuf_0__3406_/X vssd1 vssd1 vccd1 vccd1 _7041__73/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3199_ clkbuf_0__3199_/X vssd1 vssd1 vccd1 vccd1 _6478_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7365__1 _7366__2/A vssd1 vssd1 vccd1 vccd1 _8303_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7007__546 _7011__550/A vssd1 vssd1 vccd1 vccd1 _8143_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ _8330_/Q vssd1 vssd1 vccd1 vccd1 _7450_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5711_ _7779_/Q _5578_/X _5717_/S vssd1 vssd1 vccd1 vccd1 _5712_/A sky130_fd_sc_hd__mux2_1
X_3972_ _8304_/Q _3966_/X _3980_/S vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__mux2_1
X_6691_ _6744_/B vssd1 vssd1 vccd1 vccd1 _6702_/B sky130_fd_sc_hd__clkbuf_2
X_5642_ _5642_/A vssd1 vssd1 vccd1 vccd1 _7810_/D sky130_fd_sc_hd__clkbuf_1
X_6578__293 _6580__295/A vssd1 vssd1 vccd1 vccd1 _7874_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5573_ _7992_/Q vssd1 vssd1 vccd1 vccd1 _5573_/X sky130_fd_sc_hd__clkbuf_4
X_8361_ _8365_/CLK _8361_/D vssd1 vssd1 vccd1 vccd1 _8361_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_0__3371_ _6871_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3371_/X sky130_fd_sc_hd__clkbuf_16
X_4524_ _8069_/Q _4523_/X _4530_/S vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__mux2_1
X_8292_ _8292_/CLK _8292_/D vssd1 vssd1 vccd1 vccd1 _8292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7243_ _7220_/X _7167_/B _7222_/X _7223_/X _7242_/Y vssd1 vssd1 vccd1 vccd1 _7244_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4455_ _4455_/A vssd1 vssd1 vccd1 vccd1 _8098_/D sky130_fd_sc_hd__clkbuf_1
X_7303__126 _7306__129/A vssd1 vssd1 vccd1 vccd1 _8253_/CLK sky130_fd_sc_hd__inv_2
X_6097__186 _6098__187/A vssd1 vssd1 vccd1 vccd1 _7655_/CLK sky130_fd_sc_hd__inv_2
X_4386_ _7992_/Q vssd1 vssd1 vccd1 vccd1 _4386_/X sky130_fd_sc_hd__buf_2
X_7174_ _7285_/S _7174_/B _7174_/C vssd1 vssd1 vccd1 vccd1 _7175_/A sky130_fd_sc_hd__and3_1
X_6125_ _6125_/A vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__buf_2
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _7685_/Q _6048_/X _6051_/X _6055_/X vssd1 vssd1 vccd1 vccd1 _6056_/X sky130_fd_sc_hd__o22a_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _5045_/A _5007_/B vssd1 vssd1 vccd1 vccd1 _5007_/X sky130_fd_sc_hd__and2_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5909_ _5909_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__and2_1
XFILLER_10_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7358__171 _7359__172/A vssd1 vssd1 vccd1 vccd1 _8298_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _4240_/A vssd1 vssd1 vccd1 vccd1 _8183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4171_ _8211_/Q _4081_/X _4177_/S vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2972_ clkbuf_0__2972_/X vssd1 vssd1 vccd1 vccd1 _7394_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7930_ _7930_/CLK _7930_/D vssd1 vssd1 vccd1 vccd1 _7930_/Q sky130_fd_sc_hd__dfxtp_1
X_7861_ _8345_/CLK _7861_/D vssd1 vssd1 vccd1 vccd1 _7861_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7046__76 _7048__78/A vssd1 vssd1 vccd1 vccd1 _8173_/CLK sky130_fd_sc_hd__inv_2
X_6812_ _8357_/Q _6907_/C vssd1 vssd1 vccd1 vccd1 _6813_/A sky130_fd_sc_hd__and2_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7792_ _7792_/CLK _7792_/D vssd1 vssd1 vccd1 vccd1 _7792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6743_ _7410_/A _6743_/B _7409_/A _6743_/D vssd1 vssd1 vccd1 vccd1 _6763_/A sky130_fd_sc_hd__and4_1
XFILLER_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ _4220_/A vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5625_ _5558_/X _7817_/Q _5627_/S vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__mux2_1
X_3886_ _3886_/A vssd1 vssd1 vccd1 vccd1 _8368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8344_ _8345_/CLK _8344_/D vssd1 vssd1 vccd1 vccd1 _8344_/Q sky130_fd_sc_hd__dfxtp_2
X_5556_ _5555_/X _7842_/Q _5562_/S vssd1 vssd1 vccd1 vccd1 _5557_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4507_ _4507_/A _5367_/B vssd1 vssd1 vccd1 vccd1 _4530_/S sky130_fd_sc_hd__nor2_4
X_5487_ _7895_/Q _4220_/A _5491_/S vssd1 vssd1 vccd1 vccd1 _5488_/A sky130_fd_sc_hd__mux2_1
X_8275_ _8275_/CLK _8275_/D vssd1 vssd1 vccd1 vccd1 _8275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7226_ _7226_/A _7226_/B vssd1 vssd1 vccd1 vccd1 _7226_/Y sky130_fd_sc_hd__nand2_1
X_4438_ _4208_/X _8105_/Q _4444_/S vssd1 vssd1 vccd1 vccd1 _4439_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7157_ _8226_/Q _7166_/A vssd1 vssd1 vccd1 vccd1 _7164_/B sky130_fd_sc_hd__xnor2_2
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4369_ _4384_/S vssd1 vssd1 vccd1 vccd1 _4378_/S sky130_fd_sc_hd__buf_2
X_6108_ _7702_/Q _7701_/Q vssd1 vssd1 vccd1 vccd1 _6188_/B sky130_fd_sc_hd__or2b_2
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7088_ _8217_/Q vssd1 vssd1 vccd1 vccd1 _7098_/B sky130_fd_sc_hd__inv_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _6039_/A vssd1 vssd1 vccd1 vccd1 _6039_/X sky130_fd_sc_hd__buf_2
XFILLER_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6674__365 _6674__365/A vssd1 vssd1 vccd1 vccd1 _7949_/CLK sky130_fd_sc_hd__inv_2
X_8414__236 vssd1 vssd1 vccd1 vccd1 partID[10] _8414__236/LO sky130_fd_sc_hd__conb_1
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6635__338 _6635__338/A vssd1 vssd1 vccd1 vccd1 _7919_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3240_ clkbuf_0__3240_/X vssd1 vssd1 vccd1 vccd1 _6583__297/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6390_ _6390_/A vssd1 vssd1 vccd1 vccd1 _7749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5410_ _5410_/A vssd1 vssd1 vccd1 vccd1 _7930_/D sky130_fd_sc_hd__clkbuf_1
Xoutput104 _5908_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__buf_2
Xoutput115 _5915_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__buf_2
X_5341_ _5300_/X _7963_/Q _5345_/S vssd1 vssd1 vccd1 vccd1 _5342_/A sky130_fd_sc_hd__mux2_1
Xoutput159 _5823_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__buf_2
Xoutput126 _5865_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput148 _5845_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__buf_2
Xoutput137 _5887_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__buf_2
X_8060_ _8060_/CLK _8060_/D vssd1 vssd1 vccd1 vccd1 _8060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5272_ _4971_/X _5265_/A _5271_/Y _5214_/X vssd1 vssd1 vccd1 vccd1 _7994_/D sky130_fd_sc_hd__o211a_1
X_4223_ _4223_/A vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__clkbuf_2
X_4154_ _8246_/Q _4084_/X _4158_/S vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4085_ _8270_/Q _4084_/X _4091_/S vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7913_ _7913_/CLK _7913_/D vssd1 vssd1 vccd1 vccd1 _7913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7844_ _7844_/CLK _7844_/D vssd1 vssd1 vccd1 vccd1 _7844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7775_ _7775_/CLK _7775_/D vssd1 vssd1 vccd1 vccd1 _7775_/Q sky130_fd_sc_hd__dfxtp_1
X_6726_ _7421_/A _8331_/Q _8333_/Q vssd1 vssd1 vccd1 vccd1 _7423_/C sky130_fd_sc_hd__a21o_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ _4987_/A vssd1 vssd1 vccd1 vccd1 _5089_/S sky130_fd_sc_hd__buf_4
X_3938_ _8364_/Q vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__buf_2
X_3869_ _3891_/S vssd1 vssd1 vccd1 vccd1 _3882_/S sky130_fd_sc_hd__clkbuf_4
X_6657_ _6675_/A vssd1 vssd1 vccd1 vccd1 _6657_/X sky130_fd_sc_hd__buf_1
X_6931__485 _6931__485/A vssd1 vssd1 vccd1 vccd1 _8082_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3369_ clkbuf_0__3369_/X vssd1 vssd1 vccd1 vccd1 _6863__434/A sky130_fd_sc_hd__clkbuf_4
X_5608_ _5608_/A vssd1 vssd1 vccd1 vccd1 _7825_/D sky130_fd_sc_hd__clkbuf_1
X_6588_ _6650_/A vssd1 vssd1 vccd1 vccd1 _6588_/X sky130_fd_sc_hd__buf_1
X_5539_ _5296_/X _7872_/Q _5539_/S vssd1 vssd1 vccd1 vccd1 _5540_/A sky130_fd_sc_hd__mux2_1
X_8327_ _8327_/CLK _8327_/D vssd1 vssd1 vccd1 vccd1 _8327_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3406_ _7038_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3406_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3723_ clkbuf_0__3723_/X vssd1 vssd1 vccd1 vccd1 _7569__42/A sky130_fd_sc_hd__clkbuf_4
X_8258_ _8258_/CLK _8258_/D vssd1 vssd1 vccd1 vccd1 _8258_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8399_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7209_ _6198_/X _7207_/Y _7198_/X _7194_/X _7208_/Y vssd1 vssd1 vccd1 vccd1 _7210_/B
+ sky130_fd_sc_hd__o32a_1
X_8189_ _8189_/CLK _8189_/D vssd1 vssd1 vccd1 vccd1 _8189_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3199_ _6471_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3199_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3585_ clkbuf_0__3585_/X vssd1 vssd1 vccd1 vccd1 _7306__129/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6973__519 _6974__520/A vssd1 vssd1 vccd1 vccd1 _8116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__clkbuf_1
Xinput39 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__buf_4
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5890_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5899_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4910_ _8030_/Q _4410_/X _4910_/S vssd1 vssd1 vccd1 vccd1 _4911_/A sky130_fd_sc_hd__mux2_1
X_4841_ _4930_/B _4853_/A _4853_/B vssd1 vssd1 vccd1 vccd1 _4851_/B sky130_fd_sc_hd__nand3_1
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4772_ _4863_/B _4749_/X _4757_/X _4771_/X vssd1 vssd1 vccd1 vccd1 _4772_/X sky130_fd_sc_hd__a31o_2
X_7491_ _7491_/A _7491_/B vssd1 vssd1 vccd1 vccd1 _7491_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6373_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6382_/S sky130_fd_sc_hd__clkbuf_2
X_8112_ _8112_/CLK _8112_/D vssd1 vssd1 vccd1 vccd1 _8112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5324_ _5324_/A vssd1 vssd1 vccd1 vccd1 _7971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8043_ _8043_/CLK _8043_/D vssd1 vssd1 vccd1 vccd1 _8043_/Q sky130_fd_sc_hd__dfxtp_1
X_5255_ _5255_/A vssd1 vssd1 vccd1 vccd1 _8001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4206_ _3865_/X _8194_/Q _4218_/S vssd1 vssd1 vccd1 vccd1 _4207_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5186_ _8124_/Q _8132_/Q _5274_/A vssd1 vssd1 vccd1 vccd1 _5186_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_1_0_0__3370_ clkbuf_0__3370_/X vssd1 vssd1 vccd1 vccd1 _6868__438/A sky130_fd_sc_hd__clkbuf_4
X_4137_ _8360_/Q vssd1 vssd1 vccd1 vccd1 _4137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4068_ _4536_/C _4065_/Y _4066_/X _4069_/A vssd1 vssd1 vccd1 vccd1 _4068_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7827_ _7827_/CLK _7827_/D vssd1 vssd1 vccd1 vccd1 _7827_/Q sky130_fd_sc_hd__dfxtp_1
X_7758_ _7758_/CLK _7758_/D vssd1 vssd1 vccd1 vccd1 _7758_/Q sky130_fd_sc_hd__dfxtp_1
X_7689_ _8345_/CLK _7689_/D vssd1 vssd1 vccd1 vccd1 _7689_/Q sky130_fd_sc_hd__dfxtp_1
X_6709_ _8336_/Q _8335_/Q vssd1 vssd1 vccd1 vccd1 _6720_/B sky130_fd_sc_hd__and2_1
XFILLER_7_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__3583_ clkbuf_0__3583_/X vssd1 vssd1 vccd1 vccd1 _7298__123/A sky130_fd_sc_hd__clkbuf_16
XFILLER_15_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6572__288 _6574__290/A vssd1 vssd1 vccd1 vccd1 _7869_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8427__202 vssd1 vssd1 vccd1 vccd1 _8427__202/HI core1Index[2] sky130_fd_sc_hd__conb_1
XFILLER_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _4976_/X _5039_/X _5154_/A vssd1 vssd1 vccd1 vccd1 _5040_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5942_ _7854_/Q _5942_/B vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__and2_1
XFILLER_93_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5873_ _7579_/B _5877_/B vssd1 vssd1 vccd1 vccd1 _5874_/A sky130_fd_sc_hd__or2_1
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7612_ _7612_/A _7615_/B vssd1 vssd1 vccd1 vccd1 _7612_/Y sky130_fd_sc_hd__nor2_1
X_4824_ _8107_/Q _4724_/X _4725_/X _8083_/Q _4622_/A vssd1 vssd1 vccd1 vccd1 _4824_/X
+ sky130_fd_sc_hd__o221a_1
X_7543_ _7543_/A vssd1 vssd1 vccd1 vccd1 _8362_/D sky130_fd_sc_hd__clkbuf_1
X_4755_ _7791_/Q _4676_/X _4754_/X _4729_/X vssd1 vssd1 vccd1 vccd1 _4755_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7474_ _7474_/A vssd1 vssd1 vccd1 vccd1 _7474_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1_0__3206_ clkbuf_0__3206_/X vssd1 vssd1 vccd1 vccd1 _6507__279/A sky130_fd_sc_hd__clkbuf_4
X_4686_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__buf_2
XFILLER_115_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6356_ _5914_/A _7734_/Q _6360_/S vssd1 vssd1 vccd1 vccd1 _6357_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5307_ _7985_/Q vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__clkbuf_2
X_8026_ _8026_/CLK _8026_/D vssd1 vssd1 vccd1 vccd1 _8026_/Q sky130_fd_sc_hd__dfxtp_1
X_6287_ _7618_/A vssd1 vssd1 vccd1 vccd1 _6287_/X sky130_fd_sc_hd__buf_2
XFILLER_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5238_ _7952_/Q _5126_/X _5102_/A _5237_/X vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__o22a_1
X_5169_ _7954_/Q _5126_/X _5102_/A _5168_/X vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7352__166 _7356__170/A vssd1 vssd1 vccd1 vccd1 _8293_/CLK sky130_fd_sc_hd__inv_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clkbuf_opt_2_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7697_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6905__468 _6906__469/A vssd1 vssd1 vccd1 vccd1 _8063_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4540_/A vssd1 vssd1 vccd1 vccd1 _4540_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6986__529 _6987__530/A vssd1 vssd1 vccd1 vccd1 _8126_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4471_ _4486_/S vssd1 vssd1 vccd1 vccd1 _4480_/S sky130_fd_sc_hd__clkbuf_4
X_6141_ _6136_/X _7855_/Q _6134_/X _6137_/X _7679_/Q vssd1 vssd1 vccd1 vccd1 _7679_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6072_/A input2/X _6349_/D vssd1 vssd1 vccd1 vccd1 _6072_/X sky130_fd_sc_hd__or3_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_19 _5905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5023_ _8011_/Q _4955_/X _5271_/B _5022_/X vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__a22o_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _5925_/A _5931_/B vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__and2_1
XFILLER_81_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5856_ _5856_/A vssd1 vssd1 vccd1 vccd1 _5856_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3723_ _7567_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3723_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4807_ _4699_/X _7813_/Q _7797_/Q _4697_/X _4750_/X vssd1 vssd1 vccd1 vccd1 _4807_/X
+ sky130_fd_sc_hd__a221o_1
X_5787_ _7656_/Q _5561_/A _5793_/S vssd1 vssd1 vccd1 vccd1 _5788_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7526_ _8355_/Q _7529_/B _7525_/X _7519_/X vssd1 vssd1 vccd1 vccd1 _8355_/D sky130_fd_sc_hd__o211a_1
X_4738_ _4770_/A _4738_/B _4738_/C vssd1 vssd1 vccd1 vccd1 _4738_/X sky130_fd_sc_hd__or3_1
Xclkbuf_0__3585_ _7302_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3585_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7457_ _7488_/A vssd1 vssd1 vccd1 vccd1 _7470_/A sky130_fd_sc_hd__buf_2
X_4669_ _4667_/X _4668_/X _4669_/S vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__mux2_1
X_7388_ _7388_/A vssd1 vssd1 vccd1 vccd1 _7388_/X sky130_fd_sc_hd__buf_1
XFILLER_103_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ _7730_/Q _6265_/X _6307_/X vssd1 vssd1 vccd1 vccd1 _7730_/D sky130_fd_sc_hd__a21o_1
XFILLER_103_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8009_ _8009_/CLK _8009_/D vssd1 vssd1 vccd1 vccd1 _8009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3405_ clkbuf_0__3405_/X vssd1 vssd1 vccd1 vccd1 _7037__70/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3198_ clkbuf_0__3198_/X vssd1 vssd1 vccd1 vccd1 _6470__250/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7294__120 _7294__120/A vssd1 vssd1 vccd1 vccd1 _8247_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7073__99 _7073__99/A vssd1 vssd1 vccd1 vccd1 _8196_/CLK sky130_fd_sc_hd__inv_2
X_3971_ _3986_/S vssd1 vssd1 vccd1 vccd1 _3980_/S sky130_fd_sc_hd__buf_2
X_5710_ _5710_/A vssd1 vssd1 vccd1 vccd1 _7780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6690_ _8334_/Q _8333_/Q _8332_/Q _8331_/Q vssd1 vssd1 vccd1 vccd1 _6744_/B sky130_fd_sc_hd__and4_2
X_5641_ _7810_/Q _5581_/X _5645_/S vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__mux2_1
X_8360_ _8365_/CLK _8360_/D vssd1 vssd1 vccd1 vccd1 _8360_/Q sky130_fd_sc_hd__dfxtp_4
X_5572_ _5572_/A vssd1 vssd1 vccd1 vccd1 _7837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3370_ _6865_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3370_/X sky130_fd_sc_hd__clkbuf_16
X_4523_ _8360_/Q vssd1 vssd1 vccd1 vccd1 _4523_/X sky130_fd_sc_hd__clkbuf_2
X_8291_ _8291_/CLK _8291_/D vssd1 vssd1 vccd1 vccd1 _8291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7242_ _8225_/Q vssd1 vssd1 vccd1 vccd1 _7242_/Y sky130_fd_sc_hd__inv_2
X_6435__221 _6437__223/A vssd1 vssd1 vccd1 vccd1 _7778_/CLK sky130_fd_sc_hd__inv_2
X_4454_ _4249_/X _8098_/Q _4462_/S vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__mux2_1
X_6847__422 _6847__422/A vssd1 vssd1 vccd1 vccd1 _8017_/CLK sky130_fd_sc_hd__inv_2
X_7173_ _8203_/Q _7173_/B _7173_/C _7173_/D vssd1 vssd1 vccd1 vccd1 _7174_/C sky130_fd_sc_hd__nand4_4
X_4385_ _4385_/A vssd1 vssd1 vccd1 vccd1 _8123_/D sky130_fd_sc_hd__clkbuf_1
X_6124_ _6119_/X _7845_/Q _6116_/X _6120_/X _7669_/Q vssd1 vssd1 vccd1 vccd1 _7669_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__and2_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5006_ _8389_/Q _8328_/Q _8074_/Q _8106_/Q _4995_/A _5181_/A vssd1 vssd1 vccd1 vccd1
+ _5007_/B sky130_fd_sc_hd__mux4_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6957_ _6957_/A vssd1 vssd1 vccd1 vccd1 _6957_/X sky130_fd_sc_hd__buf_1
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5908_ _5908_/A vssd1 vssd1 vccd1 vccd1 _5908_/X sky130_fd_sc_hd__clkbuf_1
X_6854__426 _6858__430/A vssd1 vssd1 vccd1 vccd1 _8021_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5839_ _5839_/A vssd1 vssd1 vccd1 vccd1 _5839_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7509_ _7497_/Y _7506_/X _7508_/X vssd1 vssd1 vccd1 vccd1 _8349_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6787__391 _6791__395/A vssd1 vssd1 vccd1 vccd1 _7976_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3403_ clkbuf_0__3403_/X vssd1 vssd1 vccd1 vccd1 _7025__60/A sky130_fd_sc_hd__clkbuf_16
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4170_ _4170_/A vssd1 vssd1 vccd1 vccd1 _8212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _8349_/CLK _7860_/D vssd1 vssd1 vccd1 vccd1 _7860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6811_ _6811_/A vssd1 vssd1 vccd1 vccd1 _7991_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7791_ _7791_/CLK _7791_/D vssd1 vssd1 vccd1 vccd1 _7791_/Q sky130_fd_sc_hd__dfxtp_1
X_6742_ _6742_/A _6742_/B _6742_/C _6742_/D vssd1 vssd1 vccd1 vccd1 _6743_/D sky130_fd_sc_hd__and4_1
X_3954_ _8360_/Q vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__clkbuf_4
X_3885_ _3884_/X _8368_/Q _3891_/S vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5624_ _5624_/A vssd1 vssd1 vccd1 vccd1 _7818_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3385_ clkbuf_0__3385_/X vssd1 vssd1 vccd1 vccd1 _6937__490/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8343_ _8345_/CLK _8343_/D vssd1 vssd1 vccd1 vccd1 _8343_/Q sky130_fd_sc_hd__dfxtp_1
X_5555_ _5555_/A vssd1 vssd1 vccd1 vccd1 _5555_/X sky130_fd_sc_hd__buf_2
XFILLER_117_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8274_ _8274_/CLK _8274_/D vssd1 vssd1 vccd1 vccd1 _8274_/Q sky130_fd_sc_hd__dfxtp_1
X_4506_ _4506_/A vssd1 vssd1 vccd1 vccd1 _8075_/D sky130_fd_sc_hd__clkbuf_1
X_5486_ _5486_/A vssd1 vssd1 vccd1 vccd1 _7896_/D sky130_fd_sc_hd__clkbuf_1
X_7225_ _7244_/A _7225_/B vssd1 vssd1 vccd1 vccd1 _8219_/D sky130_fd_sc_hd__nor2_1
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4437_ _4437_/A vssd1 vssd1 vccd1 vccd1 _8106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7156_ _8393_/Q _7247_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7156_/X sky130_fd_sc_hd__and3_1
XFILLER_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6107_ _6116_/A vssd1 vssd1 vccd1 vccd1 _6107_/X sky130_fd_sc_hd__buf_6
XFILLER_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _4368_/A _4368_/B vssd1 vssd1 vccd1 vccd1 _4384_/S sky130_fd_sc_hd__or2_4
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7087_ _7110_/C vssd1 vssd1 vccd1 vccd1 _7098_/A sky130_fd_sc_hd__inv_2
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4220_/X _8157_/Q _4303_/S vssd1 vssd1 vccd1 vccd1 _4300_/A sky130_fd_sc_hd__mux2_1
X_6038_ _6051_/A vssd1 vssd1 vccd1 vccd1 _6039_/A sky130_fd_sc_hd__buf_2
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7989_ _7989_/CLK _7989_/D vssd1 vssd1 vccd1 vccd1 _7989_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput105 _5950_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput116 _5917_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__buf_2
X_5340_ _5340_/A vssd1 vssd1 vccd1 vccd1 _7964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput138 _5889_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput127 _5867_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput149 _5848_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_114_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5271_ _5271_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5271_/Y sky130_fd_sc_hd__nand2_1
X_4222_ _4222_/A vssd1 vssd1 vccd1 vccd1 _8189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ _4153_/A vssd1 vssd1 vccd1 vccd1 _8247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4084_ _7990_/Q vssd1 vssd1 vccd1 vccd1 _4084_/X sky130_fd_sc_hd__buf_2
XFILLER_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7019__55 _7019__55/A vssd1 vssd1 vccd1 vccd1 _8152_/CLK sky130_fd_sc_hd__inv_2
X_7912_ _7912_/CLK _7912_/D vssd1 vssd1 vccd1 vccd1 _7912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7843_ _7843_/CLK _7843_/D vssd1 vssd1 vccd1 vccd1 _7843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7774_ _7774_/CLK _7774_/D vssd1 vssd1 vccd1 vccd1 _7774_/Q sky130_fd_sc_hd__dfxtp_1
X_4986_ _5269_/A _4972_/X _4985_/X vssd1 vssd1 vccd1 vccd1 _4986_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6725_ _8333_/Q _7421_/A _8331_/Q vssd1 vssd1 vccd1 vccd1 _6728_/A sky130_fd_sc_hd__nand3_1
X_3937_ _3937_/A vssd1 vssd1 vccd1 vccd1 _8312_/D sky130_fd_sc_hd__clkbuf_1
X_3868_ _5511_/A _5439_/A vssd1 vssd1 vccd1 vccd1 _3891_/S sky130_fd_sc_hd__or2_2
X_3799_ _6036_/A _7538_/B _6214_/A vssd1 vssd1 vccd1 vccd1 _3799_/X sky130_fd_sc_hd__and3_1
X_5607_ _5558_/X _7825_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3368_ clkbuf_0__3368_/X vssd1 vssd1 vccd1 vccd1 _6858__430/A sky130_fd_sc_hd__clkbuf_4
X_6587_ _6851_/A vssd1 vssd1 vccd1 vccd1 _6587_/X sky130_fd_sc_hd__buf_1
XFILLER_105_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5538_ _5538_/A vssd1 vssd1 vccd1 vccd1 _7873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8326_ _8326_/CLK _8326_/D vssd1 vssd1 vccd1 vccd1 _8326_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3405_ _7032_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3405_/X sky130_fd_sc_hd__clkbuf_16
X_8257_ _8257_/CLK _8257_/D vssd1 vssd1 vccd1 vccd1 _8257_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3722_ clkbuf_0__3722_/X vssd1 vssd1 vccd1 vccd1 _7566__40/A sky130_fd_sc_hd__clkbuf_4
X_7208_ _7208_/A vssd1 vssd1 vccd1 vccd1 _7208_/Y sky130_fd_sc_hd__inv_2
X_5469_ _7903_/Q _4220_/A _5473_/S vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__mux2_1
X_8444__219 vssd1 vssd1 vccd1 vccd1 _8444__219/HI partID[1] sky130_fd_sc_hd__conb_1
X_8188_ _8188_/CLK _8188_/D vssd1 vssd1 vccd1 vccd1 _8188_/Q sky130_fd_sc_hd__dfxtp_1
X_7139_ _7207_/A _7207_/B _7422_/A vssd1 vssd1 vccd1 vccd1 _7139_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__3198_ _6465_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3198_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3584_ clkbuf_0__3584_/X vssd1 vssd1 vccd1 vccd1 _7320_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6448__231 _6452__235/A vssd1 vssd1 vccd1 vccd1 _7788_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6680__370 _6680__370/A vssd1 vssd1 vccd1 vccd1 _7954_/CLK sky130_fd_sc_hd__inv_2
X_6641__343 _6641__343/A vssd1 vssd1 vccd1 vccd1 _7924_/CLK sky130_fd_sc_hd__inv_2
X_7316__137 _7316__137/A vssd1 vssd1 vccd1 vccd1 _8264_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7576__48 _7578__50/A vssd1 vssd1 vccd1 vccd1 _8387_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _6053_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _8054_/Q vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__buf_2
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4757_/A _4760_/X _4763_/X _4770_/X _4549_/A vssd1 vssd1 vccd1 vccd1 _4771_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7490_ _7527_/B _7513_/A _7401_/B vssd1 vssd1 vccd1 vccd1 _7490_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6441_ _6453_/A vssd1 vssd1 vccd1 vccd1 _6441_/X sky130_fd_sc_hd__buf_1
X_6372_ _6372_/A vssd1 vssd1 vccd1 vccd1 _7741_/D sky130_fd_sc_hd__clkbuf_1
X_8111_ _8111_/CLK _8111_/D vssd1 vssd1 vccd1 vccd1 _8111_/Q sky130_fd_sc_hd__dfxtp_1
X_5323_ _5300_/X _7971_/Q _5327_/S vssd1 vssd1 vccd1 vccd1 _5324_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8042_ _8042_/CLK _8042_/D vssd1 vssd1 vccd1 vccd1 _8042_/Q sky130_fd_sc_hd__dfxtp_1
X_5254_ _5250_/B _5254_/B _7547_/A vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__and3b_1
X_5185_ _5271_/A _5182_/X _5184_/X vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__o21a_1
X_4205_ _4227_/S vssd1 vssd1 vccd1 vccd1 _4218_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4136_ _4136_/A vssd1 vssd1 vccd1 vccd1 _8252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4067_ _8049_/Q _8054_/Q vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__or2b_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7826_ _7826_/CLK _7826_/D vssd1 vssd1 vccd1 vccd1 _7826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4969_ _5100_/A vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__clkbuf_4
X_7757_ _7757_/CLK _7757_/D vssd1 vssd1 vccd1 vccd1 _7757_/Q sky130_fd_sc_hd__dfxtp_1
X_7688_ _8345_/CLK _7688_/D vssd1 vssd1 vccd1 vccd1 _7688_/Q sky130_fd_sc_hd__dfxtp_1
X_6708_ _7411_/A _7411_/B _8399_/Q vssd1 vssd1 vccd1 vccd1 _6742_/A sky130_fd_sc_hd__a21bo_1
XFILLER_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8309_ _8309_/CLK _8309_/D vssd1 vssd1 vccd1 vccd1 _8309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6949__500 _6949__500/A vssd1 vssd1 vccd1 vccd1 _8097_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6648__349 _6649__350/A vssd1 vssd1 vccd1 vccd1 _7930_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ _5941_/A vssd1 vssd1 vccd1 vccd1 _5941_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5872_ _5872_/A vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7012_/A
+ sky130_fd_sc_hd__clkbuf_16
X_7611_ _7614_/A _7611_/B vssd1 vssd1 vccd1 vccd1 _7611_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4823_ _8075_/Q _4716_/X _4687_/X _8038_/Q vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__a22o_1
X_7542_ _7629_/A _7629_/B _7549_/C vssd1 vssd1 vccd1 vccd1 _7543_/A sky130_fd_sc_hd__and3_1
X_4754_ _4730_/X _7887_/Q _7831_/Q _4731_/X vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7473_ _7482_/A _7473_/B vssd1 vssd1 vccd1 vccd1 _8338_/D sky130_fd_sc_hd__nor2_1
X_6590__301 _6592__303/A vssd1 vssd1 vccd1 vccd1 _7882_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3205_ clkbuf_0__3205_/X vssd1 vssd1 vccd1 vccd1 _6581_/A sky130_fd_sc_hd__clkbuf_4
X_4685_ _4750_/A vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__buf_2
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6355_ _6355_/A vssd1 vssd1 vccd1 vccd1 _7733_/D sky130_fd_sc_hd__clkbuf_1
X_6286_ _6312_/A vssd1 vssd1 vccd1 vccd1 _6337_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5306_ _5306_/A vssd1 vssd1 vccd1 vccd1 _7978_/D sky130_fd_sc_hd__clkbuf_1
X_8025_ _8025_/CLK _8025_/D vssd1 vssd1 vccd1 vccd1 _8025_/Q sky130_fd_sc_hd__dfxtp_1
X_5237_ _7917_/Q _7925_/Q _5237_/S vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6781__386 _6782__387/A vssd1 vssd1 vccd1 vccd1 _7971_/CLK sky130_fd_sc_hd__inv_2
X_5168_ _7919_/Q _7927_/Q _5237_/S vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4119_ _4119_/A vssd1 vssd1 vccd1 vccd1 _8257_/D sky130_fd_sc_hd__clkbuf_1
X_5099_ _7994_/Q _5100_/B vssd1 vssd1 vccd1 vccd1 _5115_/A sky130_fd_sc_hd__or2_1
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _7809_/CLK _7809_/D vssd1 vssd1 vccd1 vccd1 _7809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6654__353 _6655__354/A vssd1 vssd1 vccd1 vccd1 _7934_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4470_ _4912_/A _4875_/A vssd1 vssd1 vccd1 vccd1 _4486_/S sky130_fd_sc_hd__or2_2
XFILLER_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6140_ _6136_/X _7854_/Q _6134_/X _6137_/X _7678_/Q vssd1 vssd1 vccd1 vccd1 _7678_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _7692_/Q _6061_/X _6039_/A _6070_/X vssd1 vssd1 vccd1 vccd1 _6071_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _4986_/X _5000_/X _5002_/X _5021_/X vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__a31o_2
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5924_ _5924_/A vssd1 vssd1 vccd1 vccd1 _5924_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5855_ _7611_/B _5855_/B vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__or2_1
Xclkbuf_0__3722_ _7561_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3722_/X sky130_fd_sc_hd__clkbuf_16
X_4806_ _4344_/X _4538_/A _4805_/X _4774_/X vssd1 vssd1 vccd1 vccd1 _8058_/D sky130_fd_sc_hd__o211a_1
X_5786_ _5786_/A vssd1 vssd1 vccd1 vccd1 _7657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7525_ _8356_/Q _7527_/B _7513_/A vssd1 vssd1 vccd1 vccd1 _7525_/X sky130_fd_sc_hd__or3b_1
X_4737_ _7972_/Q _4681_/A _4642_/A _4736_/X vssd1 vssd1 vccd1 vccd1 _4738_/C sky130_fd_sc_hd__o211a_1
Xclkbuf_0__3584_ _7301_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3584_/X sky130_fd_sc_hd__clkbuf_16
X_7456_ _7456_/A vssd1 vssd1 vccd1 vccd1 _7488_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4668_ _8026_/Q _7981_/Q _7841_/Q _8209_/Q _4596_/A _4595_/X vssd1 vssd1 vccd1 vccd1
+ _4668_/X sky130_fd_sc_hd__mux4_1
X_6407_ _6107_/X _6188_/B _7610_/A vssd1 vssd1 vccd1 vccd1 _7756_/D sky130_fd_sc_hd__a21oi_1
XFILLER_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ _4593_/S _4598_/X _4802_/A vssd1 vssd1 vccd1 vccd1 _4599_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6338_ _7729_/Q _6320_/A _6324_/X _6337_/X vssd1 vssd1 vccd1 vccd1 _7729_/D sky130_fd_sc_hd__a211o_1
XFILLER_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6269_ _6841_/C _6254_/Y _6268_/X _6289_/B vssd1 vssd1 vccd1 vccd1 _6270_/C sky130_fd_sc_hd__a22o_1
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8008_ _8008_/CLK _8008_/D vssd1 vssd1 vccd1 vccd1 _8008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3404_ clkbuf_0__3404_/X vssd1 vssd1 vccd1 vccd1 _7029__63/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6597__307 _6597__307/A vssd1 vssd1 vccd1 vccd1 _7888_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3197_ clkbuf_0__3197_/X vssd1 vssd1 vccd1 vccd1 _6462__243/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7058__86 _7062__90/A vssd1 vssd1 vccd1 vccd1 _8183_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _3989_/B _5367_/B vssd1 vssd1 vccd1 vccd1 _3986_/S sky130_fd_sc_hd__nor2_2
XFILLER_16_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6992__534 _6993__535/A vssd1 vssd1 vccd1 vccd1 _8131_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5640_ _5640_/A vssd1 vssd1 vccd1 vccd1 _7811_/D sky130_fd_sc_hd__clkbuf_1
X_5571_ _5570_/X _7837_/Q _5571_/S vssd1 vssd1 vccd1 vccd1 _5572_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8290_ _8290_/CLK _8290_/D vssd1 vssd1 vccd1 vccd1 _8290_/Q sky130_fd_sc_hd__dfxtp_1
X_4522_ _4522_/A vssd1 vssd1 vccd1 vccd1 _8070_/D sky130_fd_sc_hd__clkbuf_1
X_7241_ _7244_/A _7241_/B vssd1 vssd1 vccd1 vccd1 _8224_/D sky130_fd_sc_hd__nor2_1
X_4453_ _4468_/S vssd1 vssd1 vccd1 vccd1 _4462_/S sky130_fd_sc_hd__buf_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7172_ _7252_/B _7202_/B _7283_/B _7262_/C vssd1 vssd1 vccd1 vccd1 _7174_/B sky130_fd_sc_hd__a211o_1
X_4384_ _4226_/X _8123_/Q _4384_/S vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__mux2_1
X_6123_ _6119_/X _7700_/Q _6116_/X _6120_/X _7668_/Q vssd1 vssd1 vccd1 vccd1 _7668_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _7684_/Q _6048_/X _6051_/X _6053_/X vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__o22a_4
XFILLER_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5005_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__buf_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6585__299 _6586__300/A vssd1 vssd1 vccd1 vccd1 _7880_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6442__226 _6443__227/A vssd1 vssd1 vccd1 vccd1 _7783_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5907_ _5907_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5908_/A sky130_fd_sc_hd__and2_1
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5838_ _6199_/B _5844_/B vssd1 vssd1 vccd1 vccd1 _5839_/A sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__3599_ clkbuf_0__3599_/X vssd1 vssd1 vccd1 vccd1 _7381__15/A sky130_fd_sc_hd__clkbuf_4
X_5769_ _5558_/X _7708_/Q _5771_/S vssd1 vssd1 vccd1 vccd1 _5770_/A sky130_fd_sc_hd__mux2_1
X_7508_ _7507_/Y _7490_/Y _7456_/A vssd1 vssd1 vccd1 vccd1 _7508_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7439_ _7450_/B _7439_/B _7439_/C vssd1 vssd1 vccd1 vccd1 _7442_/A sky130_fd_sc_hd__nand3_1
XFILLER_116_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6605__314 _6606__315/A vssd1 vssd1 vccd1 vccd1 _7895_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3402_ clkbuf_0__3402_/X vssd1 vssd1 vccd1 vccd1 _7016__52/A sky130_fd_sc_hd__clkbuf_16
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3249_ clkbuf_0__3249_/X vssd1 vssd1 vccd1 vccd1 _6622__327/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6497__271 _6501__275/A vssd1 vssd1 vccd1 vccd1 _7828_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6810_ _8356_/Q _6810_/B vssd1 vssd1 vccd1 vccd1 _6811_/A sky130_fd_sc_hd__and2_1
XFILLER_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6506__278 _6507__279/A vssd1 vssd1 vccd1 vccd1 _7835_/CLK sky130_fd_sc_hd__inv_2
X_7790_ _7790_/CLK _7790_/D vssd1 vssd1 vccd1 vccd1 _7790_/Q sky130_fd_sc_hd__dfxtp_1
X_6741_ _7621_/A _6714_/B _6718_/Y _6719_/X _6740_/X vssd1 vssd1 vccd1 vccd1 _6742_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _3953_/A vssd1 vssd1 vccd1 vccd1 _8308_/D sky130_fd_sc_hd__clkbuf_1
X_3884_ _8360_/Q vssd1 vssd1 vccd1 vccd1 _3884_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5623_ _5555_/X _7818_/Q _5627_/S vssd1 vssd1 vccd1 vccd1 _5624_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3384_ clkbuf_0__3384_/X vssd1 vssd1 vccd1 vccd1 _6931__485/A sky130_fd_sc_hd__clkbuf_4
X_6814__400 _6814__400/A vssd1 vssd1 vccd1 vccd1 _7993_/CLK sky130_fd_sc_hd__inv_2
X_8342_ _8342_/CLK _8342_/D vssd1 vssd1 vccd1 vccd1 _8342_/Q sky130_fd_sc_hd__dfxtp_1
X_5554_ _5554_/A vssd1 vssd1 vccd1 vccd1 _7843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8273_ _8273_/CLK _8273_/D vssd1 vssd1 vccd1 vccd1 _8273_/Q sky130_fd_sc_hd__dfxtp_1
X_4505_ _4347_/X _8075_/Q _4505_/S vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__mux2_1
X_5485_ _7896_/Q _4217_/A _5485_/S vssd1 vssd1 vccd1 vccd1 _5486_/A sky130_fd_sc_hd__mux2_1
X_7224_ _7220_/X _7221_/Y _7222_/X _7223_/X _7092_/A vssd1 vssd1 vccd1 vccd1 _7225_/B
+ sky130_fd_sc_hd__o32a_1
X_4436_ _4249_/X _8106_/Q _4444_/S vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7155_ _7247_/A _7247_/B _7596_/A vssd1 vssd1 vccd1 vccd1 _7155_/Y sky130_fd_sc_hd__a21oi_1
X_4367_ _4367_/A vssd1 vssd1 vccd1 vccd1 _8131_/D sky130_fd_sc_hd__clkbuf_1
X_6106_ _6125_/A vssd1 vssd1 vccd1 vccd1 _6116_/A sky130_fd_sc_hd__buf_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6860__431 _6864__435/A vssd1 vssd1 vccd1 vccd1 _8026_/CLK sky130_fd_sc_hd__inv_2
X_7086_ _8218_/Q vssd1 vssd1 vccd1 vccd1 _7110_/C sky130_fd_sc_hd__clkbuf_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4298_/A vssd1 vssd1 vccd1 vccd1 _8158_/D sky130_fd_sc_hd__clkbuf_1
X_6037_ _7730_/Q _6349_/D _7540_/A vssd1 vssd1 vccd1 vccd1 _6051_/A sky130_fd_sc_hd__a21o_2
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ _7989_/CLK _7988_/D vssd1 vssd1 vccd1 vccd1 _7988_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 _5952_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput139 _5892_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput128 _5870_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput117 _5919_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__buf_2
XFILLER_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5270_ _5187_/X _5265_/A _5269_/Y _5214_/X vssd1 vssd1 vccd1 vccd1 _7995_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4221_ _4220_/X _8189_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4152_ _8247_/Q _4081_/X _4158_/S vssd1 vssd1 vccd1 vccd1 _4153_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4083_ _4083_/A vssd1 vssd1 vccd1 vccd1 _8271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7911_ _7911_/CLK _7911_/D vssd1 vssd1 vccd1 vccd1 _7911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7842_ _7842_/CLK _7842_/D vssd1 vssd1 vccd1 vccd1 _7842_/Q sky130_fd_sc_hd__dfxtp_1
X_4985_ _4976_/X _4979_/X _5154_/A vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7773_ _7773_/CLK _7773_/D vssd1 vssd1 vccd1 vccd1 _7773_/Q sky130_fd_sc_hd__dfxtp_1
X_6724_ _8332_/Q vssd1 vssd1 vccd1 vccd1 _7421_/A sky130_fd_sc_hd__clkbuf_2
X_3936_ _8312_/Q _3772_/X _3952_/S vssd1 vssd1 vccd1 vccd1 _3937_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3867_ _3867_/A _5261_/A _3968_/B _3967_/A vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__or4b_4
X_5606_ _5606_/A vssd1 vssd1 vccd1 vccd1 _7826_/D sky130_fd_sc_hd__clkbuf_1
X_3798_ _7755_/Q _7754_/Q vssd1 vssd1 vccd1 vccd1 _6214_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1_0__3367_ clkbuf_0__3367_/X vssd1 vssd1 vccd1 vccd1 _6877_/A sky130_fd_sc_hd__clkbuf_4
X_5537_ _5292_/X _7873_/Q _5539_/S vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3404_ _7026_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3404_/X sky130_fd_sc_hd__clkbuf_16
X_8325_ _8325_/CLK _8325_/D vssd1 vssd1 vccd1 vccd1 _8325_/Q sky130_fd_sc_hd__dfxtp_1
X_8256_ _8256_/CLK _8256_/D vssd1 vssd1 vccd1 vccd1 _8256_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3721_ clkbuf_0__3721_/X vssd1 vssd1 vccd1 vccd1 _7559__34/A sky130_fd_sc_hd__clkbuf_4
X_7207_ _7207_/A _7207_/B vssd1 vssd1 vccd1 vccd1 _7207_/Y sky130_fd_sc_hd__nand2_1
X_5468_ _5468_/A vssd1 vssd1 vccd1 vccd1 _7904_/D sky130_fd_sc_hd__clkbuf_1
X_4419_ _4419_/A vssd1 vssd1 vccd1 vccd1 _8114_/D sky130_fd_sc_hd__clkbuf_1
X_5399_ _7934_/Q _4526_/X _5401_/S vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__mux2_1
X_8187_ _8187_/CLK _8187_/D vssd1 vssd1 vccd1 vccd1 _8187_/Q sky130_fd_sc_hd__dfxtp_1
X_7138_ _8405_/Q _7207_/A _7207_/B vssd1 vssd1 vccd1 vccd1 _7138_/X sky130_fd_sc_hd__and3_1
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3197_ _6459_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3197_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7069_ _7069_/A vssd1 vssd1 vccd1 vccd1 _7069_/X sky130_fd_sc_hd__buf_1
XFILLER_100_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8335_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _6055_/A sky130_fd_sc_hd__clkbuf_1
X_8418__193 vssd1 vssd1 vccd1 vccd1 _8418__193/HI core0Index[0] sky130_fd_sc_hd__conb_1
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6867__437 _6868__438/A vssd1 vssd1 vccd1 vccd1 _8032_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _4770_/A _4770_/B _4770_/C vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__or3_1
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6440_ _6471_/A vssd1 vssd1 vccd1 vccd1 _6440_/X sky130_fd_sc_hd__buf_1
X_6371_ _5929_/A _7741_/Q _6371_/S vssd1 vssd1 vccd1 vccd1 _6372_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5322_ _5322_/A vssd1 vssd1 vccd1 vccd1 _7972_/D sky130_fd_sc_hd__clkbuf_1
X_8110_ _8110_/CLK _8110_/D vssd1 vssd1 vccd1 vccd1 _8110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5253_ _6838_/A vssd1 vssd1 vccd1 vccd1 _7547_/A sky130_fd_sc_hd__clkbuf_2
X_8041_ _8041_/CLK _8041_/D vssd1 vssd1 vccd1 vccd1 _8041_/Q sky130_fd_sc_hd__dfxtp_1
X_5184_ _8092_/Q _5098_/X _5183_/X _8250_/Q _4990_/X vssd1 vssd1 vccd1 vccd1 _5184_/X
+ sky130_fd_sc_hd__o221a_1
X_4204_ _5511_/B _4204_/B vssd1 vssd1 vccd1 vccd1 _4227_/S sky130_fd_sc_hd__or2_2
XFILLER_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4135_ _8252_/Q _4134_/X _4135_/S vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4066_ _4536_/C _4063_/A vssd1 vssd1 vccd1 vccd1 _4066_/X sky130_fd_sc_hd__or2b_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7825_ _7825_/CLK _7825_/D vssd1 vssd1 vccd1 vccd1 _7825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7756_ _8391_/CLK _7756_/D vssd1 vssd1 vccd1 vccd1 _7756_/Q sky130_fd_sc_hd__dfxtp_1
X_4968_ _5231_/S vssd1 vssd1 vccd1 vccd1 _5198_/S sky130_fd_sc_hd__clkbuf_4
X_4899_ _4899_/A vssd1 vssd1 vccd1 vccd1 _8036_/D sky130_fd_sc_hd__clkbuf_1
X_7687_ _8345_/CLK _7687_/D vssd1 vssd1 vccd1 vccd1 _7687_/Q sky130_fd_sc_hd__dfxtp_1
X_6707_ _6702_/B _6702_/C _8339_/Q vssd1 vssd1 vccd1 vccd1 _7411_/B sky130_fd_sc_hd__a21o_1
X_3919_ _3919_/A vssd1 vssd1 vccd1 vccd1 _8320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6638_ _6644_/A vssd1 vssd1 vccd1 vccd1 _6638_/X sky130_fd_sc_hd__buf_1
XFILLER_118_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6569_ _6569_/A vssd1 vssd1 vccd1 vccd1 _7867_/D sky130_fd_sc_hd__clkbuf_1
X_8308_ _8308_/CLK _8308_/D vssd1 vssd1 vccd1 vccd1 _8308_/Q sky130_fd_sc_hd__dfxtp_1
X_7322__142 _7322__142/A vssd1 vssd1 vccd1 vccd1 _8269_/CLK sky130_fd_sc_hd__inv_2
X_6827__410 _6827__410/A vssd1 vssd1 vccd1 vccd1 _8003_/CLK sky130_fd_sc_hd__inv_2
X_8239_ _8239_/CLK _8239_/D vssd1 vssd1 vccd1 vccd1 _8239_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3249_ _6620_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3249_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6914__471 _6914__471/A vssd1 vssd1 vccd1 vccd1 _8068_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5940_ _7853_/Q _5942_/B vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__and2_1
XFILLER_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6956__505 _6956__505/A vssd1 vssd1 vccd1 vccd1 _8102_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5871_ _7584_/B _5877_/B vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__or2_1
X_7610_ _7610_/A _7610_/B vssd1 vssd1 vccd1 vccd1 _8397_/D sky130_fd_sc_hd__nor2_1
X_4822_ _4750_/X _4820_/X _4821_/X vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__o21a_1
X_7541_ _7549_/B vssd1 vssd1 vccd1 vccd1 _7629_/B sky130_fd_sc_hd__clkbuf_2
X_4753_ _4750_/X _4751_/X _4752_/X vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__o21a_1
X_7472_ _6711_/Y _7447_/B _7461_/X _6714_/B vssd1 vssd1 vccd1 vccd1 _7473_/B sky130_fd_sc_hd__o22a_1
Xclkbuf_1_1_0__3204_ clkbuf_0__3204_/X vssd1 vssd1 vccd1 vccd1 _6501__275/A sky130_fd_sc_hd__clkbuf_4
X_4684_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4750_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6354_ _5912_/A _6909_/A _6360_/S vssd1 vssd1 vccd1 vccd1 _6355_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6285_ _6285_/A _6285_/B vssd1 vssd1 vccd1 vccd1 _6312_/A sky130_fd_sc_hd__nor2_2
X_5305_ _5304_/X _7978_/Q _5309_/S vssd1 vssd1 vccd1 vccd1 _5306_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8024_ _8024_/CLK _8024_/D vssd1 vssd1 vccd1 vccd1 _8024_/Q sky130_fd_sc_hd__dfxtp_1
X_5236_ _5218_/A _5234_/X _5235_/X vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _5218_/A _5165_/X _5166_/X vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4118_ _8257_/Q _3963_/X _4118_/S vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__mux2_1
X_5098_ _5150_/A vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4049_ _8052_/Q vssd1 vssd1 vccd1 vccd1 _4843_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7808_ _7808_/CLK _7808_/D vssd1 vssd1 vccd1 vccd1 _7808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7739_ _8066_/CLK _7739_/D vssd1 vssd1 vccd1 vccd1 _7739_/Q sky130_fd_sc_hd__dfxtp_1
X_7554__30 _7554__30/A vssd1 vssd1 vccd1 vccd1 _8369_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6491__266 _6492__267/A vssd1 vssd1 vccd1 vccd1 _7823_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7329__148 _7329__148/A vssd1 vssd1 vccd1 vccd1 _8275_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__and2_1
XFILLER_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5021_ _5007_/X _5013_/X _5018_/X _5019_/X _5095_/A vssd1 vssd1 vccd1 vccd1 _5021_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5923_ _5923_/A _5931_/B vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__and2_1
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5854_ _5854_/A vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3721_ _7555_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3721_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4805_ _4540_/A _8058_/Q _4632_/X _4804_/X _4605_/A vssd1 vssd1 vccd1 vccd1 _4805_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7524_ _8354_/Q _7511_/X _7523_/X _7519_/X vssd1 vssd1 vccd1 vccd1 _8354_/D sky130_fd_sc_hd__o211a_1
X_5785_ _7657_/Q _5558_/A _5785_/S vssd1 vssd1 vccd1 vccd1 _5786_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4736_ _8033_/Q _4676_/A _4735_/X _4750_/A vssd1 vssd1 vccd1 vccd1 _4736_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_0__3583_ _7295_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3583_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4667_ _8119_/Q _7889_/Q _7833_/Q _7793_/Q _4579_/A _4595_/X vssd1 vssd1 vccd1 vccd1
+ _4667_/X sky130_fd_sc_hd__mux4_1
X_7455_ _3814_/X _6287_/X _7531_/C _6118_/A vssd1 vssd1 vccd1 vccd1 _7456_/A sky130_fd_sc_hd__a31o_2
X_6406_ _6406_/A vssd1 vssd1 vccd1 vccd1 _7755_/D sky130_fd_sc_hd__clkbuf_1
X_6337_ _7170_/A _6337_/B _7943_/Q _6337_/D vssd1 vssd1 vccd1 vccd1 _6337_/X sky130_fd_sc_hd__and4_1
XFILLER_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4598_ _8202_/Q _7820_/Q _7804_/Q _7788_/Q _4595_/A _4559_/A vssd1 vssd1 vccd1 vccd1
+ _4598_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6268_ _8060_/Q _6231_/A _7618_/A _6244_/A vssd1 vssd1 vccd1 vccd1 _6268_/X sky130_fd_sc_hd__a31o_1
X_6199_ _6687_/A _6199_/B _6214_/A vssd1 vssd1 vccd1 vccd1 _7533_/B sky130_fd_sc_hd__and3_2
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8007_ _8007_/CLK _8007_/D vssd1 vssd1 vccd1 vccd1 _8007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5219_ _8313_/Q _5187_/X _5125_/X _8305_/Q _5089_/S vssd1 vssd1 vccd1 vccd1 _5219_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3196_ clkbuf_0__3196_/X vssd1 vssd1 vccd1 vccd1 _6458__240/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7335__152 _7336__153/A vssd1 vssd1 vccd1 vccd1 _8279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5570_ _5570_/A vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ _8070_/Q _4520_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7240_ _7220_/X _7115_/B _7222_/X _7223_/X _7113_/Y vssd1 vssd1 vccd1 vccd1 _7241_/B
+ sky130_fd_sc_hd__o32a_1
X_4452_ _5348_/A _5457_/B vssd1 vssd1 vccd1 vccd1 _4468_/S sky130_fd_sc_hd__or2_2
X_7171_ _7265_/A _7265_/B vssd1 vssd1 vccd1 vccd1 _7283_/B sky130_fd_sc_hd__nor2_2
X_4383_ _4383_/A vssd1 vssd1 vccd1 vccd1 _8124_/D sky130_fd_sc_hd__clkbuf_1
X_6122_ _6119_/X _7699_/Q _6116_/X _6120_/X _7667_/Q vssd1 vssd1 vccd1 vccd1 _7667_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A _6062_/B vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__and2_1
XFILLER_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927__481 _6928__482/A vssd1 vssd1 vccd1 vccd1 _8078_/CLK sky130_fd_sc_hd__inv_2
X_5004_ _5237_/S vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__buf_4
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5906_ _5906_/A vssd1 vssd1 vccd1 vccd1 _5906_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5837_ _5837_/A vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3598_ clkbuf_0__3598_/X vssd1 vssd1 vccd1 vccd1 _7372__7/A sky130_fd_sc_hd__clkbuf_4
X_5768_ _5768_/A vssd1 vssd1 vccd1 vccd1 _7709_/D sky130_fd_sc_hd__clkbuf_1
X_7507_ _8349_/Q vssd1 vssd1 vccd1 vccd1 _7507_/Y sky130_fd_sc_hd__inv_2
X_4719_ _4724_/A vssd1 vssd1 vccd1 vccd1 _4719_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7438_ _7439_/B _7474_/A _7450_/B vssd1 vssd1 vccd1 vccd1 _7440_/B sky130_fd_sc_hd__a21o_1
X_5699_ _7784_/Q _5587_/X _5699_/S vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3248_ clkbuf_0__3248_/X vssd1 vssd1 vccd1 vccd1 _6632_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6794__397 _6796__399/A vssd1 vssd1 vccd1 vccd1 _7982_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6740_ _6722_/Y _6723_/X _6735_/X _6737_/X _6739_/X vssd1 vssd1 vccd1 vccd1 _6740_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3952_ _8308_/Q _3951_/X _3952_/S vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__mux2_1
X_3883_ _3883_/A vssd1 vssd1 vccd1 vccd1 _8369_/D sky130_fd_sc_hd__clkbuf_1
X_5622_ _5622_/A vssd1 vssd1 vccd1 vccd1 _7819_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3383_ clkbuf_0__3383_/X vssd1 vssd1 vccd1 vccd1 _6922__477/A sky130_fd_sc_hd__clkbuf_4
X_8341_ _8341_/CLK _8341_/D vssd1 vssd1 vccd1 vccd1 _8341_/Q sky130_fd_sc_hd__dfxtp_2
X_5553_ _5552_/X _7843_/Q _5562_/S vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__mux2_1
X_4504_ _4504_/A vssd1 vssd1 vccd1 vccd1 _8076_/D sky130_fd_sc_hd__clkbuf_1
X_8272_ _8272_/CLK _8272_/D vssd1 vssd1 vccd1 vccd1 _8272_/Q sky130_fd_sc_hd__dfxtp_1
X_5484_ _5484_/A vssd1 vssd1 vccd1 vccd1 _7897_/D sky130_fd_sc_hd__clkbuf_1
X_7223_ _7237_/B vssd1 vssd1 vccd1 vccd1 _7223_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4435_ _4450_/S vssd1 vssd1 vccd1 vccd1 _4444_/S sky130_fd_sc_hd__buf_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7154_ _8226_/Q _7166_/A _8227_/Q vssd1 vssd1 vccd1 vccd1 _7247_/B sky130_fd_sc_hd__a21o_1
X_4366_ _8131_/Q _4143_/X _4366_/S vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__mux2_1
X_6105_ _7701_/Q _7702_/Q vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__or2b_1
XFILLER_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _8219_/Q vssd1 vssd1 vccd1 vccd1 _7092_/A sky130_fd_sc_hd__inv_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4217_/X _8158_/Q _4297_/S vssd1 vssd1 vccd1 vccd1 _4298_/A sky130_fd_sc_hd__mux2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A vssd1 vssd1 vccd1 vccd1 _7540_/A sky130_fd_sc_hd__inv_2
X_6821__405 _6821__405/A vssd1 vssd1 vccd1 vccd1 _7998_/CLK sky130_fd_sc_hd__inv_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ _8065_/CLK _7987_/D vssd1 vssd1 vccd1 vccd1 _7987_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6938_ _6938_/A vssd1 vssd1 vccd1 vccd1 _6938_/X sky130_fd_sc_hd__buf_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 _5954_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput129 _5872_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput118 _5921_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__buf_2
XFILLER_114_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4220_ _4220_/A vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__clkbuf_2
X_6512__283 _6514__285/A vssd1 vssd1 vccd1 vccd1 _7840_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4151_ _4151_/A vssd1 vssd1 vccd1 vccd1 _8248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4082_ _8271_/Q _4081_/X _4091_/S vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__mux2_1
X_7910_ _7910_/CLK _7910_/D vssd1 vssd1 vccd1 vccd1 _7910_/Q sky130_fd_sc_hd__dfxtp_1
X_7841_ _7841_/CLK _7841_/D vssd1 vssd1 vccd1 vccd1 _7841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7772_ _7772_/CLK _7772_/D vssd1 vssd1 vccd1 vccd1 _7772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _5243_/A vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__clkbuf_2
X_6723_ _8402_/Q _7429_/A _7429_/B vssd1 vssd1 vccd1 vccd1 _6723_/X sky130_fd_sc_hd__and3_1
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3935_ _3964_/S vssd1 vssd1 vccd1 vccd1 _3952_/S sky130_fd_sc_hd__buf_2
X_5605_ _5555_/X _7826_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__mux2_1
X_3866_ _6340_/B _8012_/Q vssd1 vssd1 vccd1 vccd1 _3968_/B sky130_fd_sc_hd__nand2b_2
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3797_ _4052_/A vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3366_ clkbuf_0__3366_/X vssd1 vssd1 vccd1 vccd1 _6883_/A sky130_fd_sc_hd__clkbuf_4
X_5536_ _5536_/A vssd1 vssd1 vccd1 vccd1 _7874_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3403_ _7020_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3403_/X sky130_fd_sc_hd__clkbuf_16
X_8324_ _8324_/CLK _8324_/D vssd1 vssd1 vccd1 vccd1 _8324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8255_ _8255_/CLK _8255_/D vssd1 vssd1 vccd1 vccd1 _8255_/Q sky130_fd_sc_hd__dfxtp_1
X_5467_ _7904_/Q _4217_/A _5467_/S vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__mux2_1
X_4418_ _8114_/Q _4386_/X _4426_/S vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__mux2_1
X_7206_ _7218_/A _7206_/B vssd1 vssd1 vccd1 vccd1 _8214_/D sky130_fd_sc_hd__nor2_1
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8186_ _8186_/CLK _8186_/D vssd1 vssd1 vccd1 vccd1 _8186_/Q sky130_fd_sc_hd__dfxtp_1
X_5398_ _5398_/A vssd1 vssd1 vccd1 vccd1 _7935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7137_ _7204_/A _7140_/B _7208_/A vssd1 vssd1 vccd1 vccd1 _7207_/B sky130_fd_sc_hd__a21o_1
Xclkbuf_0__3196_ _6453_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3196_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4349_ _4349_/A vssd1 vssd1 vccd1 vccd1 _8139_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3582_ clkbuf_0__3582_/X vssd1 vssd1 vccd1 vccd1 _7291__117/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6019_ _7726_/Q input8/X _6025_/S vssd1 vssd1 vccd1 vccd1 _6019_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6455__237 _6457__239/A vssd1 vssd1 vccd1 vccd1 _7794_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6618__325 _6618__325/A vssd1 vssd1 vccd1 vccd1 _7906_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6370_ _6370_/A vssd1 vssd1 vccd1 vccd1 _7740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _5296_/X _7972_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5322_/A sky130_fd_sc_hd__mux2_1
X_8040_ _8040_/CLK _8040_/D vssd1 vssd1 vccd1 vccd1 _8040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5252_ _5249_/B _5261_/B _5347_/B vssd1 vssd1 vccd1 vccd1 _5254_/B sky130_fd_sc_hd__a21o_1
X_5183_ _5183_/A vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__clkbuf_2
X_4203_ _4203_/A vssd1 vssd1 vccd1 vccd1 _8195_/D sky130_fd_sc_hd__clkbuf_1
X_4134_ _8361_/Q vssd1 vssd1 vccd1 vccd1 _4134_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4065_ _4853_/A _4069_/B vssd1 vssd1 vccd1 vccd1 _4065_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7824_ _7824_/CLK _7824_/D vssd1 vssd1 vccd1 vccd1 _7824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7755_ _8065_/CLK _7755_/D vssd1 vssd1 vccd1 vccd1 _7755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _5240_/S vssd1 vssd1 vccd1 vccd1 _5231_/S sky130_fd_sc_hd__buf_2
X_4898_ _8036_/Q _4392_/X _4904_/S vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__mux2_1
X_7686_ _8345_/CLK _7686_/D vssd1 vssd1 vccd1 vccd1 _7686_/Q sky130_fd_sc_hd__dfxtp_1
X_6706_ _8395_/Q _6706_/B vssd1 vssd1 vccd1 vccd1 _7409_/A sky130_fd_sc_hd__xor2_1
X_3918_ _3865_/X _8320_/Q _3926_/S vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8450__225 vssd1 vssd1 vccd1 vccd1 _8450__225/HI partID[13] sky130_fd_sc_hd__conb_1
X_3849_ _3849_/A vssd1 vssd1 vccd1 vccd1 _8381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6568_ _7867_/Q _5901_/A _6570_/S vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5519_ _7881_/Q _4214_/A _5521_/S vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__mux2_1
X_8307_ _8307_/CLK _8307_/D vssd1 vssd1 vccd1 vccd1 _8307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8238_ _8239_/CLK _8238_/D vssd1 vssd1 vccd1 vccd1 _8238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8169_ _8169_/CLK _8169_/D vssd1 vssd1 vccd1 vccd1 _8169_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3248_ _6619_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3248_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7368__4 _7369__5/A vssd1 vssd1 vccd1 vccd1 _8306_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6873__442 _6873__442/A vssd1 vssd1 vccd1 vccd1 _8037_/CLK sky130_fd_sc_hd__inv_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6921__476 _6922__477/A vssd1 vssd1 vccd1 vccd1 _8073_/CLK sky130_fd_sc_hd__inv_2
X_5870_ _5870_/A vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4821_ _8265_/Q _4719_/Y _4720_/X _8241_/Q _4556_/A vssd1 vssd1 vccd1 vccd1 _4821_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8434__209 vssd1 vssd1 vccd1 vccd1 _8434__209/HI manufacturerID[1] sky130_fd_sc_hd__conb_1
X_7540_ _7540_/A _7540_/B vssd1 vssd1 vccd1 vccd1 _7549_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _8207_/Q _4703_/A _8024_/Q _4705_/A _4622_/A vssd1 vssd1 vccd1 vccd1 _4752_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7471_ _7488_/A vssd1 vssd1 vccd1 vccd1 _7482_/A sky130_fd_sc_hd__clkbuf_2
X_4683_ _4683_/A _4704_/A vssd1 vssd1 vccd1 vccd1 _4729_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6422_ _6422_/A vssd1 vssd1 vccd1 vccd1 _6422_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3203_ clkbuf_0__3203_/X vssd1 vssd1 vccd1 vccd1 _6495__270/A sky130_fd_sc_hd__clkbuf_4
X_6353_ _6353_/A vssd1 vssd1 vccd1 vccd1 _7732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6284_ _8401_/Q vssd1 vssd1 vccd1 vccd1 _6719_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5304_ _5567_/A vssd1 vssd1 vccd1 vccd1 _5304_/X sky130_fd_sc_hd__buf_2
X_8023_ _8023_/CLK _8023_/D vssd1 vssd1 vccd1 vccd1 _8023_/Q sky130_fd_sc_hd__dfxtp_1
X_5235_ _8366_/Q _5114_/X _5108_/B _8374_/Q _5009_/A vssd1 vssd1 vccd1 vccd1 _5235_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5166_ _8368_/Q _5114_/X _5183_/A _8376_/Q _5009_/A vssd1 vssd1 vccd1 vccd1 _5166_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4117_ _4117_/A vssd1 vssd1 vccd1 vccd1 _8258_/D sky130_fd_sc_hd__clkbuf_1
X_5097_ _5113_/A vssd1 vssd1 vccd1 vccd1 _5150_/A sky130_fd_sc_hd__inv_2
XFILLER_83_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4048_ _4387_/B _4413_/A _4414_/A vssd1 vssd1 vccd1 vccd1 _5599_/A sky130_fd_sc_hd__or3b_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _7720_/Q input33/X _6008_/S vssd1 vssd1 vccd1 vccd1 _5999_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7807_ _7807_/CLK _7807_/D vssd1 vssd1 vccd1 vccd1 _7807_/Q sky130_fd_sc_hd__dfxtp_1
X_7738_ _8066_/CLK _7738_/D vssd1 vssd1 vccd1 vccd1 _7738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7669_ _7992_/CLK _7669_/D vssd1 vssd1 vccd1 vccd1 _7669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7080__104 _7080__104/A vssd1 vssd1 vccd1 vccd1 _8201_/CLK sky130_fd_sc_hd__inv_2
X_6962__510 _6962__510/A vssd1 vssd1 vccd1 vccd1 _8107_/CLK sky130_fd_sc_hd__inv_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _7997_/Q _5020_/B vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6661__359 _6661__359/A vssd1 vssd1 vccd1 vccd1 _7940_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5922_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5931_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5853_ _7614_/B _5855_/B vssd1 vssd1 vccd1 vccd1 _5854_/A sky130_fd_sc_hd__or2_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5784_ _5784_/A vssd1 vssd1 vccd1 vccd1 _7658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4804_ _4863_/B _4782_/X _4789_/X _4803_/X vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__a31o_2
X_7523_ _8355_/Q _7523_/B _7513_/X vssd1 vssd1 vccd1 vccd1 _7523_/X sky130_fd_sc_hd__or3b_1
X_4735_ _4696_/A _7964_/Q _7768_/Q _4698_/A vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3582_ _7289_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3582_/X sky130_fd_sc_hd__clkbuf_16
X_7454_ _7454_/A vssd1 vssd1 vccd1 vccd1 _8332_/D sky130_fd_sc_hd__clkbuf_1
X_4666_ _4650_/S _4665_/X _4770_/A vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4597_ _7652_/Q _7660_/Q _7711_/Q _7812_/Q _4595_/X _4596_/X vssd1 vssd1 vccd1 vccd1
+ _4597_/X sky130_fd_sc_hd__mux4_2
X_6405_ _6404_/X _6405_/B vssd1 vssd1 vccd1 vccd1 _6406_/A sky130_fd_sc_hd__and2b_1
X_6336_ _8390_/Q vssd1 vssd1 vccd1 vccd1 _7170_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6412__202 _6413__203/A vssd1 vssd1 vccd1 vccd1 _7759_/CLK sky130_fd_sc_hd__inv_2
X_6267_ _7135_/A _6249_/A _6301_/B _6289_/A vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6198_ _7220_/A vssd1 vssd1 vccd1 vccd1 _6198_/X sky130_fd_sc_hd__clkbuf_2
X_8006_ _8006_/CLK _8006_/D vssd1 vssd1 vccd1 vccd1 _8006_/Q sky130_fd_sc_hd__dfxtp_1
X_5218_ _5218_/A _5218_/B vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__or2_1
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5149_ _8323_/Q _8069_/Q _5149_/S vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3195_ clkbuf_0__3195_/X vssd1 vssd1 vccd1 vccd1 _6451__234/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4520_ _8361_/Q vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4451_ _4451_/A vssd1 vssd1 vccd1 vccd1 _8099_/D sky130_fd_sc_hd__clkbuf_1
X_7170_ _7170_/A _7220_/A vssd1 vssd1 vccd1 vccd1 _7265_/B sky130_fd_sc_hd__nand2_1
X_6886__452 _6888__454/A vssd1 vssd1 vccd1 vccd1 _8047_/CLK sky130_fd_sc_hd__inv_2
X_6121_ _6119_/X _7698_/Q _6116_/X _6120_/X _7666_/Q vssd1 vssd1 vccd1 vccd1 _7666_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _4223_/X _8124_/Q _4384_/S vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6052_ _6052_/A vssd1 vssd1 vccd1 vccd1 _6062_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5003_/A vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__buf_2
XFILLER_39_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _5905_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5906_/A sky130_fd_sc_hd__and2_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5836_ _6687_/B _5844_/B vssd1 vssd1 vccd1 vccd1 _5837_/A sky130_fd_sc_hd__or2_1
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3597_ clkbuf_0__3597_/X vssd1 vssd1 vccd1 vccd1 _7369__5/A sky130_fd_sc_hd__clkbuf_4
X_5767_ _5555_/X _7709_/Q _5771_/S vssd1 vssd1 vccd1 vccd1 _5768_/A sky130_fd_sc_hd__mux2_1
X_7506_ _7506_/A _7506_/B vssd1 vssd1 vccd1 vccd1 _7506_/X sky130_fd_sc_hd__or2_1
X_5698_ _5698_/A vssd1 vssd1 vccd1 vccd1 _7785_/D sky130_fd_sc_hd__clkbuf_1
X_4718_ _8142_/Q _4716_/X _4717_/X _7824_/Q vssd1 vssd1 vccd1 vccd1 _4718_/X sky130_fd_sc_hd__a22o_1
X_7437_ _7489_/A _7496_/B _7439_/C vssd1 vssd1 vccd1 vccd1 _7474_/A sky130_fd_sc_hd__o21a_1
X_4649_ _8027_/Q _7982_/Q _7842_/Q _8210_/Q _4596_/A _4595_/X vssd1 vssd1 vccd1 vccd1
+ _4649_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6319_ _7723_/Q _6265_/X _6307_/X _6318_/X vssd1 vssd1 vccd1 vccd1 _7723_/D sky130_fd_sc_hd__a211o_1
XFILLER_77_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8349_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3247_ clkbuf_0__3247_/X vssd1 vssd1 vccd1 vccd1 _6618__325/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6419__208 _6421__210/A vssd1 vssd1 vccd1 vccd1 _7765_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _4217_/A vssd1 vssd1 vccd1 vccd1 _3951_/X sky130_fd_sc_hd__clkbuf_2
X_3882_ _3881_/X _8369_/Q _3882_/S vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__mux2_1
X_5621_ _5552_/X _7819_/Q _5627_/S vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3382_ clkbuf_0__3382_/X vssd1 vssd1 vccd1 vccd1 _6938_/A sky130_fd_sc_hd__clkbuf_4
X_5552_ _5552_/A vssd1 vssd1 vccd1 vccd1 _5552_/X sky130_fd_sc_hd__buf_2
X_8340_ _8341_/CLK _8340_/D vssd1 vssd1 vccd1 vccd1 _8340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8271_ _8271_/CLK _8271_/D vssd1 vssd1 vccd1 vccd1 _8271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4503_ _4344_/X _8076_/Q _4505_/S vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__mux2_1
X_5483_ _7897_/Q _4214_/A _5485_/S vssd1 vssd1 vccd1 vccd1 _5484_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7222_ _7222_/A vssd1 vssd1 vccd1 vccd1 _7222_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4434_ _4507_/A _5439_/A vssd1 vssd1 vccd1 vccd1 _4450_/S sky130_fd_sc_hd__or2_2
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7153_ _7593_/A _7153_/B vssd1 vssd1 vccd1 vccd1 _7173_/C sky130_fd_sc_hd__xor2_2
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _8132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7084_ _8401_/Q vssd1 vssd1 vccd1 vccd1 _7096_/A sky130_fd_sc_hd__inv_2
X_6104_ _7600_/A vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__buf_4
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6035_ _6036_/A _7861_/Q _5817_/C _5815_/X _7644_/Q vssd1 vssd1 vccd1 vccd1 _6349_/D
+ sky130_fd_sc_hd__a41o_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4296_/A vssd1 vssd1 vccd1 vccd1 _8159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7986_ _8365_/CLK _7986_/D vssd1 vssd1 vccd1 vccd1 _7986_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5819_ _5955_/A vssd1 vssd1 vccd1 vccd1 _5826_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6799_ _8351_/Q _6910_/A vssd1 vssd1 vccd1 vccd1 _6800_/A sky130_fd_sc_hd__and2_1
XFILLER_10_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6087__178 _6087__178/A vssd1 vssd1 vccd1 vccd1 _7647_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput108 _5957_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput119 _5924_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__buf_2
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ _8248_/Q _4044_/X _4158_/S vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__mux2_1
X_4081_ _7991_/Q vssd1 vssd1 vccd1 vccd1 _4081_/X sky130_fd_sc_hd__buf_2
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7840_ _7840_/CLK _7840_/D vssd1 vssd1 vccd1 vccd1 _7840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7771_ _7771_/CLK _7771_/D vssd1 vssd1 vccd1 vccd1 _7771_/Q sky130_fd_sc_hd__dfxtp_1
X_4983_ _5020_/B _4997_/B vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__or2_2
X_6722_ _7429_/A _7429_/B _8402_/Q vssd1 vssd1 vccd1 vccd1 _6722_/Y sky130_fd_sc_hd__a21oi_1
X_3934_ _4121_/A _3989_/B vssd1 vssd1 vccd1 vccd1 _3964_/S sky130_fd_sc_hd__nor2_2
X_3865_ _5025_/A vssd1 vssd1 vccd1 vccd1 _3865_/X sky130_fd_sc_hd__buf_2
X_5604_ _5604_/A vssd1 vssd1 vccd1 vccd1 _7827_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3365_ clkbuf_0__3365_/X vssd1 vssd1 vccd1 vccd1 _6850__425/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3796_ _7941_/Q vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__buf_2
X_7348__163 _7349__164/A vssd1 vssd1 vccd1 vccd1 _8290_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3402_ _7014_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3402_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5535_ _5288_/X _7874_/Q _5539_/S vssd1 vssd1 vccd1 vccd1 _5536_/A sky130_fd_sc_hd__mux2_1
X_8323_ _8323_/CLK _8323_/D vssd1 vssd1 vccd1 vccd1 _8323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8254_ _8254_/CLK _8254_/D vssd1 vssd1 vccd1 vccd1 _8254_/Q sky130_fd_sc_hd__dfxtp_1
X_5466_ _5466_/A vssd1 vssd1 vccd1 vccd1 _7905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7205_ _7141_/B _7238_/C _7233_/A _7204_/Y vssd1 vssd1 vccd1 vccd1 _7206_/B sky130_fd_sc_hd__o2bb2a_1
X_4417_ _4432_/S vssd1 vssd1 vccd1 vccd1 _4426_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8185_ _8185_/CLK _8185_/D vssd1 vssd1 vccd1 vccd1 _8185_/Q sky130_fd_sc_hd__dfxtp_1
X_5397_ _7935_/Q _4523_/X _5401_/S vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7136_ _7208_/A _7204_/A _7140_/B vssd1 vssd1 vccd1 vccd1 _7207_/A sky130_fd_sc_hd__nand3_1
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3195_ _6447_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3195_/X sky130_fd_sc_hd__clkbuf_16
X_4348_ _4347_/X _8139_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__mux2_1
X_4279_ _4279_/A vssd1 vssd1 vccd1 vccd1 _8166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6018_ _6018_/A vssd1 vssd1 vccd1 vccd1 _6018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _7969_/CLK _7969_/D vssd1 vssd1 vccd1 vccd1 _7969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _5320_/A vssd1 vssd1 vccd1 vccd1 _7973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5251_ _3893_/A _3968_/B _5475_/B _5250_/X _5214_/X vssd1 vssd1 vccd1 vccd1 _8002_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4202_ _8195_/Q _4099_/X _4202_/S vssd1 vssd1 vccd1 vccd1 _4203_/A sky130_fd_sc_hd__mux2_1
X_5182_ _8164_/Q _7902_/Q _5274_/A vssd1 vssd1 vccd1 vccd1 _5182_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4133_ _4133_/A vssd1 vssd1 vccd1 vccd1 _8253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4064_ _8054_/Q _8049_/Q vssd1 vssd1 vccd1 vccd1 _4069_/B sky130_fd_sc_hd__or2b_1
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7823_ _7823_/CLK _7823_/D vssd1 vssd1 vccd1 vccd1 _7823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7754_ _8065_/CLK _7754_/D vssd1 vssd1 vccd1 vccd1 _7754_/Q sky130_fd_sc_hd__dfxtp_1
X_7566__40 _7566__40/A vssd1 vssd1 vccd1 vccd1 _8379_/CLK sky130_fd_sc_hd__inv_2
X_6705_ _8343_/Q _6705_/B vssd1 vssd1 vccd1 vccd1 _6706_/B sky130_fd_sc_hd__xnor2_2
X_4966_ _5100_/B vssd1 vssd1 vccd1 vccd1 _5240_/S sky130_fd_sc_hd__clkbuf_4
X_7685_ _8345_/CLK _7685_/D vssd1 vssd1 vccd1 vccd1 _7685_/Q sky130_fd_sc_hd__dfxtp_1
X_4897_ _4897_/A vssd1 vssd1 vccd1 vccd1 _8037_/D sky130_fd_sc_hd__clkbuf_1
X_3917_ _3932_/S vssd1 vssd1 vccd1 vccd1 _3926_/S sky130_fd_sc_hd__clkbuf_4
X_7030__64 _7031__65/A vssd1 vssd1 vccd1 vccd1 _8161_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3848_ _8381_/Q _3772_/X _3856_/S vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6567_ _6567_/A vssd1 vssd1 vccd1 vccd1 _7866_/D sky130_fd_sc_hd__clkbuf_1
X_3779_ _7993_/Q _7998_/Q vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__and2b_1
X_8306_ _8306_/CLK _8306_/D vssd1 vssd1 vccd1 vccd1 _8306_/Q sky130_fd_sc_hd__dfxtp_1
X_5518_ _5518_/A vssd1 vssd1 vccd1 vccd1 _7882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8237_ _8239_/CLK _8237_/D vssd1 vssd1 vccd1 vccd1 _8237_/Q sky130_fd_sc_hd__dfxtp_1
X_5449_ _3831_/X _7912_/Q _5449_/S vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8168_ _8168_/CLK _8168_/D vssd1 vssd1 vccd1 vccd1 _8168_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3247_ _6613_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3247_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7119_ _7119_/A _7150_/C _7119_/C vssd1 vssd1 vccd1 vccd1 _7234_/A sky130_fd_sc_hd__and3_1
XFILLER_101_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8099_ _8099_/CLK _8099_/D vssd1 vssd1 vccd1 vccd1 _8099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6461__242 _6462__243/A vssd1 vssd1 vccd1 vccd1 _7799_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4820_ _8139_/Q _4697_/A _4699_/A _7821_/Q vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4697_/A _7979_/Q _7839_/Q _4699_/A vssd1 vssd1 vccd1 vccd1 _4751_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7470_ _7470_/A _7470_/B vssd1 vssd1 vccd1 vccd1 _8337_/D sky130_fd_sc_hd__nor2_1
X_4682_ _4682_/A _4682_/B vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__nand2_2
Xclkbuf_1_1_0__3202_ clkbuf_0__3202_/X vssd1 vssd1 vccd1 vccd1 _6487__263/A sky130_fd_sc_hd__clkbuf_4
X_6670__361 _6671__362/A vssd1 vssd1 vccd1 vccd1 _7945_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8410__232 vssd1 vssd1 vccd1 vccd1 partID[2] _8410__232/LO sky130_fd_sc_hd__conb_1
X_6352_ _5909_/A _7732_/Q _6360_/S vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__mux2_1
X_6283_ _7717_/Q _6216_/X _6282_/X vssd1 vssd1 vccd1 vccd1 _7717_/D sky130_fd_sc_hd__a21o_1
X_5303_ _7986_/Q vssd1 vssd1 vccd1 vccd1 _5567_/A sky130_fd_sc_hd__buf_2
XFILLER_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8022_ _8022_/CLK _8022_/D vssd1 vssd1 vccd1 vccd1 _8022_/Q sky130_fd_sc_hd__dfxtp_1
X_5234_ _7877_/Q _7944_/Q _5234_/S vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5165_ _7879_/Q _7946_/Q _5234_/S vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4116_ _8258_/Q _3959_/X _4118_/S vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _7995_/Q vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__clkbuf_2
X_4047_ _8055_/Q vssd1 vssd1 vccd1 vccd1 _4414_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ _7806_/CLK _7806_/D vssd1 vssd1 vccd1 vccd1 _7806_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4949_ _4949_/A _4949_/B _4949_/C _3782_/S vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__or4b_1
X_7737_ _8066_/CLK _7737_/D vssd1 vssd1 vccd1 vccd1 _7737_/Q sky130_fd_sc_hd__dfxtp_1
X_7668_ _7992_/CLK _7668_/D vssd1 vssd1 vccd1 vccd1 _7668_/Q sky130_fd_sc_hd__dfxtp_1
X_6619_ _6650_/A vssd1 vssd1 vccd1 vccd1 _6619_/X sky130_fd_sc_hd__buf_1
XFILLER_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7599_ _7599_/A _7599_/B vssd1 vssd1 vccd1 vccd1 _7599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7560__35 _7560__35/A vssd1 vssd1 vccd1 vccd1 _8374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6468__248 _6470__250/A vssd1 vssd1 vccd1 vccd1 _7805_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5921_ _5921_/A vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7379__13 _7379__13/A vssd1 vssd1 vccd1 vccd1 _8315_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5852_ _5852_/A vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__clkbuf_1
X_5783_ _7658_/Q _5555_/A _5785_/S vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__mux2_1
X_4803_ _4757_/A _4792_/X _4795_/X _4802_/X _4549_/A vssd1 vssd1 vccd1 vccd1 _4803_/X
+ sky130_fd_sc_hd__o311a_1
X_7522_ _8353_/Q _7511_/X _7521_/X _7519_/X vssd1 vssd1 vccd1 vccd1 _8353_/D sky130_fd_sc_hd__o211a_1
X_4734_ _4729_/X _4732_/X _4733_/X vssd1 vssd1 vccd1 vccd1 _4738_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7453_ _7493_/A _7453_/B vssd1 vssd1 vccd1 vccd1 _7454_/A sky130_fd_sc_hd__and2_1
X_4665_ _7649_/Q _7657_/Q _7708_/Q _7809_/Q _4571_/A _4596_/X vssd1 vssd1 vccd1 vccd1
+ _4665_/X sky130_fd_sc_hd__mux4_1
X_4596_ _4596_/A vssd1 vssd1 vccd1 vccd1 _4596_/X sky130_fd_sc_hd__clkbuf_4
X_6404_ _6400_/A _6185_/C _6342_/A _6403_/B vssd1 vssd1 vccd1 vccd1 _6404_/X sky130_fd_sc_hd__a31o_1
X_6335_ _7728_/Q _6320_/X _6324_/X _6334_/X vssd1 vssd1 vccd1 vccd1 _7728_/D sky130_fd_sc_hd__a211o_1
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6266_ _8404_/Q vssd1 vssd1 vccd1 vccd1 _7135_/A sky130_fd_sc_hd__buf_2
X_8005_ _8005_/CLK _8005_/D vssd1 vssd1 vccd1 vccd1 _8005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6197_ _8204_/Q _8203_/Q vssd1 vssd1 vccd1 vccd1 _7220_/A sky130_fd_sc_hd__nor2_2
XFILLER_28_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5217_ _8289_/Q _8297_/Q _5227_/S vssd1 vssd1 vccd1 vccd1 _5218_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3401_ clkbuf_0__3401_/X vssd1 vssd1 vccd1 vccd1 _7026_/A sky130_fd_sc_hd__clkbuf_4
X_5148_ _5148_/A vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__buf_2
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5079_ _7937_/Q _7929_/Q _7921_/Q _7956_/Q _4978_/X _4995_/X vssd1 vssd1 vccd1 vccd1
+ _5079_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3194_ clkbuf_0__3194_/X vssd1 vssd1 vccd1 vccd1 _6443__227/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6677__367 _6677__367/A vssd1 vssd1 vccd1 vccd1 _7951_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2978_ clkbuf_0__2978_/X vssd1 vssd1 vccd1 vccd1 _6208__195/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6474__252 _6474__252/A vssd1 vssd1 vccd1 vccd1 _7809_/CLK sky130_fd_sc_hd__inv_2
X_4450_ _4226_/X _8099_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7342__158 _7344__160/A vssd1 vssd1 vccd1 vccd1 _8285_/CLK sky130_fd_sc_hd__inv_2
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _8125_/D sky130_fd_sc_hd__clkbuf_1
X_6120_ _6129_/A vssd1 vssd1 vccd1 vccd1 _6120_/X sky130_fd_sc_hd__clkbuf_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6051_/A vssd1 vssd1 vccd1 vccd1 _6051_/X sky130_fd_sc_hd__buf_2
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A vssd1 vssd1 vccd1 vccd1 _5002_/X sky130_fd_sc_hd__buf_2
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5904_ _5904_/A vssd1 vssd1 vccd1 vccd1 _5904_/X sky130_fd_sc_hd__clkbuf_1
X_6884_ _6896_/A vssd1 vssd1 vccd1 vccd1 _6884_/X sky130_fd_sc_hd__buf_1
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5835_ _5903_/B vssd1 vssd1 vccd1 vccd1 _5844_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1_0__3596_ clkbuf_0__3596_/X vssd1 vssd1 vccd1 vccd1 _7382_/A sky130_fd_sc_hd__clkbuf_4
X_5766_ _5766_/A vssd1 vssd1 vccd1 vccd1 _7710_/D sky130_fd_sc_hd__clkbuf_1
X_6637__340 _6637__340/A vssd1 vssd1 vccd1 vccd1 _7921_/CLK sky130_fd_sc_hd__inv_2
X_6934__487 _6936__489/A vssd1 vssd1 vccd1 vccd1 _8084_/CLK sky130_fd_sc_hd__inv_2
X_7505_ _8348_/Q _7498_/A _8349_/Q vssd1 vssd1 vccd1 vccd1 _7506_/B sky130_fd_sc_hd__a21oi_1
X_5697_ _7785_/Q _5584_/X _5699_/S vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__mux2_1
X_4717_ _4717_/A vssd1 vssd1 vccd1 vccd1 _4717_/X sky130_fd_sc_hd__buf_2
X_4648_ _8120_/Q _7890_/Q _7834_/Q _7794_/Q _4579_/A _4589_/X vssd1 vssd1 vccd1 vccd1
+ _4648_/X sky130_fd_sc_hd__mux4_1
X_7436_ _7414_/X _7419_/X _7435_/X _7401_/B _8330_/Q vssd1 vssd1 vccd1 vccd1 _7439_/C
+ sky130_fd_sc_hd__a311o_2
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579_ _4579_/A vssd1 vssd1 vccd1 vccd1 _4579_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6318_ _8396_/Q _6326_/B _6322_/C _6326_/D vssd1 vssd1 vccd1 vccd1 _6318_/X sky130_fd_sc_hd__and4_1
XFILLER_39_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6249_ _6249_/A vssd1 vssd1 vccd1 vccd1 _6249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3246_ clkbuf_0__3246_/X vssd1 vssd1 vccd1 vccd1 _6611__319/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3950_ _8361_/Q vssd1 vssd1 vccd1 vccd1 _4217_/A sky130_fd_sc_hd__buf_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3881_ _8361_/Q vssd1 vssd1 vccd1 vccd1 _3881_/X sky130_fd_sc_hd__buf_2
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5620_ _5620_/A vssd1 vssd1 vccd1 vccd1 _7820_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3381_ clkbuf_0__3381_/X vssd1 vssd1 vccd1 vccd1 _6914__471/A sky130_fd_sc_hd__clkbuf_4
X_5551_ _5551_/A vssd1 vssd1 vccd1 vccd1 _7844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8270_ _8270_/CLK _8270_/D vssd1 vssd1 vccd1 vccd1 _8270_/Q sky130_fd_sc_hd__dfxtp_1
X_4502_ _4502_/A vssd1 vssd1 vccd1 vccd1 _8077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7221_ _7221_/A _7221_/B vssd1 vssd1 vccd1 vccd1 _7221_/Y sky130_fd_sc_hd__nand2_1
X_5482_ _5482_/A vssd1 vssd1 vccd1 vccd1 _7898_/D sky130_fd_sc_hd__clkbuf_1
X_4433_ _4433_/A vssd1 vssd1 vccd1 vccd1 _8107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7152_ _7152_/A _7247_/A vssd1 vssd1 vccd1 vccd1 _7153_/B sky130_fd_sc_hd__xnor2_2
X_4364_ _8132_/Q _4140_/X _4366_/S vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7083_ _8231_/Q _8230_/Q _8229_/Q _8204_/Q vssd1 vssd1 vccd1 vccd1 _7252_/B sky130_fd_sc_hd__and4_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _4214_/X _8159_/Q _4297_/S vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6034_ _6034_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6034_/X sky130_fd_sc_hd__and2_1
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7985_ _8365_/CLK _7985_/D vssd1 vssd1 vccd1 vccd1 _7985_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5818_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__inv_2
X_6798_ _6798_/A vssd1 vssd1 vccd1 vccd1 _7985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5749_ _7762_/Q _5555_/A _5753_/S vssd1 vssd1 vccd1 vccd1 _5750_/A sky130_fd_sc_hd__mux2_1
X_7419_ _7415_/Y _7416_/X _7417_/X _7418_/X _7491_/A vssd1 vssd1 vccd1 vccd1 _7419_/X
+ sky130_fd_sc_hd__o2111a_1
X_8399_ _8399_/CLK _8399_/D vssd1 vssd1 vccd1 vccd1 _8399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6425__213 _6427__215/A vssd1 vssd1 vccd1 vccd1 _7770_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput109 _5959_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__buf_2
XFILLER_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ _4080_/A vssd1 vssd1 vccd1 vccd1 _8272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7770_ _7770_/CLK _7770_/D vssd1 vssd1 vccd1 vccd1 _7770_/Q sky130_fd_sc_hd__dfxtp_1
X_4982_ _7996_/Q _4982_/B vssd1 vssd1 vccd1 vccd1 _4997_/B sky130_fd_sc_hd__nor2_1
X_6777__383 _6777__383/A vssd1 vssd1 vccd1 vccd1 _7968_/CLK sky130_fd_sc_hd__inv_2
X_6721_ _8335_/Q _6738_/B _8336_/Q vssd1 vssd1 vccd1 vccd1 _7429_/B sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8066_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3933_ _3933_/A vssd1 vssd1 vccd1 vccd1 _8313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3864_ _8365_/Q vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__buf_4
X_5603_ _5552_/X _7827_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3795_ _5261_/A _5261_/B vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__nand2_1
X_8322_ _8322_/CLK _8322_/D vssd1 vssd1 vccd1 vccd1 _8322_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3401_ _7013_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3401_/X sky130_fd_sc_hd__clkbuf_16
X_5534_ _5534_/A vssd1 vssd1 vccd1 vccd1 _7875_/D sky130_fd_sc_hd__clkbuf_1
X_8253_ _8253_/CLK _8253_/D vssd1 vssd1 vccd1 vccd1 _8253_/Q sky130_fd_sc_hd__dfxtp_1
X_5465_ _7905_/Q _4214_/A _5467_/S vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__mux2_1
X_7204_ _7204_/A vssd1 vssd1 vccd1 vccd1 _7204_/Y sky130_fd_sc_hd__clkinv_2
X_8184_ _8184_/CLK _8184_/D vssd1 vssd1 vccd1 vccd1 _8184_/Q sky130_fd_sc_hd__dfxtp_1
X_4416_ _5635_/A _4875_/A vssd1 vssd1 vccd1 vccd1 _4432_/S sky130_fd_sc_hd__nor2_2
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7135_ _7135_/A _7135_/B vssd1 vssd1 vccd1 vccd1 _7135_/X sky130_fd_sc_hd__xor2_1
X_5396_ _5396_/A vssd1 vssd1 vccd1 vccd1 _7936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3194_ _6441_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3194_/X sky130_fd_sc_hd__clkbuf_16
X_4347_ _7985_/Q vssd1 vssd1 vccd1 vccd1 _4347_/X sky130_fd_sc_hd__buf_2
XFILLER_101_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4278_ _8166_/Q _4134_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__mux2_1
X_6017_ _7674_/Q _6016_/X _6023_/S vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__mux2_4
XFILLER_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7003__543 _7004__544/A vssd1 vssd1 vccd1 vccd1 _8140_/CLK sky130_fd_sc_hd__inv_2
X_6899__463 _6901__465/A vssd1 vssd1 vccd1 vccd1 _8058_/CLK sky130_fd_sc_hd__inv_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7968_ _7968_/CLK _7968_/D vssd1 vssd1 vccd1 vccd1 _7968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2978_ _6102_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2978_/X sky130_fd_sc_hd__clkbuf_16
X_7899_ _7899_/CLK _7899_/D vssd1 vssd1 vccd1 vccd1 _7899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6919_ _6981_/A vssd1 vssd1 vccd1 vccd1 _6919_/X sky130_fd_sc_hd__buf_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6574__290 _6574__290/A vssd1 vssd1 vccd1 vccd1 _7871_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6093__183 _6093__183/A vssd1 vssd1 vccd1 vccd1 _7652_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _5347_/C _5250_/B vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__or2_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4201_ _4201_/A vssd1 vssd1 vccd1 vccd1 _8196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5181_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _8253_/Q _4131_/X _4135_/S vssd1 vssd1 vccd1 vccd1 _4133_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4063_ _4063_/A vssd1 vssd1 vccd1 vccd1 _4853_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7822_ _7822_/CLK _7822_/D vssd1 vssd1 vccd1 vccd1 _7822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7753_ _8349_/CLK _7753_/D vssd1 vssd1 vccd1 vccd1 _7753_/Q sky130_fd_sc_hd__dfxtp_1
X_4965_ _4965_/A vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__buf_2
X_7015__51 _7016__52/A vssd1 vssd1 vccd1 vccd1 _8148_/CLK sky130_fd_sc_hd__inv_2
X_6704_ _7612_/A _6704_/B vssd1 vssd1 vccd1 vccd1 _6743_/B sky130_fd_sc_hd__xor2_1
X_3916_ _5348_/A _3989_/B vssd1 vssd1 vccd1 vccd1 _3932_/S sky130_fd_sc_hd__or2_2
X_7684_ _8349_/CLK _7684_/D vssd1 vssd1 vccd1 vccd1 _7684_/Q sky130_fd_sc_hd__dfxtp_1
X_4896_ _8037_/Q _4386_/X _4904_/S vssd1 vssd1 vccd1 vccd1 _4897_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3847_ _3862_/S vssd1 vssd1 vccd1 vccd1 _3856_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6566_ _7866_/Q _5899_/A _6570_/S vssd1 vssd1 vccd1 vccd1 _6567_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3347_ clkbuf_0__3347_/X vssd1 vssd1 vccd1 vccd1 _6814__400/A sky130_fd_sc_hd__clkbuf_4
X_3778_ _7998_/Q vssd1 vssd1 vccd1 vccd1 _5261_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8305_ _8305_/CLK _8305_/D vssd1 vssd1 vccd1 vccd1 _8305_/Q sky130_fd_sc_hd__dfxtp_1
X_5517_ _7882_/Q _4211_/A _5521_/S vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8236_ _8239_/CLK _8236_/D vssd1 vssd1 vccd1 vccd1 _8236_/Q sky130_fd_sc_hd__dfxtp_1
X_5448_ _5448_/A vssd1 vssd1 vccd1 vccd1 _7913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8167_ _8167_/CLK _8167_/D vssd1 vssd1 vccd1 vccd1 _8167_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3246_ _6607_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3246_/X sky130_fd_sc_hd__clkbuf_16
X_5379_ _7946_/Q _4523_/X _5383_/S vssd1 vssd1 vccd1 vccd1 _5380_/A sky130_fd_sc_hd__mux2_1
X_7118_ _7238_/A _7238_/B _7117_/A vssd1 vssd1 vccd1 vccd1 _7118_/Y sky130_fd_sc_hd__a21oi_1
X_8098_ _8098_/CLK _8098_/D vssd1 vssd1 vccd1 vccd1 _8098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6205__192 _6208__195/A vssd1 vssd1 vccd1 vccd1 _7704_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6101__190 _6101__190/A vssd1 vssd1 vccd1 vccd1 _7659_/CLK sky130_fd_sc_hd__inv_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7297__122 _7300__125/A vssd1 vssd1 vccd1 vccd1 _8249_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6880__448 _6882__450/A vssd1 vssd1 vccd1 vccd1 _8043_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4750_/A vssd1 vssd1 vccd1 vccd1 _4750_/X sky130_fd_sc_hd__clkbuf_2
X_4681_ _4681_/A vssd1 vssd1 vccd1 vccd1 _4681_/X sky130_fd_sc_hd__buf_4
Xclkbuf_1_1_0__3201_ clkbuf_0__3201_/X vssd1 vssd1 vccd1 vccd1 _6483__260/A sky130_fd_sc_hd__clkbuf_4
X_6351_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6360_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_115_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7306__129 _7306__129/A vssd1 vssd1 vccd1 vccd1 _8256_/CLK sky130_fd_sc_hd__inv_2
X_6631__335 _6631__335/A vssd1 vssd1 vccd1 vccd1 _7916_/CLK sky130_fd_sc_hd__inv_2
X_5302_ _5302_/A vssd1 vssd1 vccd1 vccd1 _7979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6282_ _6270_/A _6278_/X _6280_/X _7642_/A vssd1 vssd1 vccd1 vccd1 _6282_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8021_ _8021_/CLK _8021_/D vssd1 vssd1 vccd1 vccd1 _8021_/Q sky130_fd_sc_hd__dfxtp_1
X_5233_ _5148_/X _5231_/X _5232_/X _5045_/A vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__o211a_1
X_5164_ _5148_/X _5162_/X _5163_/X _5045_/A vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__o211a_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4115_ _4115_/A vssd1 vssd1 vccd1 vccd1 _8259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5095_ _5095_/A vssd1 vssd1 vccd1 vccd1 _5265_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4046_ _8053_/Q vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7805_ _7805_/CLK _7805_/D vssd1 vssd1 vccd1 vccd1 _7805_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _7668_/Q _5996_/X _6006_/S vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__mux2_4
X_7736_ _8066_/CLK _7736_/D vssd1 vssd1 vccd1 vccd1 _7736_/Q sky130_fd_sc_hd__dfxtp_1
X_4948_ _4948_/A vssd1 vssd1 vccd1 vccd1 _8014_/D sky130_fd_sc_hd__clkbuf_1
X_7667_ _7846_/CLK _7667_/D vssd1 vssd1 vccd1 vccd1 _7667_/Q sky130_fd_sc_hd__dfxtp_1
X_4879_ _8044_/Q _4392_/X _4885_/S vssd1 vssd1 vccd1 vccd1 _4880_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7598_ _7614_/A _7598_/B vssd1 vssd1 vccd1 vccd1 _7598_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6549_ _6549_/A vssd1 vssd1 vccd1 vccd1 _7858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8219_ _8231_/CLK _8219_/D vssd1 vssd1 vccd1 vccd1 _8219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7184__108 _7184__108/A vssd1 vssd1 vccd1 vccd1 _8207_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8440__215 vssd1 vssd1 vccd1 vccd1 _8440__215/HI manufacturerID[7] sky130_fd_sc_hd__conb_1
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _5920_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__and2_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5851_ _7617_/A _5855_/B vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__or2_1
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5782_ _5782_/A vssd1 vssd1 vccd1 vccd1 _7659_/D sky130_fd_sc_hd__clkbuf_1
X_6817__401 _6820__404/A vssd1 vssd1 vccd1 vccd1 _7994_/CLK sky130_fd_sc_hd__inv_2
X_4802_ _4802_/A _4802_/B _4802_/C vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__or3_1
X_7521_ _8354_/Q _7523_/B _7513_/X vssd1 vssd1 vccd1 vccd1 _7521_/X sky130_fd_sc_hd__or3b_1
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4733_ _4703_/A _7760_/Q _4725_/A _8017_/Q _4726_/A vssd1 vssd1 vccd1 vccd1 _4733_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7452_ _7421_/A _7466_/A _7446_/Y _7422_/B vssd1 vssd1 vccd1 vccd1 _7453_/B sky130_fd_sc_hd__a22o_1
X_6403_ _6403_/A _6403_/B vssd1 vssd1 vccd1 vccd1 _7754_/D sky130_fd_sc_hd__nor2_1
X_4664_ _4664_/A _4664_/B vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__and2_1
X_4595_ _4595_/A vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__buf_2
X_6334_ _8391_/Q _6337_/B _7943_/Q _6337_/D vssd1 vssd1 vccd1 vccd1 _6334_/X sky130_fd_sc_hd__and4_1
X_6265_ _6320_/A vssd1 vssd1 vccd1 vccd1 _6265_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8004_ _8004_/CLK _8004_/D vssd1 vssd1 vccd1 vccd1 _8004_/Q sky130_fd_sc_hd__dfxtp_1
X_5216_ _5212_/Y _5213_/Y _5215_/Y vssd1 vssd1 vccd1 vccd1 _8005_/D sky130_fd_sc_hd__a21oi_1
X_6196_ _8231_/Q _6192_/X _6194_/X _7262_/C vssd1 vssd1 vccd1 vccd1 _6196_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0_0__3400_ clkbuf_0__3400_/X vssd1 vssd1 vccd1 vccd1 _7075_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5147_ _5103_/X _5145_/X _5146_/X vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__o21a_1
X_5078_ _4988_/X _5075_/X _5077_/X vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4029_ _4029_/A vssd1 vssd1 vccd1 vccd1 _8280_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3262_ clkbuf_0__3262_/X vssd1 vssd1 vccd1 vccd1 _6686__375/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0_0__3193_ clkbuf_0__3193_/X vssd1 vssd1 vccd1 vccd1 _6453_/A sky130_fd_sc_hd__clkbuf_4
X_8417__239 vssd1 vssd1 vccd1 vccd1 partID[15] _8417__239/LO sky130_fd_sc_hd__conb_1
XFILLER_100_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7719_ _7989_/CLK _7719_/D vssd1 vssd1 vccd1 vccd1 _7719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2977_ clkbuf_0__2977_/X vssd1 vssd1 vccd1 vccd1 _6098__187/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6771__378 _6772__379/A vssd1 vssd1 vccd1 vccd1 _7963_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4380_ _4220_/X _8125_/Q _4384_/S vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6050_ _7683_/Q _6048_/X _6039_/X _6049_/X vssd1 vssd1 vccd1 vccd1 _6050_/X sky130_fd_sc_hd__o22a_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5001_ _7997_/Q _5020_/B vssd1 vssd1 vccd1 vccd1 _5002_/A sky130_fd_sc_hd__xor2_2
XFILLER_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7049__79 _7050__80/A vssd1 vssd1 vccd1 vccd1 _8176_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5903_ _5903_/A _5903_/B vssd1 vssd1 vccd1 vccd1 _5904_/A sky130_fd_sc_hd__or2_1
X_6883_ _6883_/A vssd1 vssd1 vccd1 vccd1 _6883_/X sky130_fd_sc_hd__buf_1
X_5834_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5903_/B sky130_fd_sc_hd__clkbuf_4
X_6893__458 _6893__458/A vssd1 vssd1 vccd1 vccd1 _8053_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3595_ clkbuf_0__3595_/X vssd1 vssd1 vccd1 vccd1 _7359__172/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5765_ _5552_/X _7710_/Q _5771_/S vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__mux2_1
X_7504_ _8348_/Q _7497_/Y _7503_/X _7448_/X vssd1 vssd1 vccd1 vccd1 _8348_/D sky130_fd_sc_hd__o211a_1
X_5696_ _5696_/A vssd1 vssd1 vccd1 vccd1 _7786_/D sky130_fd_sc_hd__clkbuf_1
X_4716_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4716_/X sky130_fd_sc_hd__clkbuf_2
X_7435_ _7435_/A _7435_/B _7435_/C _7435_/D vssd1 vssd1 vccd1 vccd1 _7435_/X sky130_fd_sc_hd__and4_1
X_4647_ _4650_/S _4645_/X _4770_/A vssd1 vssd1 vccd1 vccd1 _4647_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4578_ _4682_/B vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__buf_2
X_6317_ _7722_/Q _6265_/X _6307_/X _6316_/X vssd1 vssd1 vccd1 vccd1 _7722_/D sky130_fd_sc_hd__a211o_1
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6248_ _7712_/Q _6216_/X _6247_/X vssd1 vssd1 vccd1 vccd1 _7712_/D sky130_fd_sc_hd__a21o_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6179_ _6179_/A vssd1 vssd1 vccd1 vccd1 _7699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6683__372 _6683__372/A vssd1 vssd1 vccd1 vccd1 _7956_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3245_ clkbuf_0__3245_/X vssd1 vssd1 vccd1 vccd1 _6606__315/A sky130_fd_sc_hd__clkbuf_4
XFILLER_111_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8223_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3880_ _3880_/A vssd1 vssd1 vccd1 vccd1 _8370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _5547_/X _7844_/Q _5562_/S vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5481_ _7898_/Q _4211_/A _5485_/S vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__mux2_1
X_4501_ _4341_/X _8077_/Q _4505_/S vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__mux2_1
X_7220_ _7220_/A vssd1 vssd1 vccd1 vccd1 _7220_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4432_ _8107_/Q _4410_/X _4432_/S vssd1 vssd1 vccd1 vccd1 _4433_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7151_ _7151_/A _7151_/B _7166_/A vssd1 vssd1 vccd1 vccd1 _7247_/A sky130_fd_sc_hd__or3b_2
X_4363_ _4363_/A vssd1 vssd1 vccd1 vccd1 _8133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8446__221 vssd1 vssd1 vccd1 vccd1 _8446__221/HI partID[5] sky130_fd_sc_hd__conb_1
X_7082_ _3814_/X _7533_/B _6287_/X _6118_/A vssd1 vssd1 vccd1 vccd1 _7285_/S sky130_fd_sc_hd__a31oi_4
XFILLER_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _4294_/A vssd1 vssd1 vccd1 vccd1 _8160_/D sky130_fd_sc_hd__clkbuf_1
X_6102_ _6209_/A vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__buf_1
XFILLER_113_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6033_ _6052_/A vssd1 vssd1 vccd1 vccd1 _6070_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7984_ _7984_/CLK _7984_/D vssd1 vssd1 vccd1 vccd1 _7984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6940__492 _6941__493/A vssd1 vssd1 vccd1 vccd1 _8089_/CLK sky130_fd_sc_hd__inv_2
X_6901__465 _6901__465/A vssd1 vssd1 vccd1 vccd1 _8060_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5817_ _6349_/A _6687_/A _5817_/C _5966_/A vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__nand4_4
X_6797_ _8350_/Q _6910_/A vssd1 vssd1 vccd1 vccd1 _6798_/A sky130_fd_sc_hd__and2_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5748_ _5748_/A vssd1 vssd1 vccd1 vccd1 _7763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5679_ _7793_/Q _5584_/X _5681_/S vssd1 vssd1 vccd1 vccd1 _5680_/A sky130_fd_sc_hd__mux2_1
X_7418_ _8396_/Q _7418_/B vssd1 vssd1 vccd1 vccd1 _7418_/X sky130_fd_sc_hd__xor2_1
X_8398_ _8407_/CLK _8398_/D vssd1 vssd1 vccd1 vccd1 _8398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7291__117 _7291__117/A vssd1 vssd1 vccd1 vccd1 _8244_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput92 _7703_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__buf_2
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7578__50 _7578__50/A vssd1 vssd1 vccd1 vccd1 _8389_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _4981_/A vssd1 vssd1 vccd1 vccd1 _5020_/B sky130_fd_sc_hd__buf_2
X_6720_ _6738_/B _6720_/B vssd1 vssd1 vccd1 vccd1 _7429_/A sky130_fd_sc_hd__nand2_1
X_3932_ _3890_/X _8313_/Q _3932_/S vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7042__74 _7043__75/A vssd1 vssd1 vccd1 vccd1 _8171_/CLK sky130_fd_sc_hd__inv_2
X_3863_ _3863_/A vssd1 vssd1 vccd1 vccd1 _8374_/D sky130_fd_sc_hd__clkbuf_1
X_6651_ _6681_/A vssd1 vssd1 vccd1 vccd1 _6651_/X sky130_fd_sc_hd__buf_1
XFILLER_32_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5602_ _5602_/A vssd1 vssd1 vccd1 vccd1 _7828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5533_ _5284_/X _7875_/Q _5539_/S vssd1 vssd1 vccd1 vccd1 _5534_/A sky130_fd_sc_hd__mux2_1
X_3794_ _6340_/B _8012_/Q vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__and2b_1
Xclkbuf_0__3400_ _7012_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3400_/X sky130_fd_sc_hd__clkbuf_16
X_8321_ _8321_/CLK _8321_/D vssd1 vssd1 vccd1 vccd1 _8321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5464_ _5464_/A vssd1 vssd1 vccd1 vccd1 _7906_/D sky130_fd_sc_hd__clkbuf_1
X_8252_ _8252_/CLK _8252_/D vssd1 vssd1 vccd1 vccd1 _8252_/Q sky130_fd_sc_hd__dfxtp_1
X_7203_ _7237_/B vssd1 vssd1 vccd1 vccd1 _7233_/A sky130_fd_sc_hd__clkbuf_2
X_4415_ _4387_/B _4930_/C _4930_/A vssd1 vssd1 vccd1 vccd1 _4875_/A sky130_fd_sc_hd__nand3b_2
Xclkbuf_0__3262_ _6681_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3262_/X sky130_fd_sc_hd__clkbuf_16
X_8183_ _8183_/CLK _8183_/D vssd1 vssd1 vccd1 vccd1 _8183_/Q sky130_fd_sc_hd__dfxtp_1
X_5395_ _7936_/Q _4520_/X _5395_/S vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7134_ _7134_/A _7134_/B vssd1 vssd1 vccd1 vccd1 _7135_/B sky130_fd_sc_hd__nand2_1
X_4346_ _4346_/A vssd1 vssd1 vccd1 vccd1 _8140_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3193_ _6440_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3193_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6487__263 _6487__263/A vssd1 vssd1 vccd1 vccd1 _7820_/CLK sky130_fd_sc_hd__inv_2
X_4277_ _4277_/A vssd1 vssd1 vccd1 vccd1 _8167_/D sky130_fd_sc_hd__clkbuf_1
X_6016_ _7725_/Q input7/X _6025_/S vssd1 vssd1 vccd1 vccd1 _6016_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7355__169 _7355__169/A vssd1 vssd1 vccd1 vccd1 _8296_/CLK sky130_fd_sc_hd__inv_2
X_7967_ _7967_/CLK _7967_/D vssd1 vssd1 vccd1 vccd1 _7967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2977_ _6096_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2977_/X sky130_fd_sc_hd__clkbuf_16
X_7898_ _7898_/CLK _7898_/D vssd1 vssd1 vccd1 vccd1 _7898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6947__498 _6949__500/A vssd1 vssd1 vccd1 vccd1 _8095_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _8196_/Q _4096_/X _4202_/S vssd1 vssd1 vccd1 vccd1 _4201_/A sky130_fd_sc_hd__mux2_1
X_5180_ _5191_/A vssd1 vssd1 vccd1 vccd1 _5271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4131_ _8362_/Q vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__buf_2
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4062_ _8053_/Q _8052_/Q _8051_/Q vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__and3_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ _7821_/CLK _7821_/D vssd1 vssd1 vccd1 vccd1 _7821_/Q sky130_fd_sc_hd__dfxtp_1
X_7752_ _8349_/CLK _7752_/D vssd1 vssd1 vccd1 vccd1 _7752_/Q sky130_fd_sc_hd__dfxtp_1
X_4964_ _5003_/A vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__buf_2
X_6703_ _6700_/Y _7411_/A _6753_/B vssd1 vssd1 vccd1 vccd1 _6704_/B sky130_fd_sc_hd__a21bo_1
X_3915_ _5347_/C _5347_/B _4230_/C vssd1 vssd1 vccd1 vccd1 _3989_/B sky130_fd_sc_hd__nand3b_4
X_7683_ _8349_/CLK _7683_/D vssd1 vssd1 vccd1 vccd1 _7683_/Q sky130_fd_sc_hd__dfxtp_1
X_4895_ _4910_/S vssd1 vssd1 vccd1 vccd1 _4904_/S sky130_fd_sc_hd__clkbuf_4
X_3846_ _4121_/A _5511_/A vssd1 vssd1 vccd1 vccd1 _3862_/S sky130_fd_sc_hd__nor2_2
X_6565_ _6565_/A vssd1 vssd1 vccd1 vccd1 _7865_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3346_ clkbuf_0__3346_/X vssd1 vssd1 vccd1 vccd1 _6791__395/A sky130_fd_sc_hd__clkbuf_4
X_3777_ _7999_/Q vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6496_ _6496_/A vssd1 vssd1 vccd1 vccd1 _6496_/X sky130_fd_sc_hd__buf_1
X_5516_ _5516_/A vssd1 vssd1 vccd1 vccd1 _7883_/D sky130_fd_sc_hd__clkbuf_1
X_8304_ _8304_/CLK _8304_/D vssd1 vssd1 vccd1 vccd1 _8304_/Q sky130_fd_sc_hd__dfxtp_1
X_8235_ _8235_/CLK _8235_/D vssd1 vssd1 vccd1 vccd1 _8235_/Q sky130_fd_sc_hd__dfxtp_1
X_5447_ _3828_/X _7913_/Q _5449_/S vssd1 vssd1 vccd1 vccd1 _5448_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3245_ _6601_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3245_/X sky130_fd_sc_hd__clkbuf_16
X_8166_ _8166_/CLK _8166_/D vssd1 vssd1 vccd1 vccd1 _8166_/Q sky130_fd_sc_hd__dfxtp_1
X_5378_ _5378_/A vssd1 vssd1 vccd1 vccd1 _7947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4329_ _7991_/Q vssd1 vssd1 vccd1 vccd1 _4329_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7117_ _7117_/A _7238_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7117_/X sky130_fd_sc_hd__and3_1
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8097_ _8097_/CLK _8097_/D vssd1 vssd1 vccd1 vccd1 _8097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7572__45 _7572__45/A vssd1 vssd1 vccd1 vccd1 _8384_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995__536 _6999__540/A vssd1 vssd1 vccd1 vccd1 _8133_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0__3200_ clkbuf_0__3200_/X vssd1 vssd1 vccd1 vccd1 _6477__255/A sky130_fd_sc_hd__clkbuf_4
X_4680_ _4725_/A vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__clkbuf_2
X_6438__224 _6439__225/A vssd1 vssd1 vccd1 vccd1 _7781_/CLK sky130_fd_sc_hd__inv_2
X_6350_ _7540_/A _6350_/B _6350_/C _6350_/D vssd1 vssd1 vccd1 vccd1 _6395_/A sky130_fd_sc_hd__or4_4
X_5301_ _5300_/X _7979_/Q _5309_/S vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__mux2_1
X_6281_ _6281_/A vssd1 vssd1 vccd1 vccd1 _7642_/A sky130_fd_sc_hd__clkbuf_2
X_8020_ _8020_/CLK _8020_/D vssd1 vssd1 vccd1 vccd1 _8020_/Q sky130_fd_sc_hd__dfxtp_1
X_5232_ _8281_/Q _5150_/X _5108_/B _8273_/Q vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5163_ _8283_/Q _5150_/X _5108_/B _8275_/Q vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _8259_/Q _3955_/X _4118_/S vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _3878_/X _5029_/X _5093_/X _5027_/X vssd1 vssd1 vccd1 vccd1 _8008_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4045_ _8054_/Q vssd1 vssd1 vccd1 vccd1 _4387_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7804_ _7804_/CLK _7804_/D vssd1 vssd1 vccd1 vccd1 _7804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6857__429 _6857__429/A vssd1 vssd1 vccd1 vccd1 _8024_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _7719_/Q input32/X _6008_/S vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__mux2_1
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7735_ _8066_/CLK _7735_/D vssd1 vssd1 vccd1 vccd1 _7735_/Q sky130_fd_sc_hd__dfxtp_1
X_4947_ _4347_/X _8014_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__mux2_1
X_7666_ _7992_/CLK _7666_/D vssd1 vssd1 vccd1 vccd1 _7666_/Q sky130_fd_sc_hd__dfxtp_1
X_4878_ _4878_/A vssd1 vssd1 vccd1 vccd1 _8045_/D sky130_fd_sc_hd__clkbuf_1
X_3829_ _8386_/Q _3828_/X _3832_/S vssd1 vssd1 vccd1 vccd1 _3830_/A sky130_fd_sc_hd__mux2_1
X_7597_ _7590_/X _7595_/Y _7596_/Y _6292_/X vssd1 vssd1 vccd1 vccd1 _8393_/D sky130_fd_sc_hd__a211oi_2
X_6548_ _5882_/A _7858_/Q _6552_/S vssd1 vssd1 vccd1 vccd1 _6549_/A sky130_fd_sc_hd__mux2_1
X_8218_ _8231_/CLK _8218_/D vssd1 vssd1 vccd1 vccd1 _8218_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_0 _3831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8149_ _8149_/CLK _8149_/D vssd1 vssd1 vccd1 vccd1 _8149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6608__316 _6611__319/A vssd1 vssd1 vccd1 vccd1 _7897_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5850_ _5850_/A vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__clkbuf_1
X_7312__134 _7313__135/A vssd1 vssd1 vccd1 vccd1 _8261_/CLK sky130_fd_sc_hd__inv_2
X_5781_ _7659_/Q _5552_/A _5785_/S vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__mux2_1
X_4801_ _7970_/Q _4681_/A _4642_/A _4800_/X vssd1 vssd1 vccd1 vccd1 _4802_/C sky130_fd_sc_hd__o211a_1
X_7520_ _8352_/Q _7511_/X _7518_/X _7519_/X vssd1 vssd1 vccd1 vccd1 _8352_/D sky130_fd_sc_hd__o211a_1
X_4732_ _4730_/X _7872_/Q _7776_/Q _4731_/X vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__a22o_1
X_7451_ _7491_/B vssd1 vssd1 vccd1 vccd1 _7466_/A sky130_fd_sc_hd__clkbuf_2
X_4663_ _8199_/Q _7817_/Q _7801_/Q _7785_/Q _4571_/A _4569_/X vssd1 vssd1 vccd1 vccd1
+ _4664_/B sky130_fd_sc_hd__mux4_1
X_6402_ _6342_/A _6350_/D _6347_/Y vssd1 vssd1 vccd1 vccd1 _6403_/B sky130_fd_sc_hd__a21bo_1
X_4594_ _4669_/S vssd1 vssd1 vccd1 vccd1 _4594_/X sky130_fd_sc_hd__clkbuf_2
X_7382_ _7382_/A vssd1 vssd1 vccd1 vccd1 _7382_/X sky130_fd_sc_hd__buf_1
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6333_ _7727_/Q _6320_/X _6324_/X _6332_/X vssd1 vssd1 vccd1 vccd1 _7727_/D sky130_fd_sc_hd__a211o_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6264_ _7714_/Q _6216_/X _6263_/X vssd1 vssd1 vccd1 vccd1 _7714_/D sky130_fd_sc_hd__a21o_1
X_8003_ _8003_/CLK _8003_/D vssd1 vssd1 vccd1 vccd1 _8003_/Q sky130_fd_sc_hd__dfxtp_1
X_5215_ _3887_/X _5029_/A _5214_/X vssd1 vssd1 vccd1 vccd1 _5215_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6195_ _8203_/Q vssd1 vssd1 vccd1 vccd1 _7262_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5146_ _8315_/Q _5187_/A _5125_/A _8307_/Q _4987_/A vssd1 vssd1 vccd1 vccd1 _5146_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _4965_/A _5076_/X _5090_/A vssd1 vssd1 vccd1 vccd1 _5077_/X sky130_fd_sc_hd__a21o_1
X_4028_ _8280_/Q _3966_/X _4036_/S vssd1 vssd1 vccd1 vccd1 _4029_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3261_ clkbuf_0__3261_/X vssd1 vssd1 vccd1 vccd1 _6677__367/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0_0__3192_ clkbuf_0__3192_/X vssd1 vssd1 vccd1 vccd1 _6439__225/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5979_ _7714_/Q input25/X _5991_/S vssd1 vssd1 vccd1 vccd1 _5979_/X sky130_fd_sc_hd__mux2_4
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7385__18 _7385__18/A vssd1 vssd1 vccd1 vccd1 _8320_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7718_ _8391_/CLK _7718_/D vssd1 vssd1 vccd1 vccd1 _7718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7649_ _7649_/CLK _7649_/D vssd1 vssd1 vccd1 vccd1 _7649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2976_ clkbuf_0__2976_/X vssd1 vssd1 vccd1 vccd1 _6095__185/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7190__113 _7190__113/A vssd1 vssd1 vccd1 vccd1 _8212_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6508__280 _6508__280/A vssd1 vssd1 vccd1 vccd1 _7837_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5000_ _4988_/X _4989_/X _4999_/X vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__a21o_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6951_ _6957_/A vssd1 vssd1 vccd1 vccd1 _6951_/X sky130_fd_sc_hd__buf_1
X_6481__258 _6482__259/A vssd1 vssd1 vccd1 vccd1 _7815_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5902_ _5902_/A vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__clkbuf_1
X_5833_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5833_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3594_ clkbuf_0__3594_/X vssd1 vssd1 vccd1 vccd1 _7356__170/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7503_ _7402_/B _7510_/A _7502_/X _7490_/Y vssd1 vssd1 vccd1 vccd1 _7503_/X sky130_fd_sc_hd__a211o_1
X_5764_ _5764_/A vssd1 vssd1 vccd1 vccd1 _7711_/D sky130_fd_sc_hd__clkbuf_1
X_5695_ _7786_/Q _5581_/X _5699_/S vssd1 vssd1 vccd1 vccd1 _5696_/A sky130_fd_sc_hd__mux2_1
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__clkbuf_2
X_7434_ _8394_/Q _6706_/B _6704_/B _7117_/A vssd1 vssd1 vccd1 vccd1 _7435_/D sky130_fd_sc_hd__o2bb2a_1
X_4646_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__buf_2
X_4577_ _4867_/B _4563_/X _4576_/X vssd1 vssd1 vccd1 vccd1 _4577_/X sky130_fd_sc_hd__a21o_1
X_6316_ _7117_/A _6326_/B _6322_/C _6326_/D vssd1 vssd1 vccd1 vccd1 _6316_/X sky130_fd_sc_hd__and4_1
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6247_ _6221_/X _6229_/X _6245_/X _6246_/X vssd1 vssd1 vccd1 vccd1 _6247_/X sky130_fd_sc_hd__a31o_1
X_6178_ _7546_/B _7699_/Q _6180_/S vssd1 vssd1 vccd1 vccd1 _6179_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5129_ _8276_/Q _5125_/X _5084_/A _5128_/X vssd1 vssd1 vccd1 vccd1 _5129_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3244_ clkbuf_0__3244_/X vssd1 vssd1 vccd1 vccd1 _6597__307/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952__501 _6956__505/A vssd1 vssd1 vccd1 vccd1 _8098_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7054__83 _7055__84/A vssd1 vssd1 vccd1 vccd1 _8180_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5480_ _5480_/A vssd1 vssd1 vccd1 vccd1 _7899_/D sky130_fd_sc_hd__clkbuf_1
X_4500_ _4500_/A vssd1 vssd1 vccd1 vccd1 _8078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4431_ _4431_/A vssd1 vssd1 vccd1 vccd1 _8108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7150_ _8225_/Q _7150_/B _7150_/C _7150_/D vssd1 vssd1 vccd1 vccd1 _7166_/A sky130_fd_sc_hd__and4_2
X_4362_ _8133_/Q _4137_/X _4366_/S vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4211_/X _8160_/Q _4297_/S vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__mux2_1
X_6032_ _6079_/D vssd1 vssd1 vccd1 vccd1 _6032_/X sky130_fd_sc_hd__buf_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7983_ _7983_/CLK _7983_/D vssd1 vssd1 vccd1 vccd1 _7983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6865_ _6871_/A vssd1 vssd1 vccd1 vccd1 _6865_/X sky130_fd_sc_hd__buf_1
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5816_ _6036_/A _7861_/Q _5817_/C _5815_/X _7644_/Q vssd1 vssd1 vccd1 vccd1 _5966_/A
+ sky130_fd_sc_hd__a41oi_4
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5747_ _7763_/Q _5552_/A _5753_/S vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5678_ _5678_/A vssd1 vssd1 vccd1 vccd1 _7794_/D sky130_fd_sc_hd__clkbuf_1
X_7417_ _7117_/A _6704_/B _6706_/B _8394_/Q vssd1 vssd1 vccd1 vccd1 _7417_/X sky130_fd_sc_hd__o2bb2a_1
X_8397_ _8397_/CLK _8397_/D vssd1 vssd1 vccd1 vccd1 _8397_/Q sky130_fd_sc_hd__dfxtp_1
X_4629_ _4549_/X _4614_/X _4618_/X _4628_/X vssd1 vssd1 vccd1 vccd1 _4629_/X sky130_fd_sc_hd__a31o_1
X_7279_ _8237_/Q _7283_/B vssd1 vssd1 vccd1 vccd1 _7279_/X sky130_fd_sc_hd__or2_1
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6432__219 _6432__219/A vssd1 vssd1 vccd1 vccd1 _7776_/CLK sky130_fd_sc_hd__inv_2
X_6586__300 _6586__300/A vssd1 vssd1 vccd1 vccd1 _7881_/CLK sky130_fd_sc_hd__inv_2
Xoutput93 _5906_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6959__507 _6961__509/A vssd1 vssd1 vccd1 vccd1 _8104_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7027__61 _7029__63/A vssd1 vssd1 vccd1 vccd1 _8158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _7996_/Q _4982_/B vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__and2_1
X_3931_ _3931_/A vssd1 vssd1 vccd1 vccd1 _8314_/D sky130_fd_sc_hd__clkbuf_1
X_3862_ _8374_/Q _3840_/X _3862_/S vssd1 vssd1 vccd1 vccd1 _3863_/A sky130_fd_sc_hd__mux2_1
X_6650_ _6650_/A vssd1 vssd1 vccd1 vccd1 _6650_/X sky130_fd_sc_hd__buf_1
X_6593__304 _6594__305/A vssd1 vssd1 vccd1 vccd1 _7885_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5601_ _5547_/X _7828_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__mux2_1
X_6581_ _6581_/A vssd1 vssd1 vccd1 vccd1 _6581_/X sky130_fd_sc_hd__buf_1
X_5532_ _5532_/A vssd1 vssd1 vccd1 vccd1 _7876_/D sky130_fd_sc_hd__clkbuf_1
X_3793_ _3793_/A _3793_/B _3793_/C vssd1 vssd1 vccd1 vccd1 _6340_/B sky130_fd_sc_hd__and3_2
X_8320_ _8320_/CLK _8320_/D vssd1 vssd1 vccd1 vccd1 _8320_/Q sky130_fd_sc_hd__dfxtp_1
X_5463_ _7906_/Q _4211_/A _5467_/S vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__mux2_1
X_8251_ _8251_/CLK _8251_/D vssd1 vssd1 vccd1 vccd1 _8251_/Q sky130_fd_sc_hd__dfxtp_1
X_7202_ _7202_/A _7202_/B vssd1 vssd1 vccd1 vccd1 _7238_/C sky130_fd_sc_hd__nor2_1
X_4414_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__buf_2
X_5394_ _5394_/A vssd1 vssd1 vccd1 vccd1 _7937_/D sky130_fd_sc_hd__clkbuf_1
X_8182_ _8182_/CLK _8182_/D vssd1 vssd1 vccd1 vccd1 _8182_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3261_ _6675_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3261_/X sky130_fd_sc_hd__clkbuf_16
X_7133_ _7208_/A _7204_/A _7199_/A _8216_/Q vssd1 vssd1 vccd1 vccd1 _7134_/B sky130_fd_sc_hd__a31o_1
Xclkbuf_0__3192_ _6434_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3192_/X sky130_fd_sc_hd__clkbuf_16
X_4345_ _4344_/X _8140_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6784__389 _6785__390/A vssd1 vssd1 vccd1 vccd1 _7974_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4276_ _8167_/Q _4131_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6015_ _6015_/A vssd1 vssd1 vccd1 vccd1 _6015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7966_ _7966_/CLK _7966_/D vssd1 vssd1 vccd1 vccd1 _7966_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2976_ _6090_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2976_/X sky130_fd_sc_hd__clkbuf_16
X_7897_ _7897_/CLK _7897_/D vssd1 vssd1 vccd1 vccd1 _7897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7010__549 _7010__549/A vssd1 vssd1 vccd1 vccd1 _8146_/CLK sky130_fd_sc_hd__inv_2
X_7373__8 _7374__9/A vssd1 vssd1 vccd1 vccd1 _8310_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_wb_clk_i _7717_/CLK vssd1 vssd1 vccd1 vccd1 _7989_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4130_ _4130_/A vssd1 vssd1 vccd1 vccd1 _8254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4061_ _8055_/Q _8050_/Q vssd1 vssd1 vccd1 vccd1 _4536_/C sky130_fd_sc_hd__xnor2_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7820_ _7820_/CLK _7820_/D vssd1 vssd1 vccd1 vccd1 _7820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7751_ _8348_/CLK _7751_/D vssd1 vssd1 vccd1 vccd1 _7751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _5017_/A vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__clkbuf_2
X_7682_ _8349_/CLK _7682_/D vssd1 vssd1 vccd1 vccd1 _7682_/Q sky130_fd_sc_hd__dfxtp_1
X_6702_ _6702_/A _6702_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _6753_/B sky130_fd_sc_hd__nand3_2
X_3914_ _8001_/Q vssd1 vssd1 vccd1 vccd1 _5347_/B sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3414_ clkbuf_0__3414_/X vssd1 vssd1 vccd1 vccd1 _7080__104/A sky130_fd_sc_hd__clkbuf_4
X_4894_ _5635_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _4910_/S sky130_fd_sc_hd__nor2_2
X_3845_ _4286_/B _4230_/C _5347_/C vssd1 vssd1 vccd1 vccd1 _5511_/A sky130_fd_sc_hd__nand3b_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6564_ _7865_/Q _5897_/A _6564_/S vssd1 vssd1 vccd1 vccd1 _6565_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3345_ clkbuf_0__3345_/X vssd1 vssd1 vccd1 vccd1 _6785__390/A sky130_fd_sc_hd__clkbuf_4
X_3776_ _4286_/A _4120_/C _4286_/B vssd1 vssd1 vccd1 vccd1 _4507_/A sky130_fd_sc_hd__or3b_2
XFILLER_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8303_ _8303_/CLK _8303_/D vssd1 vssd1 vccd1 vccd1 _8303_/Q sky130_fd_sc_hd__dfxtp_1
X_5515_ _7883_/Q _4208_/A _5521_/S vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8234_ _8235_/CLK _8234_/D vssd1 vssd1 vccd1 vccd1 _8234_/Q sky130_fd_sc_hd__dfxtp_1
X_5446_ _5446_/A vssd1 vssd1 vccd1 vccd1 _7914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7361__174 _7362__175/A vssd1 vssd1 vccd1 vccd1 _8301_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3244_ _6595_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3244_/X sky130_fd_sc_hd__clkbuf_16
X_5377_ _7947_/Q _4520_/X _5377_/S vssd1 vssd1 vccd1 vccd1 _5378_/A sky130_fd_sc_hd__mux2_1
X_8165_ _8165_/CLK _8165_/D vssd1 vssd1 vccd1 vccd1 _8165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7116_ _7119_/A _7150_/C _7119_/C _8223_/Q vssd1 vssd1 vccd1 vccd1 _7238_/B sky130_fd_sc_hd__a31o_1
X_4328_ _4328_/A vssd1 vssd1 vccd1 vccd1 _8146_/D sky130_fd_sc_hd__clkbuf_1
X_8096_ _8096_/CLK _8096_/D vssd1 vssd1 vccd1 vccd1 _8096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4259_ _4259_/A vssd1 vssd1 vccd1 vccd1 _8175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _7949_/CLK _7949_/D vssd1 vssd1 vccd1 vccd1 _7949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7557__32 _7559__34/A vssd1 vssd1 vccd1 vccd1 _8371_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7021__56 _7022__57/A vssd1 vssd1 vccd1 vccd1 _8153_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6212__198 _6213__199/A vssd1 vssd1 vccd1 vccd1 _7710_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5300_ _5564_/A vssd1 vssd1 vccd1 vccd1 _5300_/X sky130_fd_sc_hd__buf_2
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6280_ _8003_/Q _6254_/Y _6279_/X _6243_/X vssd1 vssd1 vccd1 vccd1 _6280_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5231_ _8187_/Q _8257_/Q _5231_/S vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5162_ _8189_/Q _8259_/Q _5224_/S vssd1 vssd1 vccd1 vccd1 _5162_/X sky130_fd_sc_hd__mux2_1
X_5093_ _8008_/Q _4955_/X _5031_/X _5092_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _5093_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4113_ _4113_/A vssd1 vssd1 vccd1 vccd1 _8260_/D sky130_fd_sc_hd__clkbuf_1
X_4044_ _7992_/Q vssd1 vssd1 vccd1 vccd1 _4044_/X sky130_fd_sc_hd__clkbuf_4
X_6445__229 _6446__230/A vssd1 vssd1 vccd1 vccd1 _7786_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7803_ _7803_/CLK _7803_/D vssd1 vssd1 vccd1 vccd1 _7803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5995_ _6029_/S vssd1 vssd1 vccd1 vccd1 _6008_/S sky130_fd_sc_hd__clkbuf_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7734_ _8066_/CLK _7734_/D vssd1 vssd1 vccd1 vccd1 _7734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _4946_/A vssd1 vssd1 vccd1 vccd1 _8015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _8045_/Q _4386_/X _4885_/S vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__mux2_1
X_7665_ _7012_/A _7665_/D vssd1 vssd1 vccd1 vccd1 _7665_/Q sky130_fd_sc_hd__dfxtp_1
X_7596_ _7596_/A _7599_/B vssd1 vssd1 vccd1 vccd1 _7596_/Y sky130_fd_sc_hd__nor2_1
X_3828_ _8362_/Q vssd1 vssd1 vccd1 vccd1 _3828_/X sky130_fd_sc_hd__buf_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6547_ _6547_/A vssd1 vssd1 vccd1 vccd1 _7857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6478_ _6478_/A vssd1 vssd1 vccd1 vccd1 _6478_/X sky130_fd_sc_hd__buf_1
X_8217_ _8239_/CLK _8217_/D vssd1 vssd1 vccd1 vccd1 _8217_/Q sky130_fd_sc_hd__dfxtp_1
X_5429_ _7921_/Q _4517_/X _5431_/S vssd1 vssd1 vccd1 vccd1 _5430_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8148_ _8148_/CLK _8148_/D vssd1 vssd1 vccd1 vccd1 _8148_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_1 _5123_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8079_ _8079_/CLK _8079_/D vssd1 vssd1 vccd1 vccd1 _8079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4800_ _8031_/Q _4676_/A _4799_/X _4729_/A vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5780_ _5780_/A vssd1 vssd1 vccd1 vccd1 _7660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4731_/A vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__clkbuf_2
X_7450_ _7450_/A _7450_/B vssd1 vssd1 vccd1 vccd1 _7491_/B sky130_fd_sc_hd__and2_1
X_4662_ _4557_/A _4659_/X _4661_/X vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6401_ _7595_/A _6185_/C _6251_/X vssd1 vssd1 vccd1 vccd1 _6403_/A sky130_fd_sc_hd__a21oi_1
X_7551__27 _7553__29/A vssd1 vssd1 vccd1 vccd1 _8366_/CLK sky130_fd_sc_hd__inv_2
X_4593_ _4590_/X _4591_/X _4593_/S vssd1 vssd1 vccd1 vccd1 _4593_/X sky130_fd_sc_hd__mux2_1
X_6332_ _7593_/A _6337_/B _6332_/C _6337_/D vssd1 vssd1 vccd1 vccd1 _6332_/X sky130_fd_sc_hd__and4_1
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6263_ _6270_/A _6260_/X _6262_/X _6246_/X vssd1 vssd1 vccd1 vccd1 _6263_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _6838_/A vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__clkbuf_2
X_8002_ _8002_/CLK _8002_/D vssd1 vssd1 vccd1 vccd1 _8002_/Q sky130_fd_sc_hd__dfxtp_1
X_6863__434 _6863__434/A vssd1 vssd1 vccd1 vccd1 _8029_/CLK sky130_fd_sc_hd__inv_2
X_6194_ _8231_/Q _6194_/B vssd1 vssd1 vccd1 vccd1 _6194_/X sky130_fd_sc_hd__and2b_1
X_6824__407 _6826__409/A vssd1 vssd1 vccd1 vccd1 _8000_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5145_ _8291_/Q _8299_/Q _5224_/S vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__mux2_1
X_5076_ _8277_/Q _8261_/Q _8191_/Q _8285_/Q _5231_/S _5010_/X vssd1 vssd1 vccd1 vccd1
+ _5076_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0_0__3260_ clkbuf_0__3260_/X vssd1 vssd1 vccd1 vccd1 _6674__365/A sky130_fd_sc_hd__clkbuf_4
X_4027_ _4042_/S vssd1 vssd1 vccd1 vccd1 _4036_/S sky130_fd_sc_hd__buf_2
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3191_ clkbuf_0__3191_/X vssd1 vssd1 vccd1 vccd1 _6432__219/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _6029_/S vssd1 vssd1 vccd1 vccd1 _5991_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7717_ _7717_/CLK _7717_/D vssd1 vssd1 vccd1 vccd1 _7717_/Q sky130_fd_sc_hd__dfxtp_1
X_4929_ _4929_/A vssd1 vssd1 vccd1 vccd1 _8022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7648_ _7648_/CLK _7648_/D vssd1 vssd1 vccd1 vccd1 _7648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7579_ _7608_/A _7579_/B vssd1 vssd1 vccd1 vccd1 _7579_/Y sky130_fd_sc_hd__nand2_1
X_6614__321 _6615__322/A vssd1 vssd1 vccd1 vccd1 _7902_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2975_ clkbuf_0__2975_/X vssd1 vssd1 vccd1 vccd1 _6087__178/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3389_ clkbuf_0__3389_/X vssd1 vssd1 vccd1 vccd1 _6956__505/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6950_ _6981_/A vssd1 vssd1 vccd1 vccd1 _6950_/X sky130_fd_sc_hd__buf_1
X_5901_ _5901_/A _5903_/B vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__or2_1
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _6554_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__and2_1
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3593_ clkbuf_0__3593_/X vssd1 vssd1 vccd1 vccd1 _7349__164/A sky130_fd_sc_hd__clkbuf_4
X_5763_ _5547_/X _7711_/Q _5771_/S vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__mux2_1
X_7502_ _8348_/Q _7498_/A _7501_/Y vssd1 vssd1 vccd1 vccd1 _7502_/X sky130_fd_sc_hd__o21a_1
X_4714_ _4714_/A vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__clkbuf_2
X_5694_ _5694_/A vssd1 vssd1 vccd1 vccd1 _7787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7390__22 _7390__22/A vssd1 vssd1 vccd1 vccd1 _8324_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4645_ _7650_/Q _7658_/Q _7709_/Q _7810_/Q _4571_/A _4596_/X vssd1 vssd1 vccd1 vccd1
+ _4645_/X sky130_fd_sc_hd__mux4_1
X_7433_ _6719_/A _7429_/Y _7430_/X _7431_/Y _7432_/Y vssd1 vssd1 vccd1 vccd1 _7435_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4576_ _4567_/X _4572_/X _4575_/X vssd1 vssd1 vccd1 vccd1 _4576_/X sky130_fd_sc_hd__a21o_1
X_7364_ _7382_/A vssd1 vssd1 vccd1 vccd1 _7364_/X sky130_fd_sc_hd__buf_1
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6315_ _8397_/Q vssd1 vssd1 vccd1 vccd1 _7117_/A sky130_fd_sc_hd__buf_2
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7295_ _7295_/A vssd1 vssd1 vccd1 vccd1 _7295_/X sky130_fd_sc_hd__buf_1
X_6246_ _6281_/A vssd1 vssd1 vccd1 vccd1 _6246_/X sky130_fd_sc_hd__clkbuf_2
X_6177_ _6177_/A vssd1 vssd1 vccd1 vccd1 _7698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5128_ _8284_/Q _5126_/X _5130_/A _5127_/X vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__o22a_1
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5059_ _4988_/X _5056_/X _5058_/X vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0_0__3243_ clkbuf_0__3243_/X vssd1 vssd1 vccd1 vccd1 _6594__305/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8430__205 vssd1 vssd1 vccd1 vccd1 _8430__205/HI core1Index[5] sky130_fd_sc_hd__conb_1
XFILLER_107_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__2973_ clkbuf_0__2973_/X vssd1 vssd1 vccd1 vccd1 _6502_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3387_ clkbuf_0__3387_/X vssd1 vssd1 vccd1 vccd1 _6945__496/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4430_ _8108_/Q _4407_/X _4432_/S vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__mux2_1
X_4361_ _4361_/A vssd1 vssd1 vccd1 vccd1 _8134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4292_/A vssd1 vssd1 vccd1 vccd1 _8161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6031_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__clkbuf_4
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7982_ _7982_/CLK _7982_/D vssd1 vssd1 vccd1 vccd1 _7982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5815_ _7862_/Q _7863_/Q _7864_/Q vssd1 vssd1 vccd1 vccd1 _5815_/X sky130_fd_sc_hd__and3_2
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5746_ _5746_/A vssd1 vssd1 vccd1 vccd1 _7764_/D sky130_fd_sc_hd__clkbuf_1
X_5677_ _7794_/Q _5581_/X _5681_/S vssd1 vssd1 vccd1 vccd1 _5678_/A sky130_fd_sc_hd__mux2_1
X_7416_ _8392_/Q _7416_/B _7416_/C vssd1 vssd1 vccd1 vccd1 _7416_/X sky130_fd_sc_hd__and3_1
X_4628_ _4588_/X _4623_/X _4627_/X _4674_/A vssd1 vssd1 vccd1 vccd1 _4628_/X sky130_fd_sc_hd__o211a_1
X_8396_ _8397_/CLK _8396_/D vssd1 vssd1 vccd1 vccd1 _8396_/Q sky130_fd_sc_hd__dfxtp_4
X_7325__145 _7325__145/A vssd1 vssd1 vccd1 vccd1 _8272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4559_ _4559_/A vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__clkbuf_4
X_7278_ _8008_/Q _7266_/X _7277_/X _7269_/X vssd1 vssd1 vccd1 vccd1 _8236_/D sky130_fd_sc_hd__o211a_1
X_6229_ _7143_/A _6839_/C _6228_/X vssd1 vssd1 vccd1 vccd1 _6229_/X sky130_fd_sc_hd__a21o_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3241_ clkbuf_0__3241_/X vssd1 vssd1 vccd1 vccd1 _6815_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6917__474 _6918__475/A vssd1 vssd1 vccd1 vccd1 _8071_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput94 _5928_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6627__331 _6628__332/A vssd1 vssd1 vccd1 vccd1 _7912_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _3887_/X _8314_/Q _3932_/S vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _3861_/A vssd1 vssd1 vccd1 vccd1 _8375_/D sky130_fd_sc_hd__clkbuf_1
X_3792_ _3893_/A _4949_/A _5249_/B _3790_/Y _3791_/X vssd1 vssd1 vccd1 vccd1 _3793_/C
+ sky130_fd_sc_hd__o221a_1
X_5600_ _5615_/S vssd1 vssd1 vccd1 vccd1 _5609_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5531_ _5278_/X _7876_/Q _5539_/S vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__mux2_1
X_8250_ _8250_/CLK _8250_/D vssd1 vssd1 vccd1 vccd1 _8250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7201_ _7219_/A vssd1 vssd1 vccd1 vccd1 _7218_/A sky130_fd_sc_hd__clkbuf_2
X_5462_ _5462_/A vssd1 vssd1 vccd1 vccd1 _7907_/D sky130_fd_sc_hd__clkbuf_1
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _4930_/C sky130_fd_sc_hd__buf_2
X_5393_ _7937_/Q _4517_/X _5395_/S vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3260_ _6669_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3260_/X sky130_fd_sc_hd__clkbuf_16
X_8181_ _8181_/CLK _8181_/D vssd1 vssd1 vccd1 vccd1 _8181_/Q sky130_fd_sc_hd__dfxtp_1
X_7132_ _7140_/B vssd1 vssd1 vccd1 vccd1 _7199_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__3191_ _6428_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3191_/X sky130_fd_sc_hd__clkbuf_16
X_4344_ _7986_/Q vssd1 vssd1 vccd1 vccd1 _4344_/X sky130_fd_sc_hd__buf_2
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7063_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7063_/X sky130_fd_sc_hd__buf_1
X_6014_ _7673_/Q _6013_/X _6023_/S vssd1 vssd1 vccd1 vccd1 _6015_/A sky130_fd_sc_hd__mux2_4
XFILLER_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _4275_/A vssd1 vssd1 vccd1 vccd1 _8168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7965_ _7965_/CLK _7965_/D vssd1 vssd1 vccd1 vccd1 _7965_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2975_ _6084_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2975_/X sky130_fd_sc_hd__clkbuf_16
X_7896_ _7896_/CLK _7896_/D vssd1 vssd1 vccd1 vccd1 _7896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5729_ _7771_/Q _5552_/A _5735_/S vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6494__269 _6495__270/A vssd1 vssd1 vccd1 vccd1 _7826_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8379_ _8379_/CLK _8379_/D vssd1 vssd1 vccd1 vccd1 _8379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3389_ _6951_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3389_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8436__211 vssd1 vssd1 vccd1 vccd1 _8436__211/HI manufacturerID[3] sky130_fd_sc_hd__conb_1
XFILLER_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6850__425 _6850__425/A vssd1 vssd1 vccd1 vccd1 _8020_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6965__512 _6966__513/A vssd1 vssd1 vccd1 vccd1 _8109_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4060_ _8052_/Q _4536_/B _4536_/A _4056_/Y vssd1 vssd1 vccd1 vccd1 _4060_/X sky130_fd_sc_hd__a211o_1
XFILLER_3_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6408__200 _6408__200/A vssd1 vssd1 vccd1 vccd1 _7757_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7750_ _8348_/CLK _7750_/D vssd1 vssd1 vccd1 vccd1 _7750_/Q sky130_fd_sc_hd__dfxtp_1
X_4962_ _4982_/B _5126_/A vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__or2_1
X_7681_ _8348_/CLK _7681_/D vssd1 vssd1 vccd1 vccd1 _7681_/Q sky130_fd_sc_hd__dfxtp_1
X_6701_ _8339_/Q _6702_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _7411_/A sky130_fd_sc_hd__nand3_2
X_3913_ _5439_/A vssd1 vssd1 vccd1 vccd1 _5348_/A sky130_fd_sc_hd__buf_2
X_4893_ _4930_/C _4930_/B _4930_/A vssd1 vssd1 vccd1 vccd1 _5725_/B sky130_fd_sc_hd__nand3b_4
X_3844_ _4286_/A vssd1 vssd1 vccd1 vccd1 _5347_/C sky130_fd_sc_hd__buf_2
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3413_ clkbuf_0__3413_/X vssd1 vssd1 vccd1 vccd1 _7295_/A sky130_fd_sc_hd__clkbuf_4
X_6632_ _6632_/A vssd1 vssd1 vccd1 vccd1 _6632_/X sky130_fd_sc_hd__buf_1
XFILLER_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3344_ clkbuf_0__3344_/X vssd1 vssd1 vccd1 vccd1 _6777__383/A sky130_fd_sc_hd__clkbuf_4
X_6563_ _6563_/A vssd1 vssd1 vccd1 vccd1 _7864_/D sky130_fd_sc_hd__clkbuf_1
X_3775_ _8001_/Q vssd1 vssd1 vccd1 vccd1 _4286_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6790__394 _6790__394/A vssd1 vssd1 vccd1 vccd1 _7979_/CLK sky130_fd_sc_hd__inv_2
X_5514_ _5514_/A vssd1 vssd1 vccd1 vccd1 _7884_/D sky130_fd_sc_hd__clkbuf_1
X_8302_ _8302_/CLK _8302_/D vssd1 vssd1 vccd1 vccd1 _8302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8233_ _8235_/CLK _8233_/D vssd1 vssd1 vccd1 vccd1 _8233_/Q sky130_fd_sc_hd__dfxtp_1
X_5445_ _3825_/X _7914_/Q _5449_/S vssd1 vssd1 vccd1 vccd1 _5446_/A sky130_fd_sc_hd__mux2_1
X_8164_ _8164_/CLK _8164_/D vssd1 vssd1 vccd1 vccd1 _8164_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3243_ _6589_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3243_/X sky130_fd_sc_hd__clkbuf_16
X_7115_ _8396_/Q _7115_/B vssd1 vssd1 vccd1 vccd1 _7146_/B sky130_fd_sc_hd__xor2_1
X_5376_ _5376_/A vssd1 vssd1 vccd1 vccd1 _7948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4327_ _4323_/X _8146_/Q _4339_/S vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__mux2_1
X_8095_ _8095_/CLK _8095_/D vssd1 vssd1 vccd1 vccd1 _8095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4258_ _4214_/X _8175_/Q _4260_/S vssd1 vssd1 vccd1 vccd1 _4259_/A sky130_fd_sc_hd__mux2_1
X_4189_ _4189_/A vssd1 vssd1 vccd1 vccd1 _8202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _7948_/CLK _7948_/D vssd1 vssd1 vccd1 vccd1 _7948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7879_ _7879_/CLK _7879_/D vssd1 vssd1 vccd1 vccd1 _7879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7338__155 _7338__155/A vssd1 vssd1 vccd1 vccd1 _8282_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5230_ _5230_/A _5230_/B _5230_/C vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__or3_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161_ _5230_/A _5161_/B _5161_/C vssd1 vssd1 vccd1 vccd1 _5161_/X sky130_fd_sc_hd__or3_1
XFILLER_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5092_ _5002_/X _5078_/X _5082_/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__a31o_2
X_4112_ _8260_/Q _3951_/X _4112_/S vssd1 vssd1 vccd1 vccd1 _4113_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4043_ _4043_/A vssd1 vssd1 vccd1 vccd1 _8273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7802_ _7802_/CLK _7802_/D vssd1 vssd1 vccd1 vccd1 _7802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5994_ _5994_/A vssd1 vssd1 vccd1 vccd1 _5994_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7733_ _8065_/CLK _7733_/D vssd1 vssd1 vccd1 vccd1 _7733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4945_ _4344_/X _8015_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__mux2_1
X_7664_ _7697_/CLK _7664_/D vssd1 vssd1 vccd1 vccd1 _7664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4891_/S vssd1 vssd1 vccd1 vccd1 _4885_/S sky130_fd_sc_hd__clkbuf_4
X_7595_ _7595_/A _7595_/B vssd1 vssd1 vccd1 vccd1 _7595_/Y sky130_fd_sc_hd__nand2_1
X_3827_ _3827_/A vssd1 vssd1 vccd1 vccd1 _8387_/D sky130_fd_sc_hd__clkbuf_1
X_6546_ _5880_/A _7857_/Q _6546_/S vssd1 vssd1 vccd1 vccd1 _6547_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8216_ _8223_/CLK _8216_/D vssd1 vssd1 vccd1 vccd1 _8216_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3189_ clkbuf_0__3189_/X vssd1 vssd1 vccd1 vccd1 _6418__207/A sky130_fd_sc_hd__clkbuf_4
X_5428_ _5428_/A vssd1 vssd1 vccd1 vccd1 _7922_/D sky130_fd_sc_hd__clkbuf_1
X_5359_ _5359_/A vssd1 vssd1 vccd1 vccd1 _7955_/D sky130_fd_sc_hd__clkbuf_1
X_8147_ _8147_/CLK _8147_/D vssd1 vssd1 vccd1 vccd1 _8147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_2 _5124_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8078_ _8078_/CLK _8078_/D vssd1 vssd1 vccd1 vccd1 _8078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4730_/A vssd1 vssd1 vccd1 vccd1 _4730_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4661_ _4594_/X _4660_/X _4575_/X vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6400_ _6400_/A vssd1 vssd1 vccd1 vccd1 _7595_/A sky130_fd_sc_hd__clkbuf_2
X_6331_ _8392_/Q vssd1 vssd1 vccd1 vccd1 _7593_/A sky130_fd_sc_hd__clkbuf_4
X_4592_ _4641_/A vssd1 vssd1 vccd1 vccd1 _4593_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_115_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6262_ _8056_/Q _6254_/Y _6261_/X _6243_/X vssd1 vssd1 vccd1 vccd1 _6262_/X sky130_fd_sc_hd__a22o_1
X_6451__234 _6451__234/A vssd1 vssd1 vccd1 vccd1 _7791_/CLK sky130_fd_sc_hd__inv_2
X_8001_ _8001_/CLK _8001_/D vssd1 vssd1 vccd1 vccd1 _8001_/Q sky130_fd_sc_hd__dfxtp_2
X_6193_ _8232_/Q _8233_/Q _8234_/Q _8235_/Q _7258_/B _8230_/Q vssd1 vssd1 vccd1 vccd1
+ _6194_/B sky130_fd_sc_hd__mux4_1
X_5213_ _8005_/Q _4955_/X _4953_/X vssd1 vssd1 vccd1 vccd1 _5213_/Y sky130_fd_sc_hd__a21oi_1
X_5144_ _3881_/X _5029_/X _5143_/X _5027_/X vssd1 vssd1 vccd1 vccd1 _8007_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5075_ _8378_/Q _7948_/Q _7881_/Q _8370_/Q _4978_/X _4995_/X vssd1 vssd1 vccd1 vccd1
+ _5075_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _4121_/A _4204_/B vssd1 vssd1 vccd1 vccd1 _4042_/S sky130_fd_sc_hd__nor2_2
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3190_ clkbuf_0__3190_/X vssd1 vssd1 vccd1 vccd1 _6424__212/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _5977_/A vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__clkbuf_1
X_7716_ _7989_/CLK _7716_/D vssd1 vssd1 vccd1 vccd1 _7716_/Q sky130_fd_sc_hd__dfxtp_1
X_4928_ _8022_/Q _4410_/X _4928_/S vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7647_ _7647_/CLK _7647_/D vssd1 vssd1 vccd1 vccd1 _7647_/Q sky130_fd_sc_hd__dfxtp_1
X_4859_ _4859_/A vssd1 vssd1 vccd1 vccd1 _8052_/D sky130_fd_sc_hd__clkbuf_1
X_6529_ _6529_/A vssd1 vssd1 vccd1 vccd1 _7849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2974_ clkbuf_0__2974_/X vssd1 vssd1 vccd1 vccd1 _6209_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7066__93 _7066__93/A vssd1 vssd1 vccd1 vccd1 _8190_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3388_ clkbuf_0__3388_/X vssd1 vssd1 vccd1 vccd1 _6957_/A sky130_fd_sc_hd__clkbuf_4
X_6621__326 _6622__327/A vssd1 vssd1 vccd1 vccd1 _7907_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5900_ _5900_/A vssd1 vssd1 vccd1 vccd1 _5900_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5831_ _5831_/A vssd1 vssd1 vccd1 vccd1 _5831_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3592_ clkbuf_0__3592_/X vssd1 vssd1 vccd1 vccd1 _7341__157/A sky130_fd_sc_hd__clkbuf_4
X_5762_ _5777_/S vssd1 vssd1 vccd1 vccd1 _5771_/S sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_6_wb_clk_i _7717_/CLK vssd1 vssd1 vccd1 vccd1 _7992_/CLK sky130_fd_sc_hd__clkbuf_16
X_7501_ _8348_/Q _7498_/A _7527_/B vssd1 vssd1 vccd1 vccd1 _7501_/Y sky130_fd_sc_hd__a21oi_1
X_4713_ _4567_/X _4709_/X _4712_/X _4588_/X vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__a211o_1
X_5693_ _7787_/Q _5578_/X _5699_/S vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__mux2_1
X_7432_ _7432_/A _7432_/B vssd1 vssd1 vccd1 vccd1 _7432_/Y sky130_fd_sc_hd__xnor2_1
X_4644_ _4664_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4644_/X sky130_fd_sc_hd__and2_1
X_6830__412 _6830__412/A vssd1 vssd1 vccd1 vccd1 _8005_/CLK sky130_fd_sc_hd__inv_2
X_4575_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4575_/X sky130_fd_sc_hd__buf_2
X_7363_ _7394_/A vssd1 vssd1 vccd1 vccd1 _7363_/X sky130_fd_sc_hd__buf_1
X_6314_ _7721_/Q _6265_/X _6307_/X _6313_/X vssd1 vssd1 vccd1 vccd1 _7721_/D sky130_fd_sc_hd__a211o_1
X_6245_ _6231_/X _6839_/C _6240_/Y _6243_/X _6244_/X vssd1 vssd1 vccd1 vccd1 _6245_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6176_ _7626_/A _7698_/Q _6180_/S vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5127_ _8190_/Q _8260_/Q _5171_/S vssd1 vssd1 vccd1 vccd1 _5127_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5058_ _4965_/A _5057_/X _5230_/A vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _4024_/S vssd1 vssd1 vccd1 vccd1 _4018_/S sky130_fd_sc_hd__buf_2
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6089__180 _6089__180/A vssd1 vssd1 vccd1 vccd1 _7649_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3242_ clkbuf_0__3242_/X vssd1 vssd1 vccd1 vccd1 _6601_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7039__71 _7041__73/A vssd1 vssd1 vccd1 vccd1 _8168_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3386_ clkbuf_0__3386_/X vssd1 vssd1 vccd1 vccd1 _6941__493/A sky130_fd_sc_hd__clkbuf_16
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4360_ _8134_/Q _4134_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4208_/X _8161_/Q _4297_/S vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__mux2_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6030_ _7678_/Q _6029_/X _7608_/A vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7981_ _7981_/CLK _7981_/D vssd1 vssd1 vccd1 vccd1 _7981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6932_ _6944_/A vssd1 vssd1 vccd1 vccd1 _6932_/X sky130_fd_sc_hd__buf_1
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5814_ _7867_/Q _7868_/Q _7865_/Q _7866_/Q vssd1 vssd1 vccd1 vccd1 _5817_/C sky130_fd_sc_hd__and4bb_4
XFILLER_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8453__228 vssd1 vssd1 vccd1 vccd1 _8453__228/HI versionID[2] sky130_fd_sc_hd__conb_1
XFILLER_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7060__88 _7061__89/A vssd1 vssd1 vccd1 vccd1 _8185_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5745_ _7764_/Q _5547_/A _5753_/S vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__mux2_1
X_5676_ _5676_/A vssd1 vssd1 vccd1 vccd1 _7795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7415_ _7416_/B _7416_/C _7593_/A vssd1 vssd1 vccd1 vccd1 _7415_/Y sky130_fd_sc_hd__a21oi_1
X_4627_ _4650_/S _4624_/X _4626_/X vssd1 vssd1 vccd1 vccd1 _4627_/X sky130_fd_sc_hd__a21o_1
X_8395_ _8399_/CLK _8395_/D vssd1 vssd1 vccd1 vccd1 _8395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4558_ _4682_/B vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7277_ _8236_/Q _7277_/B vssd1 vssd1 vccd1 vccd1 _7277_/X sky130_fd_sc_hd__or2_1
X_4489_ _5761_/A _4875_/A vssd1 vssd1 vccd1 vccd1 _4505_/S sky130_fd_sc_hd__or2_2
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6228_ _6289_/A vssd1 vssd1 vccd1 vccd1 _6228_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6159_ _7865_/Q _6157_/X _6152_/X _6154_/X _7689_/Q vssd1 vssd1 vccd1 vccd1 _7689_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6876__445 _6876__445/A vssd1 vssd1 vccd1 vccd1 _8040_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6837__418 _6837__418/A vssd1 vssd1 vccd1 vccd1 _8011_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput95 _5930_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_110_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6924__479 _6925__480/A vssd1 vssd1 vccd1 vccd1 _8076_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _8375_/Q _3837_/X _3862_/S vssd1 vssd1 vccd1 vccd1 _3861_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3583_ clkbuf_0__3583_/X vssd1 vssd1 vccd1 vccd1 _7300__125/A sky130_fd_sc_hd__clkbuf_16
X_3791_ _8001_/Q _3783_/Y _5249_/B _4950_/B vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_1_1_0__3360_ clkbuf_0__3360_/X vssd1 vssd1 vccd1 vccd1 _6833__415/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5530_ _5545_/S vssd1 vssd1 vccd1 vccd1 _5539_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_117_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5461_ _7907_/Q _4208_/A _5467_/S vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7200_ _7194_/X _7196_/X _7198_/X _7199_/Y _7219_/A vssd1 vssd1 vccd1 vccd1 _8213_/D
+ sky130_fd_sc_hd__a221oi_1
X_4412_ _4412_/A vssd1 vssd1 vccd1 vccd1 _8115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8180_ _8180_/CLK _8180_/D vssd1 vssd1 vccd1 vccd1 _8180_/Q sky130_fd_sc_hd__dfxtp_1
X_5392_ _5392_/A vssd1 vssd1 vccd1 vccd1 _7938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3190_ _6422_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3190_/X sky130_fd_sc_hd__clkbuf_16
X_7131_ _8214_/Q vssd1 vssd1 vccd1 vccd1 _7204_/A sky130_fd_sc_hd__clkbuf_2
X_4343_ _4343_/A vssd1 vssd1 vccd1 vccd1 _8141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4274_ _8168_/Q _4128_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__mux2_1
X_6013_ _7724_/Q input6/X _6025_/S vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7964_ _7964_/CLK _7964_/D vssd1 vssd1 vccd1 vccd1 _7964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7569__42 _7569__42/A vssd1 vssd1 vccd1 vccd1 _8381_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7331__150 _7331__150/A vssd1 vssd1 vccd1 vccd1 _8277_/CLK sky130_fd_sc_hd__inv_2
X_7895_ _7895_/CLK _7895_/D vssd1 vssd1 vccd1 vccd1 _7895_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2974_ _6083_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2974_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7033__66 _7035__68/A vssd1 vssd1 vccd1 vccd1 _8163_/CLK sky130_fd_sc_hd__inv_2
X_5728_ _5728_/A vssd1 vssd1 vccd1 vccd1 _7772_/D sky130_fd_sc_hd__clkbuf_1
X_3989_ _5511_/B _3989_/B vssd1 vssd1 vccd1 vccd1 _4005_/S sky130_fd_sc_hd__nor2_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5659_ _5555_/X _7802_/Q _5663_/S vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__mux2_1
X_8378_ _8378_/CLK _8378_/D vssd1 vssd1 vccd1 vccd1 _8378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3388_ _6950_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3388_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3208_ clkbuf_0__3208_/X vssd1 vssd1 vccd1 vccd1 _6574__290/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8345_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _5100_/A _5100_/B _7995_/Q vssd1 vssd1 vccd1 vccd1 _5126_/A sky130_fd_sc_hd__a21oi_1
X_7680_ _8348_/CLK _7680_/D vssd1 vssd1 vccd1 vccd1 _7680_/Q sky130_fd_sc_hd__dfxtp_1
X_6700_ _8340_/Q vssd1 vssd1 vccd1 vccd1 _6700_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3912_ _3912_/A vssd1 vssd1 vccd1 vccd1 _8321_/D sky130_fd_sc_hd__clkbuf_1
X_4892_ _4892_/A vssd1 vssd1 vccd1 vccd1 _8038_/D sky130_fd_sc_hd__clkbuf_1
X_3843_ _8000_/Q vssd1 vssd1 vccd1 vccd1 _4230_/C sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3412_ clkbuf_0__3412_/X vssd1 vssd1 vccd1 vccd1 _7071__97/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3343_ clkbuf_0__3343_/X vssd1 vssd1 vccd1 vccd1 _6773__380/A sky130_fd_sc_hd__clkbuf_4
X_6562_ _7864_/Q _5895_/A _6564_/S vssd1 vssd1 vccd1 vccd1 _6563_/A sky130_fd_sc_hd__mux2_1
X_3774_ _8000_/Q vssd1 vssd1 vccd1 vccd1 _4120_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_8301_ _8301_/CLK _8301_/D vssd1 vssd1 vccd1 vccd1 _8301_/Q sky130_fd_sc_hd__dfxtp_1
X_5513_ _7884_/Q _5025_/A _5521_/S vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__mux2_1
X_6415__205 _6415__205/A vssd1 vssd1 vccd1 vccd1 _7762_/CLK sky130_fd_sc_hd__inv_2
X_8232_ _8239_/CLK _8232_/D vssd1 vssd1 vccd1 vccd1 _8232_/Q sky130_fd_sc_hd__dfxtp_1
X_5444_ _5444_/A vssd1 vssd1 vccd1 vccd1 _7915_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3242_ _6588_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3242_/X sky130_fd_sc_hd__clkbuf_16
X_8163_ _8163_/CLK _8163_/D vssd1 vssd1 vccd1 vccd1 _8163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7114_ _7159_/A _7159_/B _7150_/D _7238_/A _7113_/Y vssd1 vssd1 vccd1 vccd1 _7115_/B
+ sky130_fd_sc_hd__a32o_1
X_5375_ _7948_/Q _4517_/X _5377_/S vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4326_ _4348_/S vssd1 vssd1 vccd1 vccd1 _4339_/S sky130_fd_sc_hd__clkbuf_4
X_8094_ _8094_/CLK _8094_/D vssd1 vssd1 vccd1 vccd1 _8094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4257_ _4257_/A vssd1 vssd1 vccd1 vccd1 _8176_/D sky130_fd_sc_hd__clkbuf_1
X_7045_ _7069_/A vssd1 vssd1 vccd1 vccd1 _7045_/X sky130_fd_sc_hd__buf_1
X_4188_ _8202_/Q _4044_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7947_ _7947_/CLK _7947_/D vssd1 vssd1 vccd1 vccd1 _7947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _7878_/CLK _7878_/D vssd1 vssd1 vccd1 vccd1 _7878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7563__37 _7564__38/A vssd1 vssd1 vccd1 vccd1 _8376_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6889__455 _6889__455/A vssd1 vssd1 vccd1 vccd1 _8050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5160_ _5103_/X _5158_/X _5159_/X vssd1 vssd1 vccd1 vccd1 _5161_/C sky130_fd_sc_hd__o21a_1
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5091_ _5084_/X _5086_/X _5089_/X _5124_/A _5095_/A vssd1 vssd1 vccd1 vccd1 _5091_/X
+ sky130_fd_sc_hd__o221a_1
X_4111_ _4111_/A vssd1 vssd1 vccd1 vccd1 _8261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4042_ _8273_/Q _3963_/X _4042_/S vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5993_ _7667_/Q _5991_/X _6006_/S vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__mux2_4
X_7801_ _7801_/CLK _7801_/D vssd1 vssd1 vccd1 vccd1 _7801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7732_ _8365_/CLK _7732_/D vssd1 vssd1 vccd1 vccd1 _7732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4944_ _4944_/A vssd1 vssd1 vccd1 vccd1 _8016_/D sky130_fd_sc_hd__clkbuf_1
X_7663_ _7697_/CLK _7663_/D vssd1 vssd1 vccd1 vccd1 _7663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4875_ _4875_/A _5725_/A vssd1 vssd1 vccd1 vccd1 _4891_/S sky130_fd_sc_hd__nor2_2
X_7594_ _7590_/X _7591_/Y _7593_/Y _6292_/X vssd1 vssd1 vccd1 vccd1 _8392_/D sky130_fd_sc_hd__a211oi_2
X_3826_ _8387_/Q _3825_/X _3832_/S vssd1 vssd1 vccd1 vccd1 _3827_/A sky130_fd_sc_hd__mux2_1
X_6545_ _6545_/A vssd1 vssd1 vccd1 vccd1 _7856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8215_ _8364_/CLK _8215_/D vssd1 vssd1 vccd1 vccd1 _8215_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3188_ clkbuf_0__3188_/X vssd1 vssd1 vccd1 vccd1 _6415__205/A sky130_fd_sc_hd__clkbuf_4
X_5427_ _7922_/Q _4514_/X _5431_/S vssd1 vssd1 vccd1 vccd1 _5428_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8146_ _8146_/CLK _8146_/D vssd1 vssd1 vccd1 vccd1 _8146_/Q sky130_fd_sc_hd__dfxtp_1
X_5358_ _3831_/X _7955_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_3 _6079_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _8153_/Q _4125_/X _4315_/S vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__mux2_1
X_8077_ _8077_/CLK _8077_/D vssd1 vssd1 vccd1 vccd1 _8077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5289_ _5288_/X _7982_/Q _5297_/S vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7344__160 _7344__160/A vssd1 vssd1 vccd1 vccd1 _8287_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3403_ clkbuf_0__3403_/X vssd1 vssd1 vccd1 vccd1 _7022__57/A sky130_fd_sc_hd__clkbuf_16
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _8018_/Q _7873_/Q _7777_/Q _7761_/Q _4582_/X _4580_/A vssd1 vssd1 vccd1 vccd1
+ _4660_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4591_ _8122_/Q _7892_/Q _7836_/Q _7796_/Q _4579_/A _4589_/X vssd1 vssd1 vccd1 vccd1
+ _4591_/X sky130_fd_sc_hd__mux4_1
X_6330_ _7726_/Q _6320_/X _6324_/X _6329_/X vssd1 vssd1 vccd1 vccd1 _7726_/D sky130_fd_sc_hd__a211o_1
X_6261_ _8059_/Q _6231_/A _6201_/X _6235_/X vssd1 vssd1 vccd1 vccd1 _6261_/X sky130_fd_sc_hd__a31o_1
X_6192_ _8236_/Q _8237_/Q _8238_/Q _8239_/Q _7258_/B _8230_/Q vssd1 vssd1 vccd1 vccd1
+ _6192_/X sky130_fd_sc_hd__mux4_1
X_8000_ _8000_/CLK _8000_/D vssd1 vssd1 vccd1 vccd1 _8000_/Q sky130_fd_sc_hd__dfxtp_1
X_5212_ _5197_/X _5211_/X _5271_/B vssd1 vssd1 vccd1 vccd1 _5212_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5143_ _8007_/Q _4956_/A _5031_/X _5142_/X _4953_/A vssd1 vssd1 vccd1 vccd1 _5143_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5074_ _3875_/X _5029_/X _5073_/X _5027_/X vssd1 vssd1 vccd1 vccd1 _8009_/D sky130_fd_sc_hd__o211a_1
X_6978__523 _6980__525/A vssd1 vssd1 vccd1 vccd1 _8120_/CLK sky130_fd_sc_hd__inv_2
X_4025_ _4025_/A vssd1 vssd1 vccd1 vccd1 _8281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8421__196 vssd1 vssd1 vccd1 vccd1 _8421__196/HI core0Index[3] sky130_fd_sc_hd__conb_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ _7662_/Q _5973_/X _5989_/S vssd1 vssd1 vccd1 vccd1 _5977_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7715_ _7991_/CLK _7715_/D vssd1 vssd1 vccd1 vccd1 _7715_/Q sky130_fd_sc_hd__dfxtp_1
X_7287__114 _7288__115/A vssd1 vssd1 vccd1 vccd1 _8241_/CLK sky130_fd_sc_hd__inv_2
X_4927_ _4927_/A vssd1 vssd1 vccd1 vccd1 _8023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _4854_/B _4858_/B _6801_/A vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__and3b_1
X_7646_ _7646_/CLK _7646_/D vssd1 vssd1 vccd1 vccd1 _7646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ _7750_/Q _7751_/Q _7752_/Q _7753_/Q vssd1 vssd1 vccd1 vccd1 _6341_/C sky130_fd_sc_hd__or4_2
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4789_ _4819_/A _4789_/B _4789_/C vssd1 vssd1 vccd1 vccd1 _4789_/X sky130_fd_sc_hd__or3_1
XFILLER_119_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _5862_/A _7849_/Q _6528_/S vssd1 vssd1 vccd1 vccd1 _6529_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6459_ _6465_/A vssd1 vssd1 vccd1 vccd1 _6459_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3208_ _6515_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3208_/X sky130_fd_sc_hd__clkbuf_16
X_8129_ _8129_/CLK _8129_/D vssd1 vssd1 vccd1 vccd1 _8129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5830_ _6536_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5831_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3591_ clkbuf_0__3591_/X vssd1 vssd1 vccd1 vccd1 _7338__155/A sky130_fd_sc_hd__clkbuf_4
X_7375__10 _7374__9/A vssd1 vssd1 vccd1 vccd1 _8312_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _5761_/A _5795_/B vssd1 vssd1 vccd1 vccd1 _5777_/S sky130_fd_sc_hd__or2_2
X_7500_ _7498_/A _7497_/Y _7499_/X _7448_/X vssd1 vssd1 vccd1 vccd1 _8347_/D sky130_fd_sc_hd__o211a_1
X_4712_ _8118_/Q _4681_/X _4664_/A _4711_/X vssd1 vssd1 vccd1 vccd1 _4712_/X sky130_fd_sc_hd__o211a_1
X_7431_ _7430_/B _7430_/C _7430_/A vssd1 vssd1 vccd1 vccd1 _7431_/Y sky130_fd_sc_hd__a21oi_1
X_5692_ _5692_/A vssd1 vssd1 vccd1 vccd1 _7788_/D sky130_fd_sc_hd__clkbuf_1
X_4643_ _8200_/Q _7818_/Q _7802_/Q _7786_/Q _4571_/A _4569_/X vssd1 vssd1 vccd1 vccd1
+ _4644_/B sky130_fd_sc_hd__mux4_1
X_4574_ _4601_/B _4584_/B vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__or2_2
X_6313_ _7612_/A _6326_/B _6322_/C _6326_/D vssd1 vssd1 vccd1 vccd1 _6313_/X sky130_fd_sc_hd__and4_1
X_6244_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6244_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6175_ _6175_/A vssd1 vssd1 vccd1 vccd1 _7697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5126_ _5126_/A vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5057_ _8278_/Q _8262_/Q _8192_/Q _8286_/Q _5231_/S _5010_/X vssd1 vssd1 vccd1 vccd1
+ _5057_/X sky130_fd_sc_hd__mux4_1
X_4008_ _5348_/A _4204_/B vssd1 vssd1 vccd1 vccd1 _4024_/S sky130_fd_sc_hd__or2_2
XFILLER_111_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5959_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6577__292 _6577__292/A vssd1 vssd1 vccd1 vccd1 _7873_/CLK sky130_fd_sc_hd__inv_2
X_7629_ _7629_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4290_ _4290_/A vssd1 vssd1 vccd1 vccd1 _8162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7980_ _7980_/CLK _7980_/D vssd1 vssd1 vccd1 vccd1 _7980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5813_ _6036_/A vssd1 vssd1 vccd1 vccd1 _6687_/A sky130_fd_sc_hd__buf_2
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5744_ _5759_/S vssd1 vssd1 vccd1 vccd1 _5753_/S sky130_fd_sc_hd__clkbuf_4
X_5675_ _7795_/Q _5578_/X _5681_/S vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7414_ _7167_/A _6699_/B _7412_/X _7413_/Y vssd1 vssd1 vccd1 vccd1 _7414_/X sky130_fd_sc_hd__o211a_1
X_8394_ _8407_/CLK _8394_/D vssd1 vssd1 vccd1 vccd1 _8394_/Q sky130_fd_sc_hd__dfxtp_2
X_4626_ _4593_/S _4625_/X _4802_/A vssd1 vssd1 vccd1 vccd1 _4626_/X sky130_fd_sc_hd__a21o_1
X_7345_ _7357_/A vssd1 vssd1 vccd1 vccd1 _7345_/X sky130_fd_sc_hd__buf_1
XFILLER_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4557_ _4557_/A vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7276_ _8007_/Q _7266_/X _7275_/X _7269_/X vssd1 vssd1 vccd1 vccd1 _8235_/D sky130_fd_sc_hd__o211a_1
X_4488_ _5653_/B vssd1 vssd1 vccd1 vccd1 _5761_/A sky130_fd_sc_hd__clkbuf_2
X_6227_ _6285_/A _6285_/B vssd1 vssd1 vccd1 vccd1 _6289_/A sky130_fd_sc_hd__or2_1
X_6158_ _7864_/Q _6157_/X _6152_/X _6154_/X _7688_/Q vssd1 vssd1 vccd1 vccd1 _7688_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _8102_/Q _5098_/X _5103_/X _5105_/X _5108_/X vssd1 vssd1 vccd1 vccd1 _5109_/X
+ sky130_fd_sc_hd__o221a_1
X_6464__245 _6464__245/A vssd1 vssd1 vccd1 vccd1 _7802_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_1_wb_clk_i clkbuf_opt_2_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput96 _5932_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__buf_2
XFILLER_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _3893_/A _4949_/A _4950_/C vssd1 vssd1 vccd1 vccd1 _3790_/Y sky130_fd_sc_hd__a21boi_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8413__235 vssd1 vssd1 vccd1 vccd1 partID[8] _8413__235/LO sky130_fd_sc_hd__conb_1
X_5460_ _5460_/A vssd1 vssd1 vccd1 vccd1 _7908_/D sky130_fd_sc_hd__clkbuf_1
X_6673__364 _6674__365/A vssd1 vssd1 vccd1 vccd1 _7948_/CLK sky130_fd_sc_hd__inv_2
X_6634__337 _6635__338/A vssd1 vssd1 vccd1 vccd1 _7918_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4411_ _8115_/Q _4410_/X _4411_/S vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _7938_/Q _4514_/X _5395_/S vssd1 vssd1 vccd1 vccd1 _5392_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7130_ _8403_/Q _7130_/B vssd1 vssd1 vccd1 vccd1 _7130_/X sky130_fd_sc_hd__xor2_1
X_4342_ _4341_/X _8141_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4343_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4273_ _4273_/A vssd1 vssd1 vccd1 vccd1 _8169_/D sky130_fd_sc_hd__clkbuf_1
X_6012_ _6029_/S vssd1 vssd1 vccd1 vccd1 _6025_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

