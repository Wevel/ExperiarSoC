magic
tech sky130A
magscale 1 2
timestamp 1653402413
<< viali >>
rect 2329 39593 2363 39627
rect 3065 39593 3099 39627
rect 3985 39593 4019 39627
rect 26433 39593 26467 39627
rect 41429 39593 41463 39627
rect 48973 39593 49007 39627
rect 56425 39593 56459 39627
rect 19257 39457 19291 39491
rect 1409 39389 1443 39423
rect 2145 39389 2179 39423
rect 2881 39389 2915 39423
rect 1593 39253 1627 39287
rect 1409 38913 1443 38947
rect 1593 38709 1627 38743
rect 1593 38505 1627 38539
rect 1409 38301 1443 38335
rect 1409 37825 1443 37859
rect 1593 37621 1627 37655
rect 1409 36737 1443 36771
rect 1593 36601 1627 36635
rect 1409 36125 1443 36159
rect 1593 35989 1627 36023
rect 1409 35037 1443 35071
rect 1593 34901 1627 34935
rect 1409 34697 1443 34731
rect 1593 34561 1627 34595
rect 1409 33949 1443 33983
rect 1593 33813 1627 33847
rect 1593 33473 1627 33507
rect 2421 33473 2455 33507
rect 1409 33337 1443 33371
rect 2237 33269 2271 33303
rect 3249 32997 3283 33031
rect 4997 32929 5031 32963
rect 5089 32929 5123 32963
rect 1869 32861 1903 32895
rect 2136 32793 2170 32827
rect 4537 32725 4571 32759
rect 4905 32725 4939 32759
rect 1593 32521 1627 32555
rect 2421 32521 2455 32555
rect 2881 32521 2915 32555
rect 5825 32521 5859 32555
rect 2789 32453 2823 32487
rect 1409 32385 1443 32419
rect 4712 32385 4746 32419
rect 3065 32317 3099 32351
rect 4445 32317 4479 32351
rect 4813 31977 4847 32011
rect 1409 31909 1443 31943
rect 1593 31773 1627 31807
rect 3065 31773 3099 31807
rect 4997 31773 5031 31807
rect 2881 31637 2915 31671
rect 3126 31365 3160 31399
rect 4721 31365 4755 31399
rect 1409 31297 1443 31331
rect 4905 31297 4939 31331
rect 4997 31297 5031 31331
rect 2881 31229 2915 31263
rect 1593 31161 1627 31195
rect 4261 31093 4295 31127
rect 4721 31093 4755 31127
rect 5181 31093 5215 31127
rect 2513 30889 2547 30923
rect 2973 30753 3007 30787
rect 3157 30753 3191 30787
rect 1593 30685 1627 30719
rect 2881 30685 2915 30719
rect 1409 30549 1443 30583
rect 4537 30345 4571 30379
rect 1409 30209 1443 30243
rect 2697 30209 2731 30243
rect 3413 30209 3447 30243
rect 3157 30141 3191 30175
rect 2513 30073 2547 30107
rect 1593 30005 1627 30039
rect 3801 29801 3835 29835
rect 4445 29665 4479 29699
rect 1593 29597 1627 29631
rect 4169 29597 4203 29631
rect 4261 29529 4295 29563
rect 1409 29461 1443 29495
rect 2881 29257 2915 29291
rect 1409 29121 1443 29155
rect 2789 29121 2823 29155
rect 2973 29053 3007 29087
rect 1593 28985 1627 29019
rect 2421 28917 2455 28951
rect 1869 28509 1903 28543
rect 2136 28441 2170 28475
rect 3249 28373 3283 28407
rect 2329 28169 2363 28203
rect 1593 28033 1627 28067
rect 2513 28033 2547 28067
rect 3893 28033 3927 28067
rect 3985 27965 4019 27999
rect 4077 27965 4111 27999
rect 1409 27829 1443 27863
rect 3525 27829 3559 27863
rect 2881 27625 2915 27659
rect 1409 27421 1443 27455
rect 2421 27421 2455 27455
rect 3065 27421 3099 27455
rect 4169 27421 4203 27455
rect 4414 27353 4448 27387
rect 1593 27285 1627 27319
rect 2237 27285 2271 27319
rect 5549 27285 5583 27319
rect 3985 27081 4019 27115
rect 2044 27013 2078 27047
rect 1777 26945 1811 26979
rect 4169 26945 4203 26979
rect 3157 26741 3191 26775
rect 2237 26537 2271 26571
rect 3801 26537 3835 26571
rect 4261 26469 4295 26503
rect 2697 26401 2731 26435
rect 2881 26401 2915 26435
rect 3893 26401 3927 26435
rect 1409 26333 1443 26367
rect 2605 26333 2639 26367
rect 4077 26333 4111 26367
rect 3801 26265 3835 26299
rect 1593 26197 1627 26231
rect 1593 25857 1627 25891
rect 3893 25857 3927 25891
rect 1409 25653 1443 25687
rect 3709 25653 3743 25687
rect 5181 25449 5215 25483
rect 1409 25245 1443 25279
rect 3801 25245 3835 25279
rect 4057 25245 4091 25279
rect 1593 25109 1627 25143
rect 3433 24905 3467 24939
rect 3801 24905 3835 24939
rect 1593 24769 1627 24803
rect 2421 24769 2455 24803
rect 3893 24769 3927 24803
rect 3985 24701 4019 24735
rect 1409 24633 1443 24667
rect 2237 24565 2271 24599
rect 1869 24157 1903 24191
rect 2136 24157 2170 24191
rect 3249 24021 3283 24055
rect 1593 23817 1627 23851
rect 2237 23817 2271 23851
rect 2697 23817 2731 23851
rect 2605 23749 2639 23783
rect 1409 23681 1443 23715
rect 3525 23681 3559 23715
rect 2789 23613 2823 23647
rect 3709 23613 3743 23647
rect 4537 23137 4571 23171
rect 1593 23069 1627 23103
rect 2237 23069 2271 23103
rect 4782 23001 4816 23035
rect 1409 22933 1443 22967
rect 2053 22933 2087 22967
rect 5917 22933 5951 22967
rect 3893 22729 3927 22763
rect 4629 22729 4663 22763
rect 3801 22661 3835 22695
rect 1409 22593 1443 22627
rect 2421 22593 2455 22627
rect 4813 22593 4847 22627
rect 3985 22525 4019 22559
rect 3433 22457 3467 22491
rect 1593 22389 1627 22423
rect 2237 22389 2271 22423
rect 3249 22185 3283 22219
rect 3801 22185 3835 22219
rect 4997 22185 5031 22219
rect 4261 22117 4295 22151
rect 1869 22049 1903 22083
rect 3985 22049 4019 22083
rect 4813 22049 4847 22083
rect 7021 22049 7055 22083
rect 2136 21981 2170 22015
rect 3801 21981 3835 22015
rect 4077 21981 4111 22015
rect 4721 21981 4755 22015
rect 4997 21981 5031 22015
rect 7288 21913 7322 21947
rect 5181 21845 5215 21879
rect 8401 21845 8435 21879
rect 2237 21641 2271 21675
rect 2605 21641 2639 21675
rect 8033 21641 8067 21675
rect 1409 21505 1443 21539
rect 2697 21505 2731 21539
rect 8217 21505 8251 21539
rect 8401 21505 8435 21539
rect 8493 21505 8527 21539
rect 9597 21505 9631 21539
rect 9864 21505 9898 21539
rect 2789 21437 2823 21471
rect 1593 21301 1627 21335
rect 10977 21301 11011 21335
rect 8217 21097 8251 21131
rect 9413 21097 9447 21131
rect 10425 21097 10459 21131
rect 13093 21097 13127 21131
rect 15761 21097 15795 21131
rect 4261 20961 4295 20995
rect 6193 20961 6227 20995
rect 8125 20961 8159 20995
rect 9505 20961 9539 20995
rect 1593 20893 1627 20927
rect 2421 20893 2455 20927
rect 4537 20893 4571 20927
rect 8033 20893 8067 20927
rect 9413 20893 9447 20927
rect 10609 20893 10643 20927
rect 10885 20893 10919 20927
rect 11713 20893 11747 20927
rect 14381 20893 14415 20927
rect 6460 20825 6494 20859
rect 11980 20825 12014 20859
rect 14648 20825 14682 20859
rect 1409 20757 1443 20791
rect 2237 20757 2271 20791
rect 7573 20757 7607 20791
rect 8401 20757 8435 20791
rect 9781 20757 9815 20791
rect 10793 20757 10827 20791
rect 3341 20553 3375 20587
rect 7297 20553 7331 20587
rect 7665 20553 7699 20587
rect 8585 20553 8619 20587
rect 12449 20553 12483 20587
rect 14657 20553 14691 20587
rect 2228 20485 2262 20519
rect 1961 20417 1995 20451
rect 7481 20417 7515 20451
rect 7757 20417 7791 20451
rect 8217 20417 8251 20451
rect 12633 20417 12667 20451
rect 12817 20417 12851 20451
rect 12909 20417 12943 20451
rect 14841 20417 14875 20451
rect 15025 20417 15059 20451
rect 15117 20417 15151 20451
rect 8309 20349 8343 20383
rect 8217 20213 8251 20247
rect 2237 20009 2271 20043
rect 7389 20009 7423 20043
rect 12541 20009 12575 20043
rect 12725 20009 12759 20043
rect 14657 20009 14691 20043
rect 15025 20009 15059 20043
rect 1593 19941 1627 19975
rect 2697 19873 2731 19907
rect 2789 19873 2823 19907
rect 1409 19805 1443 19839
rect 2605 19805 2639 19839
rect 7389 19805 7423 19839
rect 7481 19805 7515 19839
rect 12357 19805 12391 19839
rect 12541 19805 12575 19839
rect 14657 19805 14691 19839
rect 14841 19805 14875 19839
rect 7757 19669 7791 19703
rect 5365 19465 5399 19499
rect 7757 19465 7791 19499
rect 14841 19465 14875 19499
rect 15669 19465 15703 19499
rect 4252 19397 4286 19431
rect 1593 19329 1627 19363
rect 6561 19329 6595 19363
rect 7573 19329 7607 19363
rect 7849 19329 7883 19363
rect 9413 19329 9447 19363
rect 11805 19329 11839 19363
rect 12817 19329 12851 19363
rect 14473 19329 14507 19363
rect 15485 19329 15519 19363
rect 15761 19329 15795 19363
rect 3985 19261 4019 19295
rect 6653 19261 6687 19295
rect 7389 19261 7423 19295
rect 9137 19261 9171 19295
rect 11529 19261 11563 19295
rect 12909 19261 12943 19295
rect 14565 19261 14599 19295
rect 6929 19193 6963 19227
rect 1409 19125 1443 19159
rect 6745 19125 6779 19159
rect 12817 19125 12851 19159
rect 13185 19125 13219 19159
rect 14473 19125 14507 19159
rect 15301 19125 15335 19159
rect 5457 18921 5491 18955
rect 9045 18921 9079 18955
rect 12357 18921 12391 18955
rect 14289 18921 14323 18955
rect 16865 18921 16899 18955
rect 4077 18785 4111 18819
rect 10977 18785 11011 18819
rect 1409 18717 1443 18751
rect 2421 18717 2455 18751
rect 7573 18717 7607 18751
rect 7757 18717 7791 18751
rect 7849 18717 7883 18751
rect 9229 18717 9263 18751
rect 13001 18717 13035 18751
rect 13185 18717 13219 18751
rect 13277 18717 13311 18751
rect 14289 18717 14323 18751
rect 14473 18717 14507 18751
rect 15485 18717 15519 18751
rect 15741 18717 15775 18751
rect 4344 18649 4378 18683
rect 7389 18649 7423 18683
rect 11244 18649 11278 18683
rect 12817 18649 12851 18683
rect 1593 18581 1627 18615
rect 2237 18581 2271 18615
rect 14657 18581 14691 18615
rect 2237 18377 2271 18411
rect 2697 18377 2731 18411
rect 1593 18241 1627 18275
rect 2605 18241 2639 18275
rect 3525 18241 3559 18275
rect 8033 18241 8067 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 11805 18241 11839 18275
rect 13820 18241 13854 18275
rect 2789 18173 2823 18207
rect 7757 18173 7791 18207
rect 11529 18173 11563 18207
rect 13553 18173 13587 18207
rect 14933 18105 14967 18139
rect 1409 18037 1443 18071
rect 3801 18037 3835 18071
rect 7297 17833 7331 17867
rect 14381 17833 14415 17867
rect 1869 17629 1903 17663
rect 2136 17629 2170 17663
rect 5917 17629 5951 17663
rect 7941 17629 7975 17663
rect 8217 17629 8251 17663
rect 14565 17629 14599 17663
rect 14749 17629 14783 17663
rect 14841 17629 14875 17663
rect 16681 17629 16715 17663
rect 6184 17561 6218 17595
rect 7757 17561 7791 17595
rect 16948 17561 16982 17595
rect 3249 17493 3283 17527
rect 8125 17493 8159 17527
rect 18061 17493 18095 17527
rect 1593 17289 1627 17323
rect 7665 17289 7699 17323
rect 1409 17153 1443 17187
rect 7297 17153 7331 17187
rect 7389 17153 7423 17187
rect 9781 17153 9815 17187
rect 10241 17153 10275 17187
rect 17132 17153 17166 17187
rect 10333 17085 10367 17119
rect 16865 17085 16899 17119
rect 7481 16949 7515 16983
rect 9597 16949 9631 16983
rect 10333 16949 10367 16983
rect 10609 16949 10643 16983
rect 18245 16949 18279 16983
rect 7389 16745 7423 16779
rect 11529 16745 11563 16779
rect 16681 16745 16715 16779
rect 17325 16745 17359 16779
rect 18245 16745 18279 16779
rect 4077 16609 4111 16643
rect 7389 16609 7423 16643
rect 16589 16609 16623 16643
rect 18337 16609 18371 16643
rect 1409 16541 1443 16575
rect 2421 16541 2455 16575
rect 7297 16541 7331 16575
rect 9689 16541 9723 16575
rect 10149 16541 10183 16575
rect 12265 16541 12299 16575
rect 12449 16541 12483 16575
rect 12541 16541 12575 16575
rect 16497 16541 16531 16575
rect 17509 16541 17543 16575
rect 17785 16541 17819 16575
rect 18245 16541 18279 16575
rect 4344 16473 4378 16507
rect 10416 16473 10450 16507
rect 12081 16473 12115 16507
rect 1593 16405 1627 16439
rect 2237 16405 2271 16439
rect 5457 16405 5491 16439
rect 7665 16405 7699 16439
rect 9505 16405 9539 16439
rect 16865 16405 16899 16439
rect 17693 16405 17727 16439
rect 18613 16405 18647 16439
rect 7481 16201 7515 16235
rect 7849 16201 7883 16235
rect 14841 16201 14875 16235
rect 17233 16201 17267 16235
rect 17601 16201 17635 16235
rect 2298 16133 2332 16167
rect 1593 16065 1627 16099
rect 6653 16065 6687 16099
rect 6745 16065 6779 16099
rect 7665 16065 7699 16099
rect 7941 16065 7975 16099
rect 10333 16065 10367 16099
rect 11785 16065 11819 16099
rect 13728 16065 13762 16099
rect 15301 16065 15335 16099
rect 15485 16065 15519 16099
rect 15669 16065 15703 16099
rect 15761 16065 15795 16099
rect 17417 16065 17451 16099
rect 17693 16065 17727 16099
rect 2053 15997 2087 16031
rect 10425 15997 10459 16031
rect 11529 15997 11563 16031
rect 13461 15997 13495 16031
rect 1409 15861 1443 15895
rect 3433 15861 3467 15895
rect 6837 15861 6871 15895
rect 7021 15861 7055 15895
rect 10333 15861 10367 15895
rect 10701 15861 10735 15895
rect 12909 15861 12943 15895
rect 2145 15657 2179 15691
rect 6653 15657 6687 15691
rect 10793 15657 10827 15691
rect 14473 15657 14507 15691
rect 14841 15657 14875 15691
rect 17417 15657 17451 15691
rect 2605 15521 2639 15555
rect 2697 15521 2731 15555
rect 5273 15521 5307 15555
rect 14565 15521 14599 15555
rect 16957 15521 16991 15555
rect 1593 15453 1627 15487
rect 2513 15453 2547 15487
rect 7665 15453 7699 15487
rect 7849 15453 7883 15487
rect 7941 15453 7975 15487
rect 10977 15453 11011 15487
rect 11161 15453 11195 15487
rect 11253 15453 11287 15487
rect 14473 15453 14507 15487
rect 17233 15453 17267 15487
rect 17417 15453 17451 15487
rect 5540 15385 5574 15419
rect 7481 15385 7515 15419
rect 1409 15317 1443 15351
rect 17601 15317 17635 15351
rect 18613 15113 18647 15147
rect 8309 15045 8343 15079
rect 1409 14977 1443 15011
rect 2421 14977 2455 15011
rect 8125 14977 8159 15011
rect 10057 14977 10091 15011
rect 10241 14977 10275 15011
rect 10333 14977 10367 15011
rect 17500 14977 17534 15011
rect 13921 14909 13955 14943
rect 14197 14909 14231 14943
rect 17233 14909 17267 14943
rect 1593 14841 1627 14875
rect 2237 14773 2271 14807
rect 9873 14773 9907 14807
rect 1409 14569 1443 14603
rect 2329 14569 2363 14603
rect 4353 14569 4387 14603
rect 10333 14569 10367 14603
rect 10885 14569 10919 14603
rect 11253 14569 11287 14603
rect 16865 14569 16899 14603
rect 17509 14569 17543 14603
rect 13553 14501 13587 14535
rect 2789 14433 2823 14467
rect 2973 14433 3007 14467
rect 5825 14433 5859 14467
rect 5917 14433 5951 14467
rect 10977 14433 11011 14467
rect 1593 14365 1627 14399
rect 8953 14365 8987 14399
rect 9220 14365 9254 14399
rect 10885 14365 10919 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 16681 14365 16715 14399
rect 16865 14365 16899 14399
rect 17693 14365 17727 14399
rect 17877 14365 17911 14399
rect 17969 14365 18003 14399
rect 4261 14297 4295 14331
rect 13369 14297 13403 14331
rect 2697 14229 2731 14263
rect 5365 14229 5399 14263
rect 5733 14229 5767 14263
rect 17049 14229 17083 14263
rect 14105 14025 14139 14059
rect 18061 14025 18095 14059
rect 2228 13957 2262 13991
rect 3801 13889 3835 13923
rect 5733 13889 5767 13923
rect 12992 13889 13026 13923
rect 14657 13889 14691 13923
rect 14749 13889 14783 13923
rect 16681 13889 16715 13923
rect 16948 13889 16982 13923
rect 1961 13821 1995 13855
rect 10149 13821 10183 13855
rect 10425 13821 10459 13855
rect 12725 13821 12759 13855
rect 3341 13753 3375 13787
rect 3985 13685 4019 13719
rect 5549 13685 5583 13719
rect 14657 13685 14691 13719
rect 15025 13685 15059 13719
rect 1593 13481 1627 13515
rect 6837 13481 6871 13515
rect 9505 13481 9539 13515
rect 14105 13481 14139 13515
rect 16865 13481 16899 13515
rect 5457 13345 5491 13379
rect 10149 13345 10183 13379
rect 12725 13345 12759 13379
rect 1409 13277 1443 13311
rect 5713 13277 5747 13311
rect 9321 13277 9355 13311
rect 9505 13277 9539 13311
rect 10425 13277 10459 13311
rect 13001 13277 13035 13311
rect 14289 13277 14323 13311
rect 14565 13277 14599 13311
rect 17049 13277 17083 13311
rect 17233 13277 17267 13311
rect 17325 13277 17359 13311
rect 4261 13209 4295 13243
rect 14473 13209 14507 13243
rect 4353 13141 4387 13175
rect 9689 13141 9723 13175
rect 4537 12937 4571 12971
rect 6377 12937 6411 12971
rect 6837 12937 6871 12971
rect 10149 12937 10183 12971
rect 14565 12937 14599 12971
rect 18429 12937 18463 12971
rect 4629 12869 4663 12903
rect 1409 12801 1443 12835
rect 2421 12801 2455 12835
rect 3065 12801 3099 12835
rect 5825 12801 5859 12835
rect 6745 12801 6779 12835
rect 8769 12801 8803 12835
rect 9036 12801 9070 12835
rect 10793 12801 10827 12835
rect 13093 12801 13127 12835
rect 14473 12801 14507 12835
rect 15761 12801 15795 12835
rect 15853 12801 15887 12835
rect 17305 12801 17339 12835
rect 4813 12733 4847 12767
rect 6929 12733 6963 12767
rect 13369 12733 13403 12767
rect 17049 12733 17083 12767
rect 2881 12665 2915 12699
rect 1593 12597 1627 12631
rect 2237 12597 2271 12631
rect 4169 12597 4203 12631
rect 5641 12597 5675 12631
rect 10885 12597 10919 12631
rect 15761 12597 15795 12631
rect 16129 12597 16163 12631
rect 2237 12393 2271 12427
rect 10149 12393 10183 12427
rect 13093 12393 13127 12427
rect 14289 12393 14323 12427
rect 16957 12393 16991 12427
rect 2789 12257 2823 12291
rect 6285 12257 6319 12291
rect 14197 12257 14231 12291
rect 1593 12189 1627 12223
rect 4537 12189 4571 12223
rect 6541 12189 6575 12223
rect 10333 12189 10367 12223
rect 10517 12189 10551 12223
rect 10609 12189 10643 12223
rect 11713 12189 11747 12223
rect 14105 12189 14139 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 17417 12189 17451 12223
rect 2697 12121 2731 12155
rect 11980 12121 12014 12155
rect 1409 12053 1443 12087
rect 2605 12053 2639 12087
rect 4353 12053 4387 12087
rect 7665 12053 7699 12087
rect 14473 12053 14507 12087
rect 13277 11849 13311 11883
rect 13645 11849 13679 11883
rect 2136 11781 2170 11815
rect 4690 11781 4724 11815
rect 11989 11781 12023 11815
rect 1869 11713 1903 11747
rect 4445 11713 4479 11747
rect 8493 11713 8527 11747
rect 8677 11713 8711 11747
rect 13461 11713 13495 11747
rect 13737 11713 13771 11747
rect 15301 11713 15335 11747
rect 16957 11713 16991 11747
rect 17049 11713 17083 11747
rect 15393 11645 15427 11679
rect 12173 11577 12207 11611
rect 3249 11509 3283 11543
rect 5825 11509 5859 11543
rect 8861 11509 8895 11543
rect 15393 11509 15427 11543
rect 15669 11509 15703 11543
rect 16957 11509 16991 11543
rect 17325 11509 17359 11543
rect 12817 11305 12851 11339
rect 15945 11305 15979 11339
rect 18705 11305 18739 11339
rect 1593 11237 1627 11271
rect 8033 11169 8067 11203
rect 1409 11101 1443 11135
rect 8217 11101 8251 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 12633 11101 12667 11135
rect 12817 11101 12851 11135
rect 14565 11101 14599 11135
rect 17325 11101 17359 11135
rect 8401 11033 8435 11067
rect 9321 11033 9355 11067
rect 10149 11033 10183 11067
rect 14832 11033 14866 11067
rect 17592 11033 17626 11067
rect 13001 10965 13035 10999
rect 1409 10761 1443 10795
rect 3065 10761 3099 10795
rect 12909 10761 12943 10795
rect 15301 10761 15335 10795
rect 15669 10761 15703 10795
rect 17509 10761 17543 10795
rect 17877 10761 17911 10795
rect 1593 10625 1627 10659
rect 2973 10625 3007 10659
rect 8677 10625 8711 10659
rect 11529 10625 11563 10659
rect 11796 10625 11830 10659
rect 15485 10625 15519 10659
rect 15761 10625 15795 10659
rect 17693 10625 17727 10659
rect 17969 10625 18003 10659
rect 3157 10557 3191 10591
rect 8493 10557 8527 10591
rect 2605 10421 2639 10455
rect 8861 10421 8895 10455
rect 5273 10217 5307 10251
rect 5457 10217 5491 10251
rect 7941 10217 7975 10251
rect 12081 10217 12115 10251
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 2881 10013 2915 10047
rect 4997 10013 5031 10047
rect 5181 10013 5215 10047
rect 5273 10013 5307 10047
rect 6101 10013 6135 10047
rect 8125 10013 8159 10047
rect 12265 10013 12299 10047
rect 12541 10013 12575 10047
rect 6368 9945 6402 9979
rect 2697 9877 2731 9911
rect 7481 9877 7515 9911
rect 12449 9877 12483 9911
rect 6377 9673 6411 9707
rect 2780 9605 2814 9639
rect 15853 9605 15887 9639
rect 1409 9537 1443 9571
rect 6561 9537 6595 9571
rect 10057 9537 10091 9571
rect 15761 9537 15795 9571
rect 16937 9537 16971 9571
rect 2513 9469 2547 9503
rect 8493 9469 8527 9503
rect 8953 9469 8987 9503
rect 10333 9469 10367 9503
rect 15945 9469 15979 9503
rect 16681 9469 16715 9503
rect 8861 9401 8895 9435
rect 1593 9333 1627 9367
rect 3893 9333 3927 9367
rect 15393 9333 15427 9367
rect 18061 9333 18095 9367
rect 3157 9129 3191 9163
rect 6009 9129 6043 9163
rect 6193 9129 6227 9163
rect 11989 9129 12023 9163
rect 15945 9129 15979 9163
rect 1409 9061 1443 9095
rect 5641 9061 5675 9095
rect 19257 9061 19291 9095
rect 7573 8993 7607 9027
rect 9137 8993 9171 9027
rect 10057 8993 10091 9027
rect 10609 8993 10643 9027
rect 17693 8993 17727 9027
rect 1593 8925 1627 8959
rect 2237 8925 2271 8959
rect 3065 8925 3099 8959
rect 7849 8925 7883 8959
rect 9229 8925 9263 8959
rect 13369 8925 13403 8959
rect 16129 8925 16163 8959
rect 17877 8925 17911 8959
rect 18153 8925 18187 8959
rect 19441 8925 19475 8959
rect 19717 8925 19751 8959
rect 10876 8857 10910 8891
rect 2053 8789 2087 8823
rect 6009 8789 6043 8823
rect 13185 8789 13219 8823
rect 18061 8789 18095 8823
rect 19625 8789 19659 8823
rect 1777 8585 1811 8619
rect 11529 8585 11563 8619
rect 15669 8585 15703 8619
rect 16037 8585 16071 8619
rect 17049 8585 17083 8619
rect 20361 8585 20395 8619
rect 2666 8517 2700 8551
rect 6469 8517 6503 8551
rect 7757 8517 7791 8551
rect 8125 8517 8159 8551
rect 13338 8517 13372 8551
rect 16681 8517 16715 8551
rect 19809 8517 19843 8551
rect 20729 8517 20763 8551
rect 1961 8449 1995 8483
rect 2421 8449 2455 8483
rect 6377 8449 6411 8483
rect 7941 8449 7975 8483
rect 10149 8449 10183 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 13093 8449 13127 8483
rect 15853 8449 15887 8483
rect 16129 8449 16163 8483
rect 16865 8449 16899 8483
rect 17141 8449 17175 8483
rect 18153 8449 18187 8483
rect 18429 8449 18463 8483
rect 19625 8449 19659 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 20821 8449 20855 8483
rect 10425 8381 10459 8415
rect 19441 8313 19475 8347
rect 3801 8245 3835 8279
rect 14473 8245 14507 8279
rect 2513 8041 2547 8075
rect 8125 8041 8159 8075
rect 10793 8041 10827 8075
rect 11161 8041 11195 8075
rect 12817 8041 12851 8075
rect 19257 7973 19291 8007
rect 2973 7905 3007 7939
rect 3157 7905 3191 7939
rect 13277 7905 13311 7939
rect 13369 7905 13403 7939
rect 17877 7905 17911 7939
rect 1409 7837 1443 7871
rect 6745 7837 6779 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 14289 7837 14323 7871
rect 14565 7837 14599 7871
rect 17601 7837 17635 7871
rect 19441 7837 19475 7871
rect 19717 7837 19751 7871
rect 7012 7769 7046 7803
rect 14105 7769 14139 7803
rect 19625 7769 19659 7803
rect 1593 7701 1627 7735
rect 2881 7701 2915 7735
rect 13185 7701 13219 7735
rect 14473 7701 14507 7735
rect 2145 7497 2179 7531
rect 5181 7497 5215 7531
rect 7113 7497 7147 7531
rect 13185 7497 13219 7531
rect 13553 7497 13587 7531
rect 14105 7497 14139 7531
rect 15393 7497 15427 7531
rect 18797 7497 18831 7531
rect 2697 7429 2731 7463
rect 15025 7429 15059 7463
rect 2513 7361 2547 7395
rect 2605 7361 2639 7395
rect 4057 7361 4091 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6929 7361 6963 7395
rect 8585 7361 8619 7395
rect 8677 7361 8711 7395
rect 8861 7361 8895 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 13369 7361 13403 7395
rect 13645 7361 13679 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 14565 7361 14599 7395
rect 15209 7361 15243 7395
rect 15485 7361 15519 7395
rect 17417 7361 17451 7395
rect 18613 7361 18647 7395
rect 18889 7361 18923 7395
rect 1961 7293 1995 7327
rect 3801 7293 3835 7327
rect 6653 7293 6687 7327
rect 6745 7293 6779 7327
rect 17141 7293 17175 7327
rect 9229 7225 9263 7259
rect 18429 7225 18463 7259
rect 10517 7157 10551 7191
rect 10885 7157 10919 7191
rect 2881 6953 2915 6987
rect 6101 6953 6135 6987
rect 7389 6953 7423 6987
rect 7205 6817 7239 6851
rect 14289 6817 14323 6851
rect 14565 6817 14599 6851
rect 15853 6817 15887 6851
rect 17141 6817 17175 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 4537 6749 4571 6783
rect 4813 6749 4847 6783
rect 6009 6749 6043 6783
rect 7113 6749 7147 6783
rect 7297 6749 7331 6783
rect 7573 6749 7607 6783
rect 9321 6749 9355 6783
rect 9505 6749 9539 6783
rect 10057 6749 10091 6783
rect 16129 6749 16163 6783
rect 17417 6749 17451 6783
rect 2697 6681 2731 6715
rect 10324 6681 10358 6715
rect 2897 6613 2931 6647
rect 3065 6613 3099 6647
rect 6837 6613 6871 6647
rect 9413 6613 9447 6647
rect 11437 6613 11471 6647
rect 3341 6409 3375 6443
rect 7205 6409 7239 6443
rect 10425 6409 10459 6443
rect 10793 6409 10827 6443
rect 14473 6409 14507 6443
rect 14841 6409 14875 6443
rect 16865 6409 16899 6443
rect 2789 6341 2823 6375
rect 3709 6341 3743 6375
rect 7113 6341 7147 6375
rect 14197 6341 14231 6375
rect 17754 6341 17788 6375
rect 1409 6273 1443 6307
rect 2697 6273 2731 6307
rect 3525 6273 3559 6307
rect 3801 6273 3835 6307
rect 10609 6273 10643 6307
rect 10885 6273 10919 6307
rect 14657 6273 14691 6307
rect 14933 6273 14967 6307
rect 17049 6273 17083 6307
rect 17509 6205 17543 6239
rect 1593 6069 1627 6103
rect 18889 6069 18923 6103
rect 14289 5865 14323 5899
rect 15209 5865 15243 5899
rect 16405 5865 16439 5899
rect 17601 5797 17635 5831
rect 3065 5729 3099 5763
rect 16865 5729 16899 5763
rect 16957 5729 16991 5763
rect 1593 5661 1627 5695
rect 6561 5661 6595 5695
rect 6828 5661 6862 5695
rect 14473 5661 14507 5695
rect 14749 5661 14783 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 17785 5661 17819 5695
rect 18061 5661 18095 5695
rect 2881 5593 2915 5627
rect 17969 5593 18003 5627
rect 1409 5525 1443 5559
rect 2421 5525 2455 5559
rect 2789 5525 2823 5559
rect 7941 5525 7975 5559
rect 14657 5525 14691 5559
rect 15577 5525 15611 5559
rect 16773 5525 16807 5559
rect 3617 5321 3651 5355
rect 12909 5321 12943 5355
rect 14473 5321 14507 5355
rect 14841 5321 14875 5355
rect 16681 5321 16715 5355
rect 18613 5321 18647 5355
rect 18981 5253 19015 5287
rect 2237 5185 2271 5219
rect 2504 5185 2538 5219
rect 4261 5185 4295 5219
rect 4905 5185 4939 5219
rect 6561 5185 6595 5219
rect 9781 5185 9815 5219
rect 10609 5185 10643 5219
rect 10701 5185 10735 5219
rect 11785 5185 11819 5219
rect 14657 5185 14691 5219
rect 14933 5185 14967 5219
rect 16865 5185 16899 5219
rect 17049 5185 17083 5219
rect 17141 5185 17175 5219
rect 18797 5185 18831 5219
rect 19073 5185 19107 5219
rect 4721 5117 4755 5151
rect 6377 5117 6411 5151
rect 9873 5117 9907 5151
rect 11529 5117 11563 5151
rect 4077 5049 4111 5083
rect 1593 4981 1627 5015
rect 5089 4981 5123 5015
rect 6745 4981 6779 5015
rect 9965 4981 9999 5015
rect 10149 4981 10183 5015
rect 10609 4981 10643 5015
rect 10977 4981 11011 5015
rect 2421 4777 2455 4811
rect 4629 4777 4663 4811
rect 11161 4777 11195 4811
rect 15393 4777 15427 4811
rect 18245 4777 18279 4811
rect 3801 4641 3835 4675
rect 19257 4641 19291 4675
rect 1409 4573 1443 4607
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 6193 4573 6227 4607
rect 6377 4573 6411 4607
rect 8953 4573 8987 4607
rect 11345 4573 11379 4607
rect 11621 4573 11655 4607
rect 15577 4573 15611 4607
rect 15853 4573 15887 4607
rect 16313 4573 16347 4607
rect 16589 4573 16623 4607
rect 18429 4573 18463 4607
rect 18705 4573 18739 4607
rect 24593 4573 24627 4607
rect 9220 4505 9254 4539
rect 11529 4505 11563 4539
rect 1593 4437 1627 4471
rect 3065 4437 3099 4471
rect 4169 4437 4203 4471
rect 6561 4437 6595 4471
rect 10333 4437 10367 4471
rect 15761 4437 15795 4471
rect 18613 4437 18647 4471
rect 19487 4437 19521 4471
rect 24409 4437 24443 4471
rect 10149 4233 10183 4267
rect 2237 4165 2271 4199
rect 6745 4165 6779 4199
rect 19717 4165 19751 4199
rect 1409 4097 1443 4131
rect 3433 4097 3467 4131
rect 3617 4097 3651 4131
rect 3709 4097 3743 4131
rect 4353 4097 4387 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 6837 4097 6871 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 10241 4097 10275 4131
rect 16129 4097 16163 4131
rect 18429 4097 18463 4131
rect 18613 4097 18647 4131
rect 18797 4097 18831 4131
rect 18889 4097 18923 4131
rect 19349 4097 19383 4131
rect 19533 4097 19567 4131
rect 19809 4097 19843 4131
rect 6929 4029 6963 4063
rect 16681 4029 16715 4063
rect 16957 4029 16991 4063
rect 5457 3961 5491 3995
rect 1593 3893 1627 3927
rect 3249 3893 3283 3927
rect 4169 3893 4203 3927
rect 4813 3893 4847 3927
rect 6377 3893 6411 3927
rect 15945 3893 15979 3927
rect 5641 3689 5675 3723
rect 10701 3689 10735 3723
rect 16589 3689 16623 3723
rect 18245 3689 18279 3723
rect 5181 3621 5215 3655
rect 57989 3621 58023 3655
rect 3801 3553 3835 3587
rect 14657 3553 14691 3587
rect 1409 3485 1443 3519
rect 2145 3485 2179 3519
rect 2881 3485 2915 3519
rect 4057 3485 4091 3519
rect 5825 3485 5859 3519
rect 6469 3485 6503 3519
rect 7113 3485 7147 3519
rect 7757 3485 7791 3519
rect 10241 3485 10275 3519
rect 10885 3485 10919 3519
rect 11161 3485 11195 3519
rect 11805 3485 11839 3519
rect 13553 3485 13587 3519
rect 14933 3485 14967 3519
rect 16129 3485 16163 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 17785 3485 17819 3519
rect 18429 3485 18463 3519
rect 18705 3485 18739 3519
rect 19441 3485 19475 3519
rect 21373 3485 21407 3519
rect 57805 3417 57839 3451
rect 1593 3349 1627 3383
rect 2329 3349 2363 3383
rect 3065 3349 3099 3383
rect 6285 3349 6319 3383
rect 7573 3349 7607 3383
rect 10057 3349 10091 3383
rect 11069 3349 11103 3383
rect 13369 3349 13403 3383
rect 16957 3349 16991 3383
rect 18613 3349 18647 3383
rect 19257 3349 19291 3383
rect 21189 3349 21223 3383
rect 7941 3145 7975 3179
rect 10425 3145 10459 3179
rect 10793 3145 10827 3179
rect 11529 3145 11563 3179
rect 11897 3145 11931 3179
rect 14473 3145 14507 3179
rect 17141 3145 17175 3179
rect 23673 3145 23707 3179
rect 56977 3145 57011 3179
rect 6806 3077 6840 3111
rect 16773 3077 16807 3111
rect 17693 3077 17727 3111
rect 18061 3077 18095 3111
rect 1685 3009 1719 3043
rect 2697 3009 2731 3043
rect 3709 3009 3743 3043
rect 5733 3009 5767 3043
rect 6561 3009 6595 3043
rect 8585 3009 8619 3043
rect 9965 3009 9999 3043
rect 10609 3009 10643 3043
rect 10885 3009 10919 3043
rect 11713 3009 11747 3043
rect 11989 3009 12023 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 14933 3009 14967 3043
rect 16129 3009 16163 3043
rect 16957 3009 16991 3043
rect 17233 3009 17267 3043
rect 17877 3009 17911 3043
rect 18153 3009 18187 3043
rect 19073 3009 19107 3043
rect 21281 3009 21315 3043
rect 23857 3009 23891 3043
rect 27721 3009 27755 3043
rect 33701 3009 33735 3043
rect 56793 3009 56827 3043
rect 1409 2941 1443 2975
rect 4353 2941 4387 2975
rect 13185 2941 13219 2975
rect 13461 2941 13495 2975
rect 33425 2941 33459 2975
rect 4997 2873 5031 2907
rect 8401 2873 8435 2907
rect 15945 2873 15979 2907
rect 18889 2873 18923 2907
rect 21097 2873 21131 2907
rect 27537 2873 27571 2907
rect 2881 2805 2915 2839
rect 3525 2805 3559 2839
rect 5549 2805 5583 2839
rect 9229 2805 9263 2839
rect 9781 2805 9815 2839
rect 12633 2805 12667 2839
rect 19717 2805 19751 2839
rect 22017 2805 22051 2839
rect 32597 2805 32631 2839
rect 35541 2805 35575 2839
rect 37473 2805 37507 2839
rect 39957 2805 39991 2839
rect 42901 2805 42935 2839
rect 44373 2805 44407 2839
rect 47777 2805 47811 2839
rect 50169 2805 50203 2839
rect 53113 2805 53147 2839
rect 54585 2805 54619 2839
rect 58173 2805 58207 2839
rect 12541 2601 12575 2635
rect 26065 2601 26099 2635
rect 28825 2601 28859 2635
rect 30297 2601 30331 2635
rect 51181 2601 51215 2635
rect 14105 2533 14139 2567
rect 16865 2533 16899 2567
rect 48237 2533 48271 2567
rect 4537 2465 4571 2499
rect 7297 2465 7331 2499
rect 18245 2465 18279 2499
rect 32413 2465 32447 2499
rect 38117 2465 38151 2499
rect 1409 2397 1443 2431
rect 3801 2397 3835 2431
rect 6377 2397 6411 2431
rect 9045 2397 9079 2431
rect 9965 2397 9999 2431
rect 11805 2397 11839 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 14289 2397 14323 2431
rect 14933 2397 14967 2431
rect 17325 2397 17359 2431
rect 19809 2397 19843 2431
rect 20729 2397 20763 2431
rect 22201 2397 22235 2431
rect 23121 2397 23155 2431
rect 23857 2397 23891 2431
rect 24685 2397 24719 2431
rect 25605 2397 25639 2431
rect 26249 2397 26283 2431
rect 27169 2397 27203 2431
rect 28273 2397 28307 2431
rect 29009 2397 29043 2431
rect 29745 2397 29779 2431
rect 30481 2397 30515 2431
rect 31125 2397 31159 2431
rect 32137 2397 32171 2431
rect 34069 2397 34103 2431
rect 34897 2397 34931 2431
rect 35173 2397 35207 2431
rect 38761 2397 38795 2431
rect 41613 2397 41647 2431
rect 43637 2397 43671 2431
rect 45109 2397 45143 2431
rect 46029 2397 46063 2431
rect 46581 2397 46615 2431
rect 48053 2397 48087 2431
rect 48973 2397 49007 2431
rect 50169 2397 50203 2431
rect 50997 2397 51031 2431
rect 51917 2397 51951 2431
rect 52745 2397 52779 2431
rect 53941 2397 53975 2431
rect 55321 2397 55355 2431
rect 56241 2397 56275 2431
rect 58081 2397 58115 2431
rect 2605 2329 2639 2363
rect 12909 2329 12943 2363
rect 15669 2329 15703 2363
rect 36461 2329 36495 2363
rect 37933 2329 37967 2363
rect 39957 2329 39991 2363
rect 40785 2329 40819 2363
rect 42901 2329 42935 2363
rect 56977 2329 57011 2363
rect 3985 2261 4019 2295
rect 5181 2261 5215 2295
rect 6561 2261 6595 2295
rect 8033 2261 8067 2295
rect 9229 2261 9263 2295
rect 10793 2261 10827 2295
rect 11989 2261 12023 2295
rect 15117 2261 15151 2295
rect 17509 2261 17543 2295
rect 19993 2261 20027 2295
rect 22385 2261 22419 2295
rect 24869 2261 24903 2295
rect 36553 2261 36587 2295
rect 40049 2261 40083 2295
rect 40877 2261 40911 2295
rect 42993 2261 43027 2295
rect 43821 2261 43855 2295
rect 45293 2261 45327 2295
rect 46765 2261 46799 2295
rect 50353 2261 50387 2295
rect 52929 2261 52963 2295
rect 54125 2261 54159 2295
rect 55505 2261 55539 2295
rect 57069 2261 57103 2295
<< metal1 >>
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 2317 39627 2375 39633
rect 2317 39593 2329 39627
rect 2363 39624 2375 39627
rect 2774 39624 2780 39636
rect 2363 39596 2780 39624
rect 2363 39593 2375 39596
rect 2317 39587 2375 39593
rect 2774 39584 2780 39596
rect 2832 39584 2838 39636
rect 3050 39624 3056 39636
rect 3011 39596 3056 39624
rect 3050 39584 3056 39596
rect 3108 39584 3114 39636
rect 3694 39584 3700 39636
rect 3752 39624 3758 39636
rect 3973 39627 4031 39633
rect 3973 39624 3985 39627
rect 3752 39596 3985 39624
rect 3752 39584 3758 39596
rect 3973 39593 3985 39596
rect 4019 39593 4031 39627
rect 3973 39587 4031 39593
rect 26234 39584 26240 39636
rect 26292 39624 26298 39636
rect 26421 39627 26479 39633
rect 26421 39624 26433 39627
rect 26292 39596 26433 39624
rect 26292 39584 26298 39596
rect 26421 39593 26433 39596
rect 26467 39593 26479 39627
rect 41414 39624 41420 39636
rect 41375 39596 41420 39624
rect 26421 39587 26479 39593
rect 41414 39584 41420 39596
rect 41472 39584 41478 39636
rect 48682 39584 48688 39636
rect 48740 39624 48746 39636
rect 48961 39627 49019 39633
rect 48961 39624 48973 39627
rect 48740 39596 48973 39624
rect 48740 39584 48746 39596
rect 48961 39593 48973 39596
rect 49007 39593 49019 39627
rect 48961 39587 49019 39593
rect 56134 39584 56140 39636
rect 56192 39624 56198 39636
rect 56413 39627 56471 39633
rect 56413 39624 56425 39627
rect 56192 39596 56425 39624
rect 56192 39584 56198 39596
rect 56413 39593 56425 39596
rect 56459 39593 56471 39627
rect 56413 39587 56471 39593
rect 18690 39448 18696 39500
rect 18748 39488 18754 39500
rect 19245 39491 19303 39497
rect 19245 39488 19257 39491
rect 18748 39460 19257 39488
rect 18748 39448 18754 39460
rect 19245 39457 19257 39460
rect 19291 39457 19303 39491
rect 19245 39451 19303 39457
rect 1397 39423 1455 39429
rect 1397 39389 1409 39423
rect 1443 39389 1455 39423
rect 2130 39420 2136 39432
rect 2091 39392 2136 39420
rect 1397 39383 1455 39389
rect 1412 39352 1440 39383
rect 2130 39380 2136 39392
rect 2188 39380 2194 39432
rect 2869 39423 2927 39429
rect 2869 39389 2881 39423
rect 2915 39420 2927 39423
rect 9490 39420 9496 39432
rect 2915 39392 9496 39420
rect 2915 39389 2927 39392
rect 2869 39383 2927 39389
rect 9490 39380 9496 39392
rect 9548 39380 9554 39432
rect 6638 39352 6644 39364
rect 1412 39324 6644 39352
rect 6638 39312 6644 39324
rect 6696 39312 6702 39364
rect 1578 39284 1584 39296
rect 1539 39256 1584 39284
rect 1578 39244 1584 39256
rect 1636 39244 1642 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1397 38947 1455 38953
rect 1397 38913 1409 38947
rect 1443 38944 1455 38947
rect 2590 38944 2596 38956
rect 1443 38916 2596 38944
rect 1443 38913 1455 38916
rect 1397 38907 1455 38913
rect 2590 38904 2596 38916
rect 2648 38904 2654 38956
rect 1578 38740 1584 38752
rect 1539 38712 1584 38740
rect 1578 38700 1584 38712
rect 1636 38700 1642 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1581 38539 1639 38545
rect 1581 38505 1593 38539
rect 1627 38536 1639 38539
rect 2866 38536 2872 38548
rect 1627 38508 2872 38536
rect 1627 38505 1639 38508
rect 1581 38499 1639 38505
rect 2866 38496 2872 38508
rect 2924 38496 2930 38548
rect 1397 38335 1455 38341
rect 1397 38301 1409 38335
rect 1443 38332 1455 38335
rect 1486 38332 1492 38344
rect 1443 38304 1492 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 1486 38292 1492 38304
rect 1544 38292 1550 38344
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1394 37856 1400 37868
rect 1355 37828 1400 37856
rect 1394 37816 1400 37828
rect 1452 37816 1458 37868
rect 1578 37652 1584 37664
rect 1539 37624 1584 37652
rect 1578 37612 1584 37624
rect 1636 37612 1642 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1762 36768 1768 36780
rect 1443 36740 1768 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 1578 36632 1584 36644
rect 1539 36604 1584 36632
rect 1578 36592 1584 36604
rect 1636 36592 1642 36644
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1397 36159 1455 36165
rect 1397 36125 1409 36159
rect 1443 36156 1455 36159
rect 1670 36156 1676 36168
rect 1443 36128 1676 36156
rect 1443 36125 1455 36128
rect 1397 36119 1455 36125
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 1578 36020 1584 36032
rect 1539 35992 1584 36020
rect 1578 35980 1584 35992
rect 1636 35980 1642 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 5442 35068 5448 35080
rect 1443 35040 5448 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 5442 35028 5448 35040
rect 5500 35028 5506 35080
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1397 34731 1455 34737
rect 1397 34697 1409 34731
rect 1443 34728 1455 34731
rect 2866 34728 2872 34740
rect 1443 34700 2872 34728
rect 1443 34697 1455 34700
rect 1397 34691 1455 34697
rect 2866 34688 2872 34700
rect 2924 34688 2930 34740
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1397 33983 1455 33989
rect 1397 33949 1409 33983
rect 1443 33980 1455 33983
rect 2038 33980 2044 33992
rect 1443 33952 2044 33980
rect 1443 33949 1455 33952
rect 1397 33943 1455 33949
rect 2038 33940 2044 33952
rect 2096 33940 2102 33992
rect 1578 33844 1584 33856
rect 1539 33816 1584 33844
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1578 33504 1584 33516
rect 1539 33476 1584 33504
rect 1578 33464 1584 33476
rect 1636 33464 1642 33516
rect 2406 33504 2412 33516
rect 2367 33476 2412 33504
rect 2406 33464 2412 33476
rect 2464 33464 2470 33516
rect 1397 33371 1455 33377
rect 1397 33337 1409 33371
rect 1443 33368 1455 33371
rect 4982 33368 4988 33380
rect 1443 33340 4988 33368
rect 1443 33337 1455 33340
rect 1397 33331 1455 33337
rect 4982 33328 4988 33340
rect 5040 33328 5046 33380
rect 2222 33300 2228 33312
rect 2183 33272 2228 33300
rect 2222 33260 2228 33272
rect 2280 33260 2286 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 3237 33031 3295 33037
rect 3237 32997 3249 33031
rect 3283 33028 3295 33031
rect 4614 33028 4620 33040
rect 3283 33000 4620 33028
rect 3283 32997 3295 33000
rect 3237 32991 3295 32997
rect 4614 32988 4620 33000
rect 4672 32988 4678 33040
rect 4982 32960 4988 32972
rect 4943 32932 4988 32960
rect 4982 32920 4988 32932
rect 5040 32920 5046 32972
rect 5074 32920 5080 32972
rect 5132 32960 5138 32972
rect 5132 32932 5177 32960
rect 5132 32920 5138 32932
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32892 1915 32895
rect 1903 32864 2820 32892
rect 1903 32861 1915 32864
rect 1857 32855 1915 32861
rect 2792 32836 2820 32864
rect 2124 32827 2182 32833
rect 2124 32793 2136 32827
rect 2170 32824 2182 32827
rect 2222 32824 2228 32836
rect 2170 32796 2228 32824
rect 2170 32793 2182 32796
rect 2124 32787 2182 32793
rect 2222 32784 2228 32796
rect 2280 32784 2286 32836
rect 2774 32784 2780 32836
rect 2832 32784 2838 32836
rect 4525 32759 4583 32765
rect 4525 32725 4537 32759
rect 4571 32756 4583 32759
rect 4798 32756 4804 32768
rect 4571 32728 4804 32756
rect 4571 32725 4583 32728
rect 4525 32719 4583 32725
rect 4798 32716 4804 32728
rect 4856 32716 4862 32768
rect 4890 32716 4896 32768
rect 4948 32756 4954 32768
rect 4948 32728 4993 32756
rect 4948 32716 4954 32728
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1578 32552 1584 32564
rect 1539 32524 1584 32552
rect 1578 32512 1584 32524
rect 1636 32512 1642 32564
rect 2406 32552 2412 32564
rect 2367 32524 2412 32552
rect 2406 32512 2412 32524
rect 2464 32512 2470 32564
rect 2866 32552 2872 32564
rect 2827 32524 2872 32552
rect 2866 32512 2872 32524
rect 2924 32512 2930 32564
rect 4890 32512 4896 32564
rect 4948 32552 4954 32564
rect 5813 32555 5871 32561
rect 5813 32552 5825 32555
rect 4948 32524 5825 32552
rect 4948 32512 4954 32524
rect 5813 32521 5825 32524
rect 5859 32521 5871 32555
rect 5813 32515 5871 32521
rect 2777 32487 2835 32493
rect 2777 32453 2789 32487
rect 2823 32484 2835 32487
rect 4614 32484 4620 32496
rect 2823 32456 4620 32484
rect 2823 32453 2835 32456
rect 2777 32447 2835 32453
rect 4614 32444 4620 32456
rect 4672 32444 4678 32496
rect 1397 32419 1455 32425
rect 1397 32385 1409 32419
rect 1443 32416 1455 32419
rect 3326 32416 3332 32428
rect 1443 32388 3332 32416
rect 1443 32385 1455 32388
rect 1397 32379 1455 32385
rect 3326 32376 3332 32388
rect 3384 32376 3390 32428
rect 4706 32425 4712 32428
rect 4700 32379 4712 32425
rect 4764 32416 4770 32428
rect 4764 32388 4800 32416
rect 4706 32376 4712 32379
rect 4764 32376 4770 32388
rect 3053 32351 3111 32357
rect 3053 32317 3065 32351
rect 3099 32348 3111 32351
rect 3142 32348 3148 32360
rect 3099 32320 3148 32348
rect 3099 32317 3111 32320
rect 3053 32311 3111 32317
rect 3142 32308 3148 32320
rect 3200 32308 3206 32360
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32317 4491 32351
rect 4433 32311 4491 32317
rect 2774 32240 2780 32292
rect 2832 32280 2838 32292
rect 4448 32280 4476 32311
rect 2832 32252 4476 32280
rect 2832 32240 2838 32252
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 4706 31968 4712 32020
rect 4764 32008 4770 32020
rect 4801 32011 4859 32017
rect 4801 32008 4813 32011
rect 4764 31980 4813 32008
rect 4764 31968 4770 31980
rect 4801 31977 4813 31980
rect 4847 31977 4859 32011
rect 4801 31971 4859 31977
rect 1397 31943 1455 31949
rect 1397 31909 1409 31943
rect 1443 31940 1455 31943
rect 2958 31940 2964 31952
rect 1443 31912 2964 31940
rect 1443 31909 1455 31912
rect 1397 31903 1455 31909
rect 2958 31900 2964 31912
rect 3016 31900 3022 31952
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 3050 31804 3056 31816
rect 3011 31776 3056 31804
rect 3050 31764 3056 31776
rect 3108 31764 3114 31816
rect 4798 31764 4804 31816
rect 4856 31804 4862 31816
rect 4985 31807 5043 31813
rect 4985 31804 4997 31807
rect 4856 31776 4997 31804
rect 4856 31764 4862 31776
rect 4985 31773 4997 31776
rect 5031 31773 5043 31807
rect 4985 31767 5043 31773
rect 2866 31668 2872 31680
rect 2827 31640 2872 31668
rect 2866 31628 2872 31640
rect 2924 31628 2930 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 2866 31356 2872 31408
rect 2924 31396 2930 31408
rect 3114 31399 3172 31405
rect 3114 31396 3126 31399
rect 2924 31368 3126 31396
rect 2924 31356 2930 31368
rect 3114 31365 3126 31368
rect 3160 31365 3172 31399
rect 3114 31359 3172 31365
rect 4614 31356 4620 31408
rect 4672 31396 4678 31408
rect 4709 31399 4767 31405
rect 4709 31396 4721 31399
rect 4672 31368 4721 31396
rect 4672 31356 4678 31368
rect 4709 31365 4721 31368
rect 4755 31365 4767 31399
rect 4709 31359 4767 31365
rect 1397 31331 1455 31337
rect 1397 31297 1409 31331
rect 1443 31328 1455 31331
rect 3694 31328 3700 31340
rect 1443 31300 3700 31328
rect 1443 31297 1455 31300
rect 1397 31291 1455 31297
rect 3694 31288 3700 31300
rect 3752 31288 3758 31340
rect 4890 31328 4896 31340
rect 4851 31300 4896 31328
rect 4890 31288 4896 31300
rect 4948 31288 4954 31340
rect 4982 31288 4988 31340
rect 5040 31328 5046 31340
rect 5040 31300 5085 31328
rect 5040 31288 5046 31300
rect 2774 31220 2780 31272
rect 2832 31260 2838 31272
rect 2869 31263 2927 31269
rect 2869 31260 2881 31263
rect 2832 31232 2881 31260
rect 2832 31220 2838 31232
rect 2869 31229 2881 31232
rect 2915 31229 2927 31263
rect 2869 31223 2927 31229
rect 1578 31192 1584 31204
rect 1539 31164 1584 31192
rect 1578 31152 1584 31164
rect 1636 31152 1642 31204
rect 1394 31084 1400 31136
rect 1452 31124 1458 31136
rect 1854 31124 1860 31136
rect 1452 31096 1860 31124
rect 1452 31084 1458 31096
rect 1854 31084 1860 31096
rect 1912 31084 1918 31136
rect 2866 31084 2872 31136
rect 2924 31124 2930 31136
rect 4249 31127 4307 31133
rect 4249 31124 4261 31127
rect 2924 31096 4261 31124
rect 2924 31084 2930 31096
rect 4249 31093 4261 31096
rect 4295 31124 4307 31127
rect 4709 31127 4767 31133
rect 4709 31124 4721 31127
rect 4295 31096 4721 31124
rect 4295 31093 4307 31096
rect 4249 31087 4307 31093
rect 4709 31093 4721 31096
rect 4755 31093 4767 31127
rect 4709 31087 4767 31093
rect 4798 31084 4804 31136
rect 4856 31124 4862 31136
rect 5169 31127 5227 31133
rect 5169 31124 5181 31127
rect 4856 31096 5181 31124
rect 4856 31084 4862 31096
rect 5169 31093 5181 31096
rect 5215 31093 5227 31127
rect 5169 31087 5227 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 2501 30923 2559 30929
rect 2501 30889 2513 30923
rect 2547 30920 2559 30923
rect 3050 30920 3056 30932
rect 2547 30892 3056 30920
rect 2547 30889 2559 30892
rect 2501 30883 2559 30889
rect 3050 30880 3056 30892
rect 3108 30880 3114 30932
rect 2958 30784 2964 30796
rect 2919 30756 2964 30784
rect 2958 30744 2964 30756
rect 3016 30744 3022 30796
rect 3142 30744 3148 30796
rect 3200 30784 3206 30796
rect 4706 30784 4712 30796
rect 3200 30756 4712 30784
rect 3200 30744 3206 30756
rect 4706 30744 4712 30756
rect 4764 30784 4770 30796
rect 5074 30784 5080 30796
rect 4764 30756 5080 30784
rect 4764 30744 4770 30756
rect 5074 30744 5080 30756
rect 5132 30744 5138 30796
rect 1578 30716 1584 30728
rect 1539 30688 1584 30716
rect 1578 30676 1584 30688
rect 1636 30676 1642 30728
rect 2866 30716 2872 30728
rect 2827 30688 2872 30716
rect 2866 30676 2872 30688
rect 2924 30676 2930 30728
rect 1397 30583 1455 30589
rect 1397 30549 1409 30583
rect 1443 30580 1455 30583
rect 4614 30580 4620 30592
rect 1443 30552 4620 30580
rect 1443 30549 1455 30552
rect 1397 30543 1455 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 4525 30379 4583 30385
rect 4525 30345 4537 30379
rect 4571 30376 4583 30379
rect 4982 30376 4988 30388
rect 4571 30348 4988 30376
rect 4571 30345 4583 30348
rect 4525 30339 4583 30345
rect 4982 30336 4988 30348
rect 5040 30336 5046 30388
rect 7558 30308 7564 30320
rect 1412 30280 7564 30308
rect 1412 30249 1440 30280
rect 7558 30268 7564 30280
rect 7616 30268 7622 30320
rect 1397 30243 1455 30249
rect 1397 30209 1409 30243
rect 1443 30209 1455 30243
rect 2682 30240 2688 30252
rect 2643 30212 2688 30240
rect 1397 30203 1455 30209
rect 2682 30200 2688 30212
rect 2740 30200 2746 30252
rect 3401 30243 3459 30249
rect 3401 30240 3413 30243
rect 2976 30212 3413 30240
rect 2976 30172 3004 30212
rect 3401 30209 3413 30212
rect 3447 30209 3459 30243
rect 3401 30203 3459 30209
rect 2516 30144 3004 30172
rect 3145 30175 3203 30181
rect 2516 30113 2544 30144
rect 3145 30141 3157 30175
rect 3191 30141 3203 30175
rect 3145 30135 3203 30141
rect 2501 30107 2559 30113
rect 2501 30073 2513 30107
rect 2547 30073 2559 30107
rect 2501 30067 2559 30073
rect 2774 30064 2780 30116
rect 2832 30104 2838 30116
rect 3160 30104 3188 30135
rect 2832 30076 3188 30104
rect 2832 30064 2838 30076
rect 1578 30036 1584 30048
rect 1539 30008 1584 30036
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 2682 29792 2688 29844
rect 2740 29832 2746 29844
rect 3789 29835 3847 29841
rect 3789 29832 3801 29835
rect 2740 29804 3801 29832
rect 2740 29792 2746 29804
rect 3789 29801 3801 29804
rect 3835 29801 3847 29835
rect 3789 29795 3847 29801
rect 4433 29699 4491 29705
rect 4433 29665 4445 29699
rect 4479 29696 4491 29699
rect 4706 29696 4712 29708
rect 4479 29668 4712 29696
rect 4479 29665 4491 29668
rect 4433 29659 4491 29665
rect 4706 29656 4712 29668
rect 4764 29656 4770 29708
rect 1578 29628 1584 29640
rect 1539 29600 1584 29628
rect 1578 29588 1584 29600
rect 1636 29588 1642 29640
rect 4157 29631 4215 29637
rect 4157 29597 4169 29631
rect 4203 29628 4215 29631
rect 4982 29628 4988 29640
rect 4203 29600 4988 29628
rect 4203 29597 4215 29600
rect 4157 29591 4215 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 4249 29563 4307 29569
rect 4249 29529 4261 29563
rect 4295 29560 4307 29563
rect 4614 29560 4620 29572
rect 4295 29532 4620 29560
rect 4295 29529 4307 29532
rect 4249 29523 4307 29529
rect 4614 29520 4620 29532
rect 4672 29520 4678 29572
rect 1397 29495 1455 29501
rect 1397 29461 1409 29495
rect 1443 29492 1455 29495
rect 2866 29492 2872 29504
rect 1443 29464 2872 29492
rect 1443 29461 1455 29464
rect 1397 29455 1455 29461
rect 2866 29452 2872 29464
rect 2924 29452 2930 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 2866 29288 2872 29300
rect 2827 29260 2872 29288
rect 2866 29248 2872 29260
rect 2924 29248 2930 29300
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29152 1455 29155
rect 2406 29152 2412 29164
rect 1443 29124 2412 29152
rect 1443 29121 1455 29124
rect 1397 29115 1455 29121
rect 2406 29112 2412 29124
rect 2464 29112 2470 29164
rect 2774 29152 2780 29164
rect 2735 29124 2780 29152
rect 2774 29112 2780 29124
rect 2832 29112 2838 29164
rect 2222 29044 2228 29096
rect 2280 29084 2286 29096
rect 2961 29087 3019 29093
rect 2961 29084 2973 29087
rect 2280 29056 2973 29084
rect 2280 29044 2286 29056
rect 2961 29053 2973 29056
rect 3007 29053 3019 29087
rect 2961 29047 3019 29053
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 2409 28951 2467 28957
rect 2409 28917 2421 28951
rect 2455 28948 2467 28951
rect 2498 28948 2504 28960
rect 2455 28920 2504 28948
rect 2455 28917 2467 28920
rect 2409 28911 2467 28917
rect 2498 28908 2504 28920
rect 2556 28908 2562 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1857 28543 1915 28549
rect 1857 28509 1869 28543
rect 1903 28540 1915 28543
rect 2682 28540 2688 28552
rect 1903 28512 2688 28540
rect 1903 28509 1915 28512
rect 1857 28503 1915 28509
rect 2682 28500 2688 28512
rect 2740 28500 2746 28552
rect 2124 28475 2182 28481
rect 2124 28441 2136 28475
rect 2170 28472 2182 28475
rect 2314 28472 2320 28484
rect 2170 28444 2320 28472
rect 2170 28441 2182 28444
rect 2124 28435 2182 28441
rect 2314 28432 2320 28444
rect 2372 28432 2378 28484
rect 2774 28364 2780 28416
rect 2832 28404 2838 28416
rect 3237 28407 3295 28413
rect 3237 28404 3249 28407
rect 2832 28376 3249 28404
rect 2832 28364 2838 28376
rect 3237 28373 3249 28376
rect 3283 28404 3295 28407
rect 3786 28404 3792 28416
rect 3283 28376 3792 28404
rect 3283 28373 3295 28376
rect 3237 28367 3295 28373
rect 3786 28364 3792 28376
rect 3844 28364 3850 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 2314 28200 2320 28212
rect 2275 28172 2320 28200
rect 2314 28160 2320 28172
rect 2372 28160 2378 28212
rect 1394 28024 1400 28076
rect 1452 28064 1458 28076
rect 1581 28067 1639 28073
rect 1581 28064 1593 28067
rect 1452 28036 1593 28064
rect 1452 28024 1458 28036
rect 1581 28033 1593 28036
rect 1627 28033 1639 28067
rect 2498 28064 2504 28076
rect 2459 28036 2504 28064
rect 1581 28027 1639 28033
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 3878 28064 3884 28076
rect 3839 28036 3884 28064
rect 3878 28024 3884 28036
rect 3936 28024 3942 28076
rect 3970 27996 3976 28008
rect 3931 27968 3976 27996
rect 3970 27956 3976 27968
rect 4028 27956 4034 28008
rect 4065 27999 4123 28005
rect 4065 27965 4077 27999
rect 4111 27965 4123 27999
rect 4065 27959 4123 27965
rect 2314 27888 2320 27940
rect 2372 27928 2378 27940
rect 4080 27928 4108 27959
rect 2372 27900 4108 27928
rect 2372 27888 2378 27900
rect 1397 27863 1455 27869
rect 1397 27829 1409 27863
rect 1443 27860 1455 27863
rect 2682 27860 2688 27872
rect 1443 27832 2688 27860
rect 1443 27829 1455 27832
rect 1397 27823 1455 27829
rect 2682 27820 2688 27832
rect 2740 27820 2746 27872
rect 3513 27863 3571 27869
rect 3513 27829 3525 27863
rect 3559 27860 3571 27863
rect 4062 27860 4068 27872
rect 3559 27832 4068 27860
rect 3559 27829 3571 27832
rect 3513 27823 3571 27829
rect 4062 27820 4068 27832
rect 4120 27820 4126 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 2869 27659 2927 27665
rect 2869 27625 2881 27659
rect 2915 27656 2927 27659
rect 3970 27656 3976 27668
rect 2915 27628 3976 27656
rect 2915 27625 2927 27628
rect 2869 27619 2927 27625
rect 3970 27616 3976 27628
rect 4028 27616 4034 27668
rect 1412 27492 4292 27520
rect 1412 27461 1440 27492
rect 1397 27455 1455 27461
rect 1397 27421 1409 27455
rect 1443 27421 1455 27455
rect 2406 27452 2412 27464
rect 2367 27424 2412 27452
rect 1397 27415 1455 27421
rect 2406 27412 2412 27424
rect 2464 27412 2470 27464
rect 3050 27452 3056 27464
rect 3011 27424 3056 27452
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 4157 27455 4215 27461
rect 4157 27452 4169 27455
rect 3160 27424 4169 27452
rect 2774 27344 2780 27396
rect 2832 27384 2838 27396
rect 3160 27384 3188 27424
rect 4157 27421 4169 27424
rect 4203 27421 4215 27455
rect 4264 27452 4292 27492
rect 13078 27452 13084 27464
rect 4264 27424 13084 27452
rect 4157 27415 4215 27421
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 2832 27356 3188 27384
rect 2832 27344 2838 27356
rect 3970 27344 3976 27396
rect 4028 27384 4034 27396
rect 4402 27387 4460 27393
rect 4402 27384 4414 27387
rect 4028 27356 4414 27384
rect 4028 27344 4034 27356
rect 4402 27353 4414 27356
rect 4448 27353 4460 27387
rect 4402 27347 4460 27353
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 2222 27316 2228 27328
rect 2183 27288 2228 27316
rect 2222 27276 2228 27288
rect 2280 27276 2286 27328
rect 3878 27276 3884 27328
rect 3936 27316 3942 27328
rect 5537 27319 5595 27325
rect 5537 27316 5549 27319
rect 3936 27288 5549 27316
rect 3936 27276 3942 27288
rect 5537 27285 5549 27288
rect 5583 27285 5595 27319
rect 5537 27279 5595 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1946 27072 1952 27124
rect 2004 27072 2010 27124
rect 3970 27112 3976 27124
rect 3931 27084 3976 27112
rect 3970 27072 3976 27084
rect 4028 27072 4034 27124
rect 1765 26979 1823 26985
rect 1765 26945 1777 26979
rect 1811 26976 1823 26979
rect 1964 26976 1992 27072
rect 2032 27047 2090 27053
rect 2032 27013 2044 27047
rect 2078 27044 2090 27047
rect 2222 27044 2228 27056
rect 2078 27016 2228 27044
rect 2078 27013 2090 27016
rect 2032 27007 2090 27013
rect 2222 27004 2228 27016
rect 2280 27004 2286 27056
rect 2774 26976 2780 26988
rect 1811 26948 2780 26976
rect 1811 26945 1823 26948
rect 1765 26939 1823 26945
rect 2774 26936 2780 26948
rect 2832 26936 2838 26988
rect 4154 26976 4160 26988
rect 4115 26948 4160 26976
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 3142 26772 3148 26784
rect 3103 26744 3148 26772
rect 3142 26732 3148 26744
rect 3200 26732 3206 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 2225 26571 2283 26577
rect 2225 26537 2237 26571
rect 2271 26568 2283 26571
rect 2406 26568 2412 26580
rect 2271 26540 2412 26568
rect 2271 26537 2283 26540
rect 2225 26531 2283 26537
rect 2406 26528 2412 26540
rect 2464 26528 2470 26580
rect 2516 26540 2728 26568
rect 2516 26500 2544 26540
rect 2424 26472 2544 26500
rect 2700 26500 2728 26540
rect 3142 26528 3148 26580
rect 3200 26568 3206 26580
rect 3789 26571 3847 26577
rect 3789 26568 3801 26571
rect 3200 26540 3801 26568
rect 3200 26528 3206 26540
rect 3789 26537 3801 26540
rect 3835 26537 3847 26571
rect 3789 26531 3847 26537
rect 2700 26472 2912 26500
rect 2424 26444 2452 26472
rect 2406 26392 2412 26444
rect 2464 26392 2470 26444
rect 2682 26392 2688 26444
rect 2740 26432 2746 26444
rect 2884 26441 2912 26472
rect 2869 26435 2927 26441
rect 2740 26404 2785 26432
rect 2740 26392 2746 26404
rect 2869 26401 2881 26435
rect 2915 26401 2927 26435
rect 2869 26395 2927 26401
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 2593 26367 2651 26373
rect 2593 26333 2605 26367
rect 2639 26364 2651 26367
rect 3160 26364 3188 26528
rect 4249 26503 4307 26509
rect 4249 26469 4261 26503
rect 4295 26500 4307 26503
rect 4890 26500 4896 26512
rect 4295 26472 4896 26500
rect 4295 26469 4307 26472
rect 4249 26463 4307 26469
rect 4890 26460 4896 26472
rect 4948 26460 4954 26512
rect 3878 26432 3884 26444
rect 3839 26404 3884 26432
rect 3878 26392 3884 26404
rect 3936 26392 3942 26444
rect 15746 26432 15752 26444
rect 3988 26404 15752 26432
rect 3988 26364 4016 26404
rect 15746 26392 15752 26404
rect 15804 26392 15810 26444
rect 2639 26336 3188 26364
rect 3620 26336 4016 26364
rect 4065 26367 4123 26373
rect 2639 26333 2651 26336
rect 2593 26327 2651 26333
rect 1412 26296 1440 26327
rect 3620 26296 3648 26336
rect 4065 26333 4077 26367
rect 4111 26333 4123 26367
rect 4065 26327 4123 26333
rect 3786 26296 3792 26308
rect 1412 26268 3648 26296
rect 3747 26268 3792 26296
rect 3786 26256 3792 26268
rect 3844 26256 3850 26308
rect 3970 26256 3976 26308
rect 4028 26296 4034 26308
rect 4080 26296 4108 26327
rect 4028 26268 4108 26296
rect 4028 26256 4034 26268
rect 1578 26228 1584 26240
rect 1539 26200 1584 26228
rect 1578 26188 1584 26200
rect 1636 26188 1642 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 3418 25848 3424 25900
rect 3476 25888 3482 25900
rect 3881 25891 3939 25897
rect 3881 25888 3893 25891
rect 3476 25860 3893 25888
rect 3476 25848 3482 25860
rect 3881 25857 3893 25860
rect 3927 25857 3939 25891
rect 3881 25851 3939 25857
rect 1397 25687 1455 25693
rect 1397 25653 1409 25687
rect 1443 25684 1455 25687
rect 3602 25684 3608 25696
rect 1443 25656 3608 25684
rect 1443 25653 1455 25656
rect 1397 25647 1455 25653
rect 3602 25644 3608 25656
rect 3660 25644 3666 25696
rect 3697 25687 3755 25693
rect 3697 25653 3709 25687
rect 3743 25684 3755 25687
rect 3878 25684 3884 25696
rect 3743 25656 3884 25684
rect 3743 25653 3755 25656
rect 3697 25647 3755 25653
rect 3878 25644 3884 25656
rect 3936 25644 3942 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 5169 25483 5227 25489
rect 5169 25480 5181 25483
rect 4120 25452 5181 25480
rect 4120 25440 4126 25452
rect 5169 25449 5181 25452
rect 5215 25449 5227 25483
rect 5169 25443 5227 25449
rect 1397 25279 1455 25285
rect 1397 25245 1409 25279
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 1412 25208 1440 25239
rect 1946 25236 1952 25288
rect 2004 25276 2010 25288
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 2004 25248 3801 25276
rect 2004 25236 2010 25248
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 3878 25236 3884 25288
rect 3936 25276 3942 25288
rect 4045 25279 4103 25285
rect 4045 25276 4057 25279
rect 3936 25248 4057 25276
rect 3936 25236 3942 25248
rect 4045 25245 4057 25248
rect 4091 25245 4103 25279
rect 4045 25239 4103 25245
rect 7926 25208 7932 25220
rect 1412 25180 7932 25208
rect 7926 25168 7932 25180
rect 7984 25168 7990 25220
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 3418 24936 3424 24948
rect 3379 24908 3424 24936
rect 3418 24896 3424 24908
rect 3476 24896 3482 24948
rect 3789 24939 3847 24945
rect 3789 24905 3801 24939
rect 3835 24936 3847 24939
rect 4062 24936 4068 24948
rect 3835 24908 4068 24936
rect 3835 24905 3847 24908
rect 3789 24899 3847 24905
rect 4062 24896 4068 24908
rect 4120 24896 4126 24948
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 2222 24760 2228 24812
rect 2280 24800 2286 24812
rect 2409 24803 2467 24809
rect 2409 24800 2421 24803
rect 2280 24772 2421 24800
rect 2280 24760 2286 24772
rect 2409 24769 2421 24772
rect 2455 24769 2467 24803
rect 2409 24763 2467 24769
rect 3602 24760 3608 24812
rect 3660 24800 3666 24812
rect 3881 24803 3939 24809
rect 3881 24800 3893 24803
rect 3660 24772 3893 24800
rect 3660 24760 3666 24772
rect 3881 24769 3893 24772
rect 3927 24769 3939 24803
rect 3881 24763 3939 24769
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24701 4031 24735
rect 3973 24695 4031 24701
rect 1397 24667 1455 24673
rect 1397 24633 1409 24667
rect 1443 24664 1455 24667
rect 2682 24664 2688 24676
rect 1443 24636 2688 24664
rect 1443 24633 1455 24636
rect 1397 24627 1455 24633
rect 2682 24624 2688 24636
rect 2740 24624 2746 24676
rect 2130 24556 2136 24608
rect 2188 24596 2194 24608
rect 2225 24599 2283 24605
rect 2225 24596 2237 24599
rect 2188 24568 2237 24596
rect 2188 24556 2194 24568
rect 2225 24565 2237 24568
rect 2271 24565 2283 24599
rect 2225 24559 2283 24565
rect 2406 24556 2412 24608
rect 2464 24596 2470 24608
rect 3988 24596 4016 24695
rect 2464 24568 4016 24596
rect 2464 24556 2470 24568
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 1946 24188 1952 24200
rect 1903 24160 1952 24188
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 1946 24148 1952 24160
rect 2004 24148 2010 24200
rect 2130 24197 2136 24200
rect 2124 24188 2136 24197
rect 2091 24160 2136 24188
rect 2124 24151 2136 24160
rect 2130 24148 2136 24151
rect 2188 24148 2194 24200
rect 1394 24012 1400 24064
rect 1452 24052 1458 24064
rect 1670 24052 1676 24064
rect 1452 24024 1676 24052
rect 1452 24012 1458 24024
rect 1670 24012 1676 24024
rect 1728 24012 1734 24064
rect 3237 24055 3295 24061
rect 3237 24021 3249 24055
rect 3283 24052 3295 24055
rect 3786 24052 3792 24064
rect 3283 24024 3792 24052
rect 3283 24021 3295 24024
rect 3237 24015 3295 24021
rect 3786 24012 3792 24024
rect 3844 24012 3850 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 2222 23848 2228 23860
rect 2183 23820 2228 23848
rect 2222 23808 2228 23820
rect 2280 23808 2286 23860
rect 2682 23848 2688 23860
rect 2643 23820 2688 23848
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 2593 23783 2651 23789
rect 2593 23749 2605 23783
rect 2639 23780 2651 23783
rect 3786 23780 3792 23792
rect 2639 23752 3792 23780
rect 2639 23749 2651 23752
rect 2593 23743 2651 23749
rect 3786 23740 3792 23752
rect 3844 23740 3850 23792
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23712 1455 23715
rect 1670 23712 1676 23724
rect 1443 23684 1676 23712
rect 1443 23681 1455 23684
rect 1397 23675 1455 23681
rect 1670 23672 1676 23684
rect 1728 23672 1734 23724
rect 3510 23712 3516 23724
rect 3471 23684 3516 23712
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 2406 23604 2412 23656
rect 2464 23644 2470 23656
rect 2777 23647 2835 23653
rect 2777 23644 2789 23647
rect 2464 23616 2789 23644
rect 2464 23604 2470 23616
rect 2777 23613 2789 23616
rect 2823 23644 2835 23647
rect 3697 23647 3755 23653
rect 3697 23644 3709 23647
rect 2823 23616 3709 23644
rect 2823 23613 2835 23616
rect 2777 23607 2835 23613
rect 3697 23613 3709 23616
rect 3743 23613 3755 23647
rect 3697 23607 3755 23613
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 1578 23264 1584 23316
rect 1636 23304 1642 23316
rect 1762 23304 1768 23316
rect 1636 23276 1768 23304
rect 1636 23264 1642 23276
rect 1762 23264 1768 23276
rect 1820 23264 1826 23316
rect 1762 23128 1768 23180
rect 1820 23168 1826 23180
rect 1946 23168 1952 23180
rect 1820 23140 1952 23168
rect 1820 23128 1826 23140
rect 1946 23128 1952 23140
rect 2004 23168 2010 23180
rect 4525 23171 4583 23177
rect 4525 23168 4537 23171
rect 2004 23140 4537 23168
rect 2004 23128 2010 23140
rect 4525 23137 4537 23140
rect 4571 23137 4583 23171
rect 4525 23131 4583 23137
rect 1394 23060 1400 23112
rect 1452 23100 1458 23112
rect 1581 23103 1639 23109
rect 1581 23100 1593 23103
rect 1452 23072 1593 23100
rect 1452 23060 1458 23072
rect 1581 23069 1593 23072
rect 1627 23069 1639 23103
rect 2222 23100 2228 23112
rect 2183 23072 2228 23100
rect 1581 23063 1639 23069
rect 2222 23060 2228 23072
rect 2280 23060 2286 23112
rect 4540 23100 4568 23131
rect 5534 23100 5540 23112
rect 4540 23072 5540 23100
rect 5534 23060 5540 23072
rect 5592 23060 5598 23112
rect 4614 22992 4620 23044
rect 4672 23032 4678 23044
rect 4770 23035 4828 23041
rect 4770 23032 4782 23035
rect 4672 23004 4782 23032
rect 4672 22992 4678 23004
rect 4770 23001 4782 23004
rect 4816 23001 4828 23035
rect 4770 22995 4828 23001
rect 1397 22967 1455 22973
rect 1397 22933 1409 22967
rect 1443 22964 1455 22967
rect 1946 22964 1952 22976
rect 1443 22936 1952 22964
rect 1443 22933 1455 22936
rect 1397 22927 1455 22933
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 2041 22967 2099 22973
rect 2041 22933 2053 22967
rect 2087 22964 2099 22967
rect 3878 22964 3884 22976
rect 2087 22936 3884 22964
rect 2087 22933 2099 22936
rect 2041 22927 2099 22933
rect 3878 22924 3884 22936
rect 3936 22924 3942 22976
rect 3970 22924 3976 22976
rect 4028 22964 4034 22976
rect 5905 22967 5963 22973
rect 5905 22964 5917 22967
rect 4028 22936 5917 22964
rect 4028 22924 4034 22936
rect 5905 22933 5917 22936
rect 5951 22933 5963 22967
rect 5905 22927 5963 22933
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 3878 22760 3884 22772
rect 3839 22732 3884 22760
rect 3878 22720 3884 22732
rect 3936 22720 3942 22772
rect 4614 22760 4620 22772
rect 4575 22732 4620 22760
rect 4614 22720 4620 22732
rect 4672 22720 4678 22772
rect 3789 22695 3847 22701
rect 3789 22661 3801 22695
rect 3835 22692 3847 22695
rect 3970 22692 3976 22704
rect 3835 22664 3976 22692
rect 3835 22661 3847 22664
rect 3789 22655 3847 22661
rect 3970 22652 3976 22664
rect 4028 22652 4034 22704
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22624 1455 22627
rect 2038 22624 2044 22636
rect 1443 22596 2044 22624
rect 1443 22593 1455 22596
rect 1397 22587 1455 22593
rect 2038 22584 2044 22596
rect 2096 22584 2102 22636
rect 2406 22624 2412 22636
rect 2367 22596 2412 22624
rect 2406 22584 2412 22596
rect 2464 22584 2470 22636
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 2682 22516 2688 22568
rect 2740 22556 2746 22568
rect 3973 22559 4031 22565
rect 3973 22556 3985 22559
rect 2740 22528 3985 22556
rect 2740 22516 2746 22528
rect 3973 22525 3985 22528
rect 4019 22525 4031 22559
rect 3973 22519 4031 22525
rect 3421 22491 3479 22497
rect 3421 22457 3433 22491
rect 3467 22488 3479 22491
rect 4816 22488 4844 22587
rect 3467 22460 4844 22488
rect 3467 22457 3479 22460
rect 3421 22451 3479 22457
rect 1210 22380 1216 22432
rect 1268 22420 1274 22432
rect 1581 22423 1639 22429
rect 1581 22420 1593 22423
rect 1268 22392 1593 22420
rect 1268 22380 1274 22392
rect 1581 22389 1593 22392
rect 1627 22389 1639 22423
rect 1581 22383 1639 22389
rect 2130 22380 2136 22432
rect 2188 22420 2194 22432
rect 2225 22423 2283 22429
rect 2225 22420 2237 22423
rect 2188 22392 2237 22420
rect 2188 22380 2194 22392
rect 2225 22389 2237 22392
rect 2271 22389 2283 22423
rect 2225 22383 2283 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 3234 22216 3240 22228
rect 3147 22188 3240 22216
rect 3234 22176 3240 22188
rect 3292 22216 3298 22228
rect 3789 22219 3847 22225
rect 3789 22216 3801 22219
rect 3292 22188 3801 22216
rect 3292 22176 3298 22188
rect 3789 22185 3801 22188
rect 3835 22185 3847 22219
rect 3789 22179 3847 22185
rect 4985 22219 5043 22225
rect 4985 22185 4997 22219
rect 5031 22216 5043 22219
rect 5350 22216 5356 22228
rect 5031 22188 5356 22216
rect 5031 22185 5043 22188
rect 4985 22179 5043 22185
rect 5350 22176 5356 22188
rect 5408 22176 5414 22228
rect 4249 22151 4307 22157
rect 4249 22117 4261 22151
rect 4295 22117 4307 22151
rect 4249 22111 4307 22117
rect 1762 22040 1768 22092
rect 1820 22080 1826 22092
rect 1857 22083 1915 22089
rect 1857 22080 1869 22083
rect 1820 22052 1869 22080
rect 1820 22040 1826 22052
rect 1857 22049 1869 22052
rect 1903 22049 1915 22083
rect 3970 22080 3976 22092
rect 3931 22052 3976 22080
rect 1857 22043 1915 22049
rect 3970 22040 3976 22052
rect 4028 22040 4034 22092
rect 2130 22021 2136 22024
rect 2124 22012 2136 22021
rect 2091 21984 2136 22012
rect 2124 21975 2136 21984
rect 2130 21972 2136 21975
rect 2188 21972 2194 22024
rect 3786 22012 3792 22024
rect 3747 21984 3792 22012
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 4062 22012 4068 22024
rect 4023 21984 4068 22012
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 4264 21944 4292 22111
rect 4798 22080 4804 22092
rect 4759 22052 4804 22080
rect 4798 22040 4804 22052
rect 4856 22040 4862 22092
rect 5534 22040 5540 22092
rect 5592 22080 5598 22092
rect 7009 22083 7067 22089
rect 7009 22080 7021 22083
rect 5592 22052 7021 22080
rect 5592 22040 5598 22052
rect 7009 22049 7021 22052
rect 7055 22049 7067 22083
rect 7009 22043 7067 22049
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 22012 4767 22015
rect 4890 22012 4896 22024
rect 4755 21984 4896 22012
rect 4755 21981 4767 21984
rect 4709 21975 4767 21981
rect 4890 21972 4896 21984
rect 4948 21972 4954 22024
rect 4985 22015 5043 22021
rect 4985 21981 4997 22015
rect 5031 21981 5043 22015
rect 7024 22012 7052 22043
rect 9674 22012 9680 22024
rect 7024 21984 9680 22012
rect 4985 21975 5043 21981
rect 5000 21944 5028 21975
rect 9674 21972 9680 21984
rect 9732 22012 9738 22024
rect 10870 22012 10876 22024
rect 9732 21984 10876 22012
rect 9732 21972 9738 21984
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 7276 21947 7334 21953
rect 4264 21916 5028 21944
rect 5092 21916 6500 21944
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 5092 21876 5120 21916
rect 2280 21848 5120 21876
rect 5169 21879 5227 21885
rect 2280 21836 2286 21848
rect 5169 21845 5181 21879
rect 5215 21876 5227 21879
rect 5258 21876 5264 21888
rect 5215 21848 5264 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 6472 21876 6500 21916
rect 7276 21913 7288 21947
rect 7322 21944 7334 21947
rect 8018 21944 8024 21956
rect 7322 21916 8024 21944
rect 7322 21913 7334 21916
rect 7276 21907 7334 21913
rect 8018 21904 8024 21916
rect 8076 21904 8082 21956
rect 8110 21876 8116 21888
rect 6472 21848 8116 21876
rect 8110 21836 8116 21848
rect 8168 21876 8174 21888
rect 8389 21879 8447 21885
rect 8389 21876 8401 21879
rect 8168 21848 8401 21876
rect 8168 21836 8174 21848
rect 8389 21845 8401 21848
rect 8435 21845 8447 21879
rect 8389 21839 8447 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 2130 21672 2136 21684
rect 1636 21644 2136 21672
rect 1636 21632 1642 21644
rect 2130 21632 2136 21644
rect 2188 21632 2194 21684
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 2406 21672 2412 21684
rect 2271 21644 2412 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 2406 21632 2412 21644
rect 2464 21632 2470 21684
rect 2593 21675 2651 21681
rect 2593 21641 2605 21675
rect 2639 21672 2651 21675
rect 3234 21672 3240 21684
rect 2639 21644 3240 21672
rect 2639 21641 2651 21644
rect 2593 21635 2651 21641
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 8018 21672 8024 21684
rect 7979 21644 8024 21672
rect 8018 21632 8024 21644
rect 8076 21632 8082 21684
rect 17310 21604 17316 21616
rect 1412 21576 17316 21604
rect 1412 21545 1440 21576
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 1670 21496 1676 21548
rect 1728 21496 1734 21548
rect 1946 21496 1952 21548
rect 2004 21536 2010 21548
rect 2685 21539 2743 21545
rect 2685 21536 2697 21539
rect 2004 21508 2697 21536
rect 2004 21496 2010 21508
rect 2685 21505 2697 21508
rect 2731 21505 2743 21539
rect 2685 21499 2743 21505
rect 7466 21496 7472 21548
rect 7524 21536 7530 21548
rect 8205 21539 8263 21545
rect 8205 21536 8217 21539
rect 7524 21508 8217 21536
rect 7524 21496 7530 21508
rect 8205 21505 8217 21508
rect 8251 21505 8263 21539
rect 8205 21499 8263 21505
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21505 8447 21539
rect 8389 21499 8447 21505
rect 1394 21360 1400 21412
rect 1452 21400 1458 21412
rect 1688 21400 1716 21496
rect 2777 21471 2835 21477
rect 2777 21468 2789 21471
rect 2700 21440 2789 21468
rect 2700 21412 2728 21440
rect 2777 21437 2789 21440
rect 2823 21437 2835 21471
rect 8404 21468 8432 21499
rect 8478 21496 8484 21548
rect 8536 21536 8542 21548
rect 9585 21539 9643 21545
rect 8536 21508 8581 21536
rect 8536 21496 8542 21508
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9674 21536 9680 21548
rect 9631 21508 9680 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9674 21496 9680 21508
rect 9732 21496 9738 21548
rect 9852 21539 9910 21545
rect 9852 21505 9864 21539
rect 9898 21536 9910 21539
rect 10410 21536 10416 21548
rect 9898 21508 10416 21536
rect 9898 21505 9910 21508
rect 9852 21499 9910 21505
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 8570 21468 8576 21480
rect 8404 21440 8576 21468
rect 2777 21431 2835 21437
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 1452 21372 1716 21400
rect 1452 21360 1458 21372
rect 2682 21360 2688 21412
rect 2740 21360 2746 21412
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 10962 21332 10968 21344
rect 10923 21304 10968 21332
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1762 21088 1768 21140
rect 1820 21128 1826 21140
rect 1946 21128 1952 21140
rect 1820 21100 1952 21128
rect 1820 21088 1826 21100
rect 1946 21088 1952 21100
rect 2004 21088 2010 21140
rect 8202 21128 8208 21140
rect 8163 21100 8208 21128
rect 8202 21088 8208 21100
rect 8260 21128 8266 21140
rect 9401 21131 9459 21137
rect 9401 21128 9413 21131
rect 8260 21100 9413 21128
rect 8260 21088 8266 21100
rect 9401 21097 9413 21100
rect 9447 21097 9459 21131
rect 10410 21128 10416 21140
rect 10371 21100 10416 21128
rect 9401 21091 9459 21097
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 13078 21128 13084 21140
rect 13039 21100 13084 21128
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 15746 21128 15752 21140
rect 15707 21100 15752 21128
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 1486 21020 1492 21072
rect 1544 21060 1550 21072
rect 1854 21060 1860 21072
rect 1544 21032 1860 21060
rect 1544 21020 1550 21032
rect 1854 21020 1860 21032
rect 1912 21020 1918 21072
rect 7558 21020 7564 21072
rect 7616 21060 7622 21072
rect 10962 21060 10968 21072
rect 7616 21032 10968 21060
rect 7616 21020 7622 21032
rect 2130 20952 2136 21004
rect 2188 20952 2194 21004
rect 4249 20995 4307 21001
rect 4249 20961 4261 20995
rect 4295 20992 4307 20995
rect 5258 20992 5264 21004
rect 4295 20964 5264 20992
rect 4295 20961 4307 20964
rect 4249 20955 4307 20961
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 6181 20995 6239 21001
rect 6181 20992 6193 20995
rect 5592 20964 6193 20992
rect 5592 20952 5598 20964
rect 6181 20961 6193 20964
rect 6227 20961 6239 20995
rect 8110 20992 8116 21004
rect 8071 20964 8116 20992
rect 6181 20955 6239 20961
rect 8110 20952 8116 20964
rect 8168 20952 8174 21004
rect 9508 21001 9536 21032
rect 10962 21020 10968 21032
rect 11020 21020 11026 21072
rect 9493 20995 9551 21001
rect 9493 20961 9505 20995
rect 9539 20961 9551 20995
rect 9493 20955 9551 20961
rect 10612 20964 11836 20992
rect 1578 20924 1584 20936
rect 1539 20896 1584 20924
rect 1578 20884 1584 20896
rect 1636 20884 1642 20936
rect 1854 20884 1860 20936
rect 1912 20924 1918 20936
rect 2148 20924 2176 20952
rect 10612 20936 10640 20964
rect 2406 20924 2412 20936
rect 1912 20896 2176 20924
rect 2367 20896 2412 20924
rect 1912 20884 1918 20896
rect 2406 20884 2412 20896
rect 2464 20884 2470 20936
rect 4525 20927 4583 20933
rect 4525 20893 4537 20927
rect 4571 20924 4583 20927
rect 4706 20924 4712 20936
rect 4571 20896 4712 20924
rect 4571 20893 4583 20896
rect 4525 20887 4583 20893
rect 4706 20884 4712 20896
rect 4764 20884 4770 20936
rect 8021 20927 8079 20933
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 8386 20924 8392 20936
rect 8067 20896 8392 20924
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 8386 20884 8392 20896
rect 8444 20924 8450 20936
rect 9401 20927 9459 20933
rect 9401 20924 9413 20927
rect 8444 20896 9413 20924
rect 8444 20884 8450 20896
rect 9401 20893 9413 20896
rect 9447 20893 9459 20927
rect 10594 20924 10600 20936
rect 10555 20896 10600 20924
rect 9401 20887 9459 20893
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20893 10931 20927
rect 10873 20887 10931 20893
rect 1302 20816 1308 20868
rect 1360 20856 1366 20868
rect 1762 20856 1768 20868
rect 1360 20828 1768 20856
rect 1360 20816 1366 20828
rect 1762 20816 1768 20828
rect 1820 20816 1826 20868
rect 6448 20859 6506 20865
rect 6448 20825 6460 20859
rect 6494 20856 6506 20859
rect 7282 20856 7288 20868
rect 6494 20828 7288 20856
rect 6494 20825 6506 20828
rect 6448 20819 6506 20825
rect 7282 20816 7288 20828
rect 7340 20816 7346 20868
rect 10888 20856 10916 20887
rect 10962 20884 10968 20936
rect 11020 20924 11026 20936
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 11020 20896 11713 20924
rect 11020 20884 11026 20896
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11808 20924 11836 20964
rect 12526 20924 12532 20936
rect 11808 20896 12532 20924
rect 11701 20887 11759 20893
rect 11606 20856 11612 20868
rect 10888 20828 11612 20856
rect 11606 20816 11612 20828
rect 11664 20816 11670 20868
rect 1397 20791 1455 20797
rect 1397 20757 1409 20791
rect 1443 20788 1455 20791
rect 2038 20788 2044 20800
rect 1443 20760 2044 20788
rect 1443 20757 1455 20760
rect 1397 20751 1455 20757
rect 2038 20748 2044 20760
rect 2096 20748 2102 20800
rect 2222 20788 2228 20800
rect 2183 20760 2228 20788
rect 2222 20748 2228 20760
rect 2280 20748 2286 20800
rect 3326 20748 3332 20800
rect 3384 20788 3390 20800
rect 7561 20791 7619 20797
rect 7561 20788 7573 20791
rect 3384 20760 7573 20788
rect 3384 20748 3390 20760
rect 7561 20757 7573 20760
rect 7607 20788 7619 20791
rect 8294 20788 8300 20800
rect 7607 20760 8300 20788
rect 7607 20757 7619 20760
rect 7561 20751 7619 20757
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 8570 20788 8576 20800
rect 8435 20760 8576 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 9769 20791 9827 20797
rect 9769 20757 9781 20791
rect 9815 20788 9827 20791
rect 10781 20791 10839 20797
rect 10781 20788 10793 20791
rect 9815 20760 10793 20788
rect 9815 20757 9827 20760
rect 9769 20751 9827 20757
rect 10781 20757 10793 20760
rect 10827 20757 10839 20791
rect 11716 20788 11744 20887
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20893 14427 20927
rect 14369 20887 14427 20893
rect 11968 20859 12026 20865
rect 11968 20825 11980 20859
rect 12014 20856 12026 20859
rect 12434 20856 12440 20868
rect 12014 20828 12440 20856
rect 12014 20825 12026 20828
rect 11968 20819 12026 20825
rect 12434 20816 12440 20828
rect 12492 20816 12498 20868
rect 14384 20788 14412 20887
rect 14642 20865 14648 20868
rect 14636 20819 14648 20865
rect 14700 20856 14706 20868
rect 14700 20828 14736 20856
rect 14642 20816 14648 20819
rect 14700 20816 14706 20828
rect 11716 20760 14412 20788
rect 10781 20751 10839 20757
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 3326 20584 3332 20596
rect 3239 20556 3332 20584
rect 3326 20544 3332 20556
rect 3384 20584 3390 20596
rect 4062 20584 4068 20596
rect 3384 20556 4068 20584
rect 3384 20544 3390 20556
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 7282 20584 7288 20596
rect 7243 20556 7288 20584
rect 7282 20544 7288 20556
rect 7340 20544 7346 20596
rect 7653 20587 7711 20593
rect 7653 20553 7665 20587
rect 7699 20584 7711 20587
rect 8573 20587 8631 20593
rect 8573 20584 8585 20587
rect 7699 20556 8585 20584
rect 7699 20553 7711 20556
rect 7653 20547 7711 20553
rect 8573 20553 8585 20556
rect 8619 20553 8631 20587
rect 12434 20584 12440 20596
rect 12395 20556 12440 20584
rect 8573 20547 8631 20553
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 14642 20584 14648 20596
rect 14603 20556 14648 20584
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 2222 20525 2228 20528
rect 2216 20516 2228 20525
rect 2183 20488 2228 20516
rect 2216 20479 2228 20488
rect 2222 20476 2228 20479
rect 2280 20476 2286 20528
rect 12636 20488 14872 20516
rect 1946 20448 1952 20460
rect 1907 20420 1952 20448
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 7466 20448 7472 20460
rect 7427 20420 7472 20448
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 7745 20451 7803 20457
rect 7745 20417 7757 20451
rect 7791 20448 7803 20451
rect 7926 20448 7932 20460
rect 7791 20420 7932 20448
rect 7791 20417 7803 20420
rect 7745 20411 7803 20417
rect 7926 20408 7932 20420
rect 7984 20408 7990 20460
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20448 8263 20451
rect 8386 20448 8392 20460
rect 8251 20420 8392 20448
rect 8251 20417 8263 20420
rect 8205 20411 8263 20417
rect 8386 20408 8392 20420
rect 8444 20448 8450 20460
rect 9030 20448 9036 20460
rect 8444 20420 9036 20448
rect 8444 20408 8450 20420
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 12526 20408 12532 20460
rect 12584 20448 12590 20460
rect 12636 20457 12664 20488
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 12584 20420 12633 20448
rect 12584 20408 12590 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 12805 20451 12863 20457
rect 12805 20448 12817 20451
rect 12768 20420 12817 20448
rect 12768 20408 12774 20420
rect 12805 20417 12817 20420
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 13446 20448 13452 20460
rect 12943 20420 13452 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 14844 20457 14872 20488
rect 14829 20451 14887 20457
rect 14829 20417 14841 20451
rect 14875 20417 14887 20451
rect 15010 20448 15016 20460
rect 14971 20420 15016 20448
rect 14829 20411 14887 20417
rect 15010 20408 15016 20420
rect 15068 20408 15074 20460
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15160 20420 15205 20448
rect 15160 20408 15166 20420
rect 8294 20380 8300 20392
rect 8255 20352 8300 20380
rect 8294 20340 8300 20352
rect 8352 20340 8358 20392
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 8202 20244 8208 20256
rect 7432 20216 8208 20244
rect 7432 20204 7438 20216
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 2225 20043 2283 20049
rect 2225 20009 2237 20043
rect 2271 20040 2283 20043
rect 2406 20040 2412 20052
rect 2271 20012 2412 20040
rect 2271 20009 2283 20012
rect 2225 20003 2283 20009
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 2682 20000 2688 20052
rect 2740 20000 2746 20052
rect 7374 20040 7380 20052
rect 7335 20012 7380 20040
rect 7374 20000 7380 20012
rect 7432 20000 7438 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20009 12587 20043
rect 12710 20040 12716 20052
rect 12671 20012 12716 20040
rect 12529 20003 12587 20009
rect 1578 19972 1584 19984
rect 1539 19944 1584 19972
rect 1578 19932 1584 19944
rect 1636 19932 1642 19984
rect 2498 19932 2504 19984
rect 2556 19972 2562 19984
rect 2700 19972 2728 20000
rect 12544 19972 12572 20003
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 14645 20043 14703 20049
rect 14645 20009 14657 20043
rect 14691 20009 14703 20043
rect 15010 20040 15016 20052
rect 14971 20012 15016 20040
rect 14645 20003 14703 20009
rect 12802 19972 12808 19984
rect 2556 19944 2820 19972
rect 12544 19944 12808 19972
rect 2556 19932 2562 19944
rect 2038 19864 2044 19916
rect 2096 19904 2102 19916
rect 2792 19913 2820 19944
rect 12802 19932 12808 19944
rect 12860 19972 12866 19984
rect 14660 19972 14688 20003
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 12860 19944 14688 19972
rect 12860 19932 12866 19944
rect 2685 19907 2743 19913
rect 2685 19904 2697 19907
rect 2096 19876 2697 19904
rect 2096 19864 2102 19876
rect 2685 19873 2697 19876
rect 2731 19873 2743 19907
rect 2685 19867 2743 19873
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19873 2835 19907
rect 8386 19904 8392 19916
rect 2777 19867 2835 19873
rect 7392 19876 8392 19904
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19836 1455 19839
rect 2406 19836 2412 19848
rect 1443 19808 2412 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 2406 19796 2412 19808
rect 2464 19796 2470 19848
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19836 2651 19839
rect 3326 19836 3332 19848
rect 2639 19808 3332 19836
rect 2639 19805 2651 19808
rect 2593 19799 2651 19805
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 6546 19796 6552 19848
rect 6604 19836 6610 19848
rect 7392 19845 7420 19876
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 6604 19808 7389 19836
rect 6604 19796 6610 19808
rect 7377 19805 7389 19808
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 7469 19839 7527 19845
rect 7469 19805 7481 19839
rect 7515 19805 7527 19839
rect 12342 19836 12348 19848
rect 12303 19808 12348 19836
rect 7469 19799 7527 19805
rect 7282 19728 7288 19780
rect 7340 19768 7346 19780
rect 7484 19768 7512 19799
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 13078 19836 13084 19848
rect 12575 19808 13084 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 14642 19836 14648 19848
rect 14603 19808 14648 19836
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 15746 19836 15752 19848
rect 14875 19808 15752 19836
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 7340 19740 7512 19768
rect 7340 19728 7346 19740
rect 7742 19700 7748 19712
rect 7703 19672 7748 19700
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 3694 19456 3700 19508
rect 3752 19496 3758 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 3752 19468 5365 19496
rect 3752 19456 3758 19468
rect 5353 19465 5365 19468
rect 5399 19496 5411 19499
rect 7282 19496 7288 19508
rect 5399 19468 7288 19496
rect 5399 19465 5411 19468
rect 5353 19459 5411 19465
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 7742 19496 7748 19508
rect 7703 19468 7748 19496
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 13998 19496 14004 19508
rect 7852 19468 14004 19496
rect 4240 19431 4298 19437
rect 4240 19397 4252 19431
rect 4286 19428 4298 19431
rect 4286 19400 6776 19428
rect 4286 19397 4298 19400
rect 4240 19391 4298 19397
rect 1578 19360 1584 19372
rect 1539 19332 1584 19360
rect 1578 19320 1584 19332
rect 1636 19320 1642 19372
rect 6546 19360 6552 19372
rect 6507 19332 6552 19360
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 3970 19292 3976 19304
rect 3931 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 5442 19252 5448 19304
rect 5500 19292 5506 19304
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 5500 19264 6653 19292
rect 5500 19252 5506 19264
rect 6641 19261 6653 19264
rect 6687 19261 6699 19295
rect 6748 19292 6776 19400
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7852 19369 7880 19468
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 14829 19499 14887 19505
rect 14829 19465 14841 19499
rect 14875 19496 14887 19499
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 14875 19468 15669 19496
rect 14875 19465 14887 19468
rect 14829 19459 14887 19465
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 12526 19388 12532 19440
rect 12584 19428 12590 19440
rect 12584 19400 15516 19428
rect 12584 19388 12590 19400
rect 7561 19363 7619 19369
rect 7561 19360 7573 19363
rect 7524 19332 7573 19360
rect 7524 19320 7530 19332
rect 7561 19329 7573 19332
rect 7607 19329 7619 19363
rect 7561 19323 7619 19329
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 8202 19320 8208 19372
rect 8260 19360 8266 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 8260 19332 9413 19360
rect 8260 19320 8266 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19360 11851 19363
rect 12342 19360 12348 19372
rect 11839 19332 12348 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 12342 19320 12348 19332
rect 12400 19360 12406 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12400 19332 12817 19360
rect 12400 19320 12406 19332
rect 12805 19329 12817 19332
rect 12851 19360 12863 19363
rect 14274 19360 14280 19372
rect 12851 19332 14280 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 14274 19320 14280 19332
rect 14332 19360 14338 19372
rect 14461 19363 14519 19369
rect 14461 19360 14473 19363
rect 14332 19332 14473 19360
rect 14332 19320 14338 19332
rect 14461 19329 14473 19332
rect 14507 19360 14519 19363
rect 14642 19360 14648 19372
rect 14507 19332 14648 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 15488 19369 15516 19400
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 15804 19332 15849 19360
rect 15804 19320 15810 19332
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 6748 19264 7389 19292
rect 6641 19255 6699 19261
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7377 19255 7435 19261
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19261 9183 19295
rect 9125 19255 9183 19261
rect 6917 19227 6975 19233
rect 6917 19193 6929 19227
rect 6963 19224 6975 19227
rect 7742 19224 7748 19236
rect 6963 19196 7748 19224
rect 6963 19193 6975 19196
rect 6917 19187 6975 19193
rect 7742 19184 7748 19196
rect 7800 19184 7806 19236
rect 9140 19224 9168 19255
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 9732 19264 11529 19292
rect 9732 19252 9738 19264
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 12894 19292 12900 19304
rect 12855 19264 12900 19292
rect 11517 19255 11575 19261
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 14553 19295 14611 19301
rect 14553 19261 14565 19295
rect 14599 19261 14611 19295
rect 14553 19255 14611 19261
rect 9766 19224 9772 19236
rect 9140 19196 9772 19224
rect 9766 19184 9772 19196
rect 9824 19184 9830 19236
rect 14568 19224 14596 19255
rect 16850 19224 16856 19236
rect 12636 19196 16856 19224
rect 1397 19159 1455 19165
rect 1397 19125 1409 19159
rect 1443 19156 1455 19159
rect 2682 19156 2688 19168
rect 1443 19128 2688 19156
rect 1443 19125 1455 19128
rect 1397 19119 1455 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 6733 19159 6791 19165
rect 6733 19125 6745 19159
rect 6779 19156 6791 19159
rect 7374 19156 7380 19168
rect 6779 19128 7380 19156
rect 6779 19125 6791 19128
rect 6733 19119 6791 19125
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 8018 19116 8024 19168
rect 8076 19156 8082 19168
rect 12636 19156 12664 19196
rect 16850 19184 16856 19196
rect 16908 19184 16914 19236
rect 12802 19156 12808 19168
rect 8076 19128 12664 19156
rect 12763 19128 12808 19156
rect 8076 19116 8082 19128
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13170 19156 13176 19168
rect 13131 19128 13176 19156
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 14458 19156 14464 19168
rect 14419 19128 14464 19156
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15562 19156 15568 19168
rect 15335 19128 15568 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 2222 18912 2228 18964
rect 2280 18952 2286 18964
rect 5442 18952 5448 18964
rect 2280 18924 5304 18952
rect 5403 18924 5448 18952
rect 2280 18912 2286 18924
rect 5276 18884 5304 18924
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 9030 18952 9036 18964
rect 8991 18924 9036 18952
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 12345 18955 12403 18961
rect 12345 18952 12357 18955
rect 9140 18924 12357 18952
rect 9140 18884 9168 18924
rect 12345 18921 12357 18924
rect 12391 18952 12403 18955
rect 12894 18952 12900 18964
rect 12391 18924 12900 18952
rect 12391 18921 12403 18924
rect 12345 18915 12403 18921
rect 12894 18912 12900 18924
rect 12952 18912 12958 18964
rect 14277 18955 14335 18961
rect 14277 18921 14289 18955
rect 14323 18952 14335 18955
rect 14458 18952 14464 18964
rect 14323 18924 14464 18952
rect 14323 18921 14335 18924
rect 14277 18915 14335 18921
rect 5276 18856 9168 18884
rect 12802 18844 12808 18896
rect 12860 18884 12866 18896
rect 14292 18884 14320 18915
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 16850 18952 16856 18964
rect 16811 18924 16856 18952
rect 16850 18912 16856 18924
rect 16908 18912 16914 18964
rect 12860 18856 14320 18884
rect 12860 18844 12866 18856
rect 1946 18776 1952 18828
rect 2004 18816 2010 18828
rect 3970 18816 3976 18828
rect 2004 18788 3976 18816
rect 2004 18776 2010 18788
rect 3970 18776 3976 18788
rect 4028 18816 4034 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 4028 18788 4077 18816
rect 4028 18776 4034 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 7466 18776 7472 18828
rect 7524 18816 7530 18828
rect 10962 18816 10968 18828
rect 7524 18788 7604 18816
rect 10923 18788 10968 18816
rect 7524 18776 7530 18788
rect 7576 18760 7604 18788
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 1397 18751 1455 18757
rect 1397 18717 1409 18751
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1412 18680 1440 18711
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 2409 18751 2467 18757
rect 2409 18748 2421 18751
rect 2280 18720 2421 18748
rect 2280 18708 2286 18720
rect 2409 18717 2421 18720
rect 2455 18717 2467 18751
rect 7558 18748 7564 18760
rect 7471 18720 7564 18748
rect 2409 18711 2467 18717
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7742 18748 7748 18760
rect 7703 18720 7748 18748
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 7837 18751 7895 18757
rect 7837 18717 7849 18751
rect 7883 18717 7895 18751
rect 7837 18711 7895 18717
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18748 9275 18751
rect 9674 18748 9680 18760
rect 9263 18720 9680 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 4154 18680 4160 18692
rect 1412 18652 4160 18680
rect 4154 18640 4160 18652
rect 4212 18640 4218 18692
rect 4332 18683 4390 18689
rect 4332 18649 4344 18683
rect 4378 18680 4390 18683
rect 7377 18683 7435 18689
rect 7377 18680 7389 18683
rect 4378 18652 7389 18680
rect 4378 18649 4390 18652
rect 4332 18643 4390 18649
rect 7377 18649 7389 18652
rect 7423 18649 7435 18683
rect 7377 18643 7435 18649
rect 7466 18640 7472 18692
rect 7524 18680 7530 18692
rect 7852 18680 7880 18711
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 12989 18751 13047 18757
rect 12989 18748 13001 18751
rect 12584 18720 13001 18748
rect 12584 18708 12590 18720
rect 12989 18717 13001 18720
rect 13035 18717 13047 18751
rect 13170 18748 13176 18760
rect 13131 18720 13176 18748
rect 12989 18711 13047 18717
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 14274 18748 14280 18760
rect 13320 18720 13365 18748
rect 14235 18720 14280 18748
rect 13320 18708 13326 18720
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 14458 18748 14464 18760
rect 14419 18720 14464 18748
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 7524 18652 7880 18680
rect 11232 18683 11290 18689
rect 7524 18640 7530 18652
rect 11232 18649 11244 18683
rect 11278 18680 11290 18683
rect 12805 18683 12863 18689
rect 12805 18680 12817 18683
rect 11278 18652 12817 18680
rect 11278 18649 11290 18652
rect 11232 18643 11290 18649
rect 12805 18649 12817 18652
rect 12851 18649 12863 18683
rect 12805 18643 12863 18649
rect 13538 18640 13544 18692
rect 13596 18680 13602 18692
rect 15488 18680 15516 18711
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 15729 18751 15787 18757
rect 15729 18748 15741 18751
rect 15620 18720 15741 18748
rect 15620 18708 15626 18720
rect 15729 18717 15741 18720
rect 15775 18717 15787 18751
rect 15729 18711 15787 18717
rect 13596 18652 15516 18680
rect 13596 18640 13602 18652
rect 1578 18612 1584 18624
rect 1539 18584 1584 18612
rect 1578 18572 1584 18584
rect 1636 18572 1642 18624
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 2225 18615 2283 18621
rect 2225 18612 2237 18615
rect 2188 18584 2237 18612
rect 2188 18572 2194 18584
rect 2225 18581 2237 18584
rect 2271 18581 2283 18615
rect 14642 18612 14648 18624
rect 14603 18584 14648 18612
rect 2225 18575 2283 18581
rect 14642 18572 14648 18584
rect 14700 18572 14706 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 2222 18408 2228 18420
rect 2183 18380 2228 18408
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 2682 18408 2688 18420
rect 2643 18380 2688 18408
rect 2682 18368 2688 18380
rect 2740 18368 2746 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 15194 18408 15200 18420
rect 4212 18380 15200 18408
rect 4212 18368 4218 18380
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 1394 18300 1400 18352
rect 1452 18340 1458 18352
rect 14458 18340 14464 18352
rect 1452 18312 14464 18340
rect 1452 18300 1458 18312
rect 14458 18300 14464 18312
rect 14516 18300 14522 18352
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 3234 18272 3240 18284
rect 2639 18244 3240 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 3510 18272 3516 18284
rect 3471 18244 3516 18272
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 7558 18232 7564 18284
rect 7616 18272 7622 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 7616 18244 8033 18272
rect 7616 18232 7622 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 10413 18275 10471 18281
rect 10413 18272 10425 18275
rect 8021 18235 8079 18241
rect 8864 18244 10425 18272
rect 2498 18164 2504 18216
rect 2556 18204 2562 18216
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2556 18176 2789 18204
rect 2556 18164 2562 18176
rect 2777 18173 2789 18176
rect 2823 18173 2835 18207
rect 7742 18204 7748 18216
rect 7703 18176 7748 18204
rect 2777 18167 2835 18173
rect 7742 18164 7748 18176
rect 7800 18204 7806 18216
rect 8864 18204 8892 18244
rect 10413 18241 10425 18244
rect 10459 18241 10471 18275
rect 10594 18272 10600 18284
rect 10555 18244 10600 18272
rect 10413 18235 10471 18241
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 11793 18275 11851 18281
rect 11020 18244 11652 18272
rect 11020 18232 11026 18244
rect 7800 18176 8892 18204
rect 7800 18164 7806 18176
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 9824 18176 11529 18204
rect 9824 18164 9830 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 11624 18204 11652 18244
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 12802 18272 12808 18284
rect 11839 18244 12808 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 13808 18275 13866 18281
rect 13808 18241 13820 18275
rect 13854 18272 13866 18275
rect 14366 18272 14372 18284
rect 13854 18244 14372 18272
rect 13854 18241 13866 18244
rect 13808 18235 13866 18241
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14476 18272 14504 18300
rect 14476 18244 14964 18272
rect 13538 18204 13544 18216
rect 11624 18176 13544 18204
rect 11517 18167 11575 18173
rect 13538 18164 13544 18176
rect 13596 18164 13602 18216
rect 14936 18145 14964 18244
rect 14921 18139 14979 18145
rect 14921 18105 14933 18139
rect 14967 18105 14979 18139
rect 14921 18099 14979 18105
rect 1397 18071 1455 18077
rect 1397 18037 1409 18071
rect 1443 18068 1455 18071
rect 2682 18068 2688 18080
rect 1443 18040 2688 18068
rect 1443 18037 1455 18040
rect 1397 18031 1455 18037
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 3789 18071 3847 18077
rect 3789 18037 3801 18071
rect 3835 18068 3847 18071
rect 4614 18068 4620 18080
rect 3835 18040 4620 18068
rect 3835 18037 3847 18040
rect 3789 18031 3847 18037
rect 4614 18028 4620 18040
rect 4672 18068 4678 18080
rect 5166 18068 5172 18080
rect 4672 18040 5172 18068
rect 4672 18028 4678 18040
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 1820 17836 7297 17864
rect 1820 17824 1826 17836
rect 7285 17833 7297 17836
rect 7331 17864 7343 17867
rect 7374 17864 7380 17876
rect 7331 17836 7380 17864
rect 7331 17833 7343 17836
rect 7285 17827 7343 17833
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 14366 17864 14372 17876
rect 14327 17836 14372 17864
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 7190 17688 7196 17740
rect 7248 17728 7254 17740
rect 7248 17700 8248 17728
rect 7248 17688 7254 17700
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 1946 17660 1952 17672
rect 1903 17632 1952 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2130 17669 2136 17672
rect 2124 17660 2136 17669
rect 2091 17632 2136 17660
rect 2124 17623 2136 17632
rect 2130 17620 2136 17623
rect 2188 17620 2194 17672
rect 5905 17663 5963 17669
rect 5905 17660 5917 17663
rect 2746 17632 5917 17660
rect 1964 17592 1992 17620
rect 2746 17592 2774 17632
rect 5905 17629 5917 17632
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 8220 17669 8248 17700
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7616 17632 7941 17660
rect 7616 17620 7622 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 14424 17632 14565 17660
rect 14424 17620 14430 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 14553 17623 14611 17629
rect 14642 17620 14648 17672
rect 14700 17660 14706 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 14700 17632 14749 17660
rect 14700 17620 14706 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16758 17660 16764 17672
rect 16715 17632 16764 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 1964 17564 2774 17592
rect 6172 17595 6230 17601
rect 6172 17561 6184 17595
rect 6218 17592 6230 17595
rect 7745 17595 7803 17601
rect 7745 17592 7757 17595
rect 6218 17564 7757 17592
rect 6218 17561 6230 17564
rect 6172 17555 6230 17561
rect 7745 17561 7757 17564
rect 7791 17561 7803 17595
rect 7745 17555 7803 17561
rect 14182 17552 14188 17604
rect 14240 17592 14246 17604
rect 14844 17592 14872 17623
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 14240 17564 14872 17592
rect 16936 17595 16994 17601
rect 14240 17552 14246 17564
rect 16936 17561 16948 17595
rect 16982 17592 16994 17595
rect 17218 17592 17224 17604
rect 16982 17564 17224 17592
rect 16982 17561 16994 17564
rect 16936 17555 16994 17561
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 3234 17524 3240 17536
rect 3195 17496 3240 17524
rect 3234 17484 3240 17496
rect 3292 17484 3298 17536
rect 7650 17484 7656 17536
rect 7708 17524 7714 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7708 17496 8125 17524
rect 7708 17484 7714 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 18046 17524 18052 17536
rect 18007 17496 18052 17524
rect 8113 17487 8171 17493
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 7650 17320 7656 17332
rect 7611 17292 7656 17320
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 2406 17212 2412 17264
rect 2464 17252 2470 17264
rect 18046 17252 18052 17264
rect 2464 17224 18052 17252
rect 2464 17212 2470 17224
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 1397 17187 1455 17193
rect 1397 17153 1409 17187
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 1412 17048 1440 17147
rect 2314 17144 2320 17196
rect 2372 17184 2378 17196
rect 5718 17184 5724 17196
rect 2372 17156 5724 17184
rect 2372 17144 2378 17156
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 7282 17184 7288 17196
rect 7243 17156 7288 17184
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 9766 17184 9772 17196
rect 7432 17156 7477 17184
rect 9727 17156 9772 17184
rect 7432 17144 7438 17156
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10226 17184 10232 17196
rect 10187 17156 10232 17184
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 17126 17193 17132 17196
rect 17120 17147 17132 17193
rect 17184 17184 17190 17196
rect 17184 17156 17220 17184
rect 17126 17144 17132 17147
rect 17184 17144 17190 17156
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 1912 17088 10333 17116
rect 1912 17076 1918 17088
rect 10321 17085 10333 17088
rect 10367 17116 10379 17119
rect 11514 17116 11520 17128
rect 10367 17088 11520 17116
rect 10367 17085 10379 17088
rect 10321 17079 10379 17085
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16816 17088 16865 17116
rect 16816 17076 16822 17088
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 11054 17048 11060 17060
rect 1412 17020 11060 17048
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 7469 16983 7527 16989
rect 7469 16980 7481 16983
rect 7432 16952 7481 16980
rect 7432 16940 7438 16952
rect 7469 16949 7481 16952
rect 7515 16980 7527 16983
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 7515 16952 9597 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 9585 16949 9597 16952
rect 9631 16980 9643 16983
rect 10318 16980 10324 16992
rect 9631 16952 10324 16980
rect 9631 16949 9643 16952
rect 9585 16943 9643 16949
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 10597 16983 10655 16989
rect 10597 16949 10609 16983
rect 10643 16980 10655 16983
rect 12342 16980 12348 16992
rect 10643 16952 12348 16980
rect 10643 16949 10655 16952
rect 10597 16943 10655 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 16390 16980 16396 16992
rect 15252 16952 16396 16980
rect 15252 16940 15258 16952
rect 16390 16940 16396 16952
rect 16448 16980 16454 16992
rect 18233 16983 18291 16989
rect 18233 16980 18245 16983
rect 16448 16952 18245 16980
rect 16448 16940 16454 16952
rect 18233 16949 18245 16952
rect 18279 16949 18291 16983
rect 18233 16943 18291 16949
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 7374 16776 7380 16788
rect 7335 16748 7380 16776
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 11514 16776 11520 16788
rect 11475 16748 11520 16776
rect 11514 16736 11520 16748
rect 11572 16736 11578 16788
rect 16669 16779 16727 16785
rect 16669 16745 16681 16779
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 2406 16668 2412 16720
rect 2464 16708 2470 16720
rect 2682 16708 2688 16720
rect 2464 16680 2688 16708
rect 2464 16668 2470 16680
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 16684 16708 16712 16739
rect 17126 16736 17132 16788
rect 17184 16776 17190 16788
rect 17313 16779 17371 16785
rect 17313 16776 17325 16779
rect 17184 16748 17325 16776
rect 17184 16736 17190 16748
rect 17313 16745 17325 16748
rect 17359 16745 17371 16779
rect 17313 16739 17371 16745
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16745 18291 16779
rect 18233 16739 18291 16745
rect 17402 16708 17408 16720
rect 16684 16680 17408 16708
rect 17402 16668 17408 16680
rect 17460 16708 17466 16720
rect 18248 16708 18276 16739
rect 17460 16680 18276 16708
rect 17460 16668 17466 16680
rect 1946 16600 1952 16652
rect 2004 16640 2010 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 2004 16612 4077 16640
rect 2004 16600 2010 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 7377 16643 7435 16649
rect 7377 16609 7389 16643
rect 7423 16609 7435 16643
rect 7377 16603 7435 16609
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 1412 16504 1440 16535
rect 2130 16532 2136 16584
rect 2188 16572 2194 16584
rect 2409 16575 2467 16581
rect 2409 16572 2421 16575
rect 2188 16544 2421 16572
rect 2188 16532 2194 16544
rect 2409 16541 2421 16544
rect 2455 16541 2467 16575
rect 2409 16535 2467 16541
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 7282 16572 7288 16584
rect 6696 16544 7288 16572
rect 6696 16532 6702 16544
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 4062 16504 4068 16516
rect 1412 16476 4068 16504
rect 4062 16464 4068 16476
rect 4120 16464 4126 16516
rect 4332 16507 4390 16513
rect 4332 16473 4344 16507
rect 4378 16504 4390 16507
rect 5350 16504 5356 16516
rect 4378 16476 5356 16504
rect 4378 16473 4390 16476
rect 4332 16467 4390 16473
rect 5350 16464 5356 16476
rect 5408 16464 5414 16516
rect 7392 16504 7420 16603
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16577 16643 16635 16649
rect 16577 16640 16589 16643
rect 16448 16612 16589 16640
rect 16448 16600 16454 16612
rect 16577 16609 16589 16612
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 18046 16600 18052 16652
rect 18104 16640 18110 16652
rect 18325 16643 18383 16649
rect 18325 16640 18337 16643
rect 18104 16612 18337 16640
rect 18104 16600 18110 16612
rect 18325 16609 18337 16612
rect 18371 16609 18383 16643
rect 18325 16603 18383 16609
rect 9674 16572 9680 16584
rect 9635 16544 9680 16572
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16572 10195 16575
rect 10962 16572 10968 16584
rect 10183 16544 10968 16572
rect 10183 16541 10195 16544
rect 10137 16535 10195 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 10226 16504 10232 16516
rect 5460 16476 7420 16504
rect 7576 16476 10232 16504
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 2222 16436 2228 16448
rect 2183 16408 2228 16436
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 5460 16445 5488 16476
rect 5445 16439 5503 16445
rect 5445 16436 5457 16439
rect 2556 16408 5457 16436
rect 2556 16396 2562 16408
rect 5445 16405 5457 16408
rect 5491 16405 5503 16439
rect 5445 16399 5503 16405
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 7576 16436 7604 16476
rect 7340 16408 7604 16436
rect 7653 16439 7711 16445
rect 7340 16396 7346 16408
rect 7653 16405 7665 16439
rect 7699 16436 7711 16439
rect 7834 16436 7840 16448
rect 7699 16408 7840 16436
rect 7699 16405 7711 16408
rect 7653 16399 7711 16405
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 9508 16445 9536 16476
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 10404 16507 10462 16513
rect 10404 16473 10416 16507
rect 10450 16504 10462 16507
rect 12069 16507 12127 16513
rect 12069 16504 12081 16507
rect 10450 16476 12081 16504
rect 10450 16473 10462 16476
rect 10404 16467 10462 16473
rect 12069 16473 12081 16476
rect 12115 16473 12127 16507
rect 12069 16467 12127 16473
rect 9493 16439 9551 16445
rect 9493 16405 9505 16439
rect 9539 16405 9551 16439
rect 9493 16399 9551 16405
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 12268 16436 12296 16535
rect 12342 16532 12348 16584
rect 12400 16572 12406 16584
rect 12437 16575 12495 16581
rect 12437 16572 12449 16575
rect 12400 16544 12449 16572
rect 12400 16532 12406 16544
rect 12437 16541 12449 16544
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16572 12587 16575
rect 15194 16572 15200 16584
rect 12575 16544 15200 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 17586 16572 17592 16584
rect 17543 16544 17592 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 16500 16504 16528 16535
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 17770 16572 17776 16584
rect 17731 16544 17776 16572
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 17126 16504 17132 16516
rect 16500 16476 17132 16504
rect 17126 16464 17132 16476
rect 17184 16504 17190 16516
rect 18248 16504 18276 16535
rect 17184 16476 18276 16504
rect 17184 16464 17190 16476
rect 10928 16408 12296 16436
rect 16853 16439 16911 16445
rect 10928 16396 10934 16408
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 17681 16439 17739 16445
rect 17681 16436 17693 16439
rect 16899 16408 17693 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 17681 16405 17693 16408
rect 17727 16405 17739 16439
rect 18598 16436 18604 16448
rect 18559 16408 18604 16436
rect 17681 16399 17739 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2096 16204 2452 16232
rect 2096 16192 2102 16204
rect 1486 16124 1492 16176
rect 1544 16164 1550 16176
rect 1544 16136 1716 16164
rect 1544 16124 1550 16136
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 1452 16068 1593 16096
rect 1452 16056 1458 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 1688 16096 1716 16136
rect 2222 16124 2228 16176
rect 2280 16173 2286 16176
rect 2280 16167 2344 16173
rect 2280 16133 2298 16167
rect 2332 16133 2344 16167
rect 2424 16164 2452 16204
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 7469 16235 7527 16241
rect 7469 16232 7481 16235
rect 5408 16204 7481 16232
rect 5408 16192 5414 16204
rect 7469 16201 7481 16204
rect 7515 16201 7527 16235
rect 7834 16232 7840 16244
rect 7795 16204 7840 16232
rect 7469 16195 7527 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16201 14887 16235
rect 17218 16232 17224 16244
rect 17179 16204 17224 16232
rect 14829 16195 14887 16201
rect 14550 16164 14556 16176
rect 2424 16136 14556 16164
rect 2280 16127 2344 16133
rect 2280 16124 2286 16127
rect 14550 16124 14556 16136
rect 14608 16164 14614 16176
rect 14844 16164 14872 16195
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 17589 16235 17647 16241
rect 17589 16201 17601 16235
rect 17635 16232 17647 16235
rect 18598 16232 18604 16244
rect 17635 16204 18604 16232
rect 17635 16201 17647 16204
rect 17589 16195 17647 16201
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 14608 16136 14872 16164
rect 14608 16124 14614 16136
rect 6638 16096 6644 16108
rect 1688 16068 6500 16096
rect 6599 16068 6644 16096
rect 1581 16059 1639 16065
rect 1946 15988 1952 16040
rect 2004 16028 2010 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 2004 16000 2053 16028
rect 2004 15988 2010 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 6472 16028 6500 16068
rect 6638 16056 6644 16068
rect 6696 16056 6702 16108
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 7650 16096 7656 16108
rect 6788 16068 6833 16096
rect 7611 16068 7656 16096
rect 6788 16056 6794 16068
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 8202 16096 8208 16108
rect 7975 16068 8208 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10284 16068 10333 16096
rect 10284 16056 10290 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 11773 16099 11831 16105
rect 11773 16096 11785 16099
rect 10836 16068 11785 16096
rect 10836 16056 10842 16068
rect 11773 16065 11785 16068
rect 11819 16065 11831 16099
rect 11773 16059 11831 16065
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 13716 16099 13774 16105
rect 13716 16065 13728 16099
rect 13762 16096 13774 16099
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 13762 16068 15301 16096
rect 13762 16065 13774 16068
rect 13716 16059 13774 16065
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15289 16059 15347 16065
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16065 15531 16099
rect 15654 16096 15660 16108
rect 15615 16068 15660 16096
rect 15473 16059 15531 16065
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 6472 16000 10425 16028
rect 2041 15991 2099 15997
rect 10413 15997 10425 16000
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 5810 15960 5816 15972
rect 3344 15932 5816 15960
rect 1397 15895 1455 15901
rect 1397 15861 1409 15895
rect 1443 15892 1455 15895
rect 3344 15892 3372 15932
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 7374 15960 7380 15972
rect 6840 15932 7380 15960
rect 1443 15864 3372 15892
rect 1443 15861 1455 15864
rect 1397 15855 1455 15861
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 5074 15892 5080 15904
rect 3476 15864 5080 15892
rect 3476 15852 3482 15864
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 6840 15901 6868 15932
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 10428 15960 10456 15991
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 11020 16000 11529 16028
rect 11020 15988 11026 16000
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 12526 15988 12532 16040
rect 12584 16028 12590 16040
rect 13449 16031 13507 16037
rect 13449 16028 13461 16031
rect 12584 16000 13461 16028
rect 12584 15988 12590 16000
rect 13449 15997 13461 16000
rect 13495 16028 13507 16031
rect 13556 16028 13584 16056
rect 13495 16000 13584 16028
rect 13495 15997 13507 16000
rect 13449 15991 13507 15997
rect 14458 15988 14464 16040
rect 14516 16028 14522 16040
rect 14918 16028 14924 16040
rect 14516 16000 14924 16028
rect 14516 15988 14522 16000
rect 14918 15988 14924 16000
rect 14976 16028 14982 16040
rect 15488 16028 15516 16059
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 15838 16096 15844 16108
rect 15795 16068 15844 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 16546 16068 17417 16096
rect 16546 16028 16574 16068
rect 17405 16065 17417 16068
rect 17451 16065 17463 16099
rect 17678 16096 17684 16108
rect 17639 16068 17684 16096
rect 17405 16059 17463 16065
rect 14976 16000 16574 16028
rect 17420 16028 17448 16059
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 17586 16028 17592 16040
rect 17420 16000 17592 16028
rect 14976 15988 14982 16000
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 10428 15932 11284 15960
rect 6825 15895 6883 15901
rect 6825 15861 6837 15895
rect 6871 15861 6883 15895
rect 7006 15892 7012 15904
rect 6967 15864 7012 15892
rect 6825 15855 6883 15861
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 11146 15892 11152 15904
rect 10735 15864 11152 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11256 15892 11284 15932
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 11256 15864 12909 15892
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 6641 15691 6699 15697
rect 4120 15660 6224 15688
rect 4120 15648 4126 15660
rect 1946 15580 1952 15632
rect 2004 15620 2010 15632
rect 6196 15620 6224 15660
rect 6641 15657 6653 15691
rect 6687 15688 6699 15691
rect 6730 15688 6736 15700
rect 6687 15660 6736 15688
rect 6687 15657 6699 15660
rect 6641 15651 6699 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 12526 15688 12532 15700
rect 11020 15660 12532 15688
rect 11020 15648 11026 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 14274 15648 14280 15700
rect 14332 15688 14338 15700
rect 14461 15691 14519 15697
rect 14461 15688 14473 15691
rect 14332 15660 14473 15688
rect 14332 15648 14338 15660
rect 14461 15657 14473 15660
rect 14507 15657 14519 15691
rect 14461 15651 14519 15657
rect 14829 15691 14887 15697
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 15654 15688 15660 15700
rect 14875 15660 15660 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 17402 15688 17408 15700
rect 17363 15660 17408 15688
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 12434 15620 12440 15632
rect 2004 15592 5304 15620
rect 6196 15592 12440 15620
rect 2004 15580 2010 15592
rect 5276 15564 5304 15592
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 2590 15552 2596 15564
rect 2551 15524 2596 15552
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 5258 15552 5264 15564
rect 2740 15524 2785 15552
rect 5171 15524 5264 15552
rect 2740 15512 2746 15524
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 7006 15512 7012 15564
rect 7064 15552 7070 15564
rect 14550 15552 14556 15564
rect 7064 15524 7880 15552
rect 14511 15524 14556 15552
rect 7064 15512 7070 15524
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 3418 15484 3424 15496
rect 2547 15456 3424 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 7650 15484 7656 15496
rect 7563 15456 7656 15484
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 7852 15493 7880 15524
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 16945 15555 17003 15561
rect 16945 15521 16957 15555
rect 16991 15552 17003 15555
rect 17310 15552 17316 15564
rect 16991 15524 17316 15552
rect 16991 15521 17003 15524
rect 16945 15515 17003 15521
rect 17310 15512 17316 15524
rect 17368 15552 17374 15564
rect 17368 15524 17448 15552
rect 17368 15512 17374 15524
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8018 15484 8024 15496
rect 7975 15456 8024 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10928 15456 10977 15484
rect 10928 15444 10934 15456
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 11146 15484 11152 15496
rect 11107 15456 11152 15484
rect 10965 15447 11023 15453
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11974 15484 11980 15496
rect 11287 15456 11980 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 14458 15484 14464 15496
rect 14419 15456 14464 15484
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 17126 15444 17132 15496
rect 17184 15484 17190 15496
rect 17420 15493 17448 15524
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 17184 15456 17233 15484
rect 17184 15444 17190 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 18598 15484 18604 15496
rect 17451 15456 18604 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 18598 15444 18604 15456
rect 18656 15444 18662 15496
rect 5528 15419 5586 15425
rect 5528 15385 5540 15419
rect 5574 15416 5586 15419
rect 7469 15419 7527 15425
rect 7469 15416 7481 15419
rect 5574 15388 7481 15416
rect 5574 15385 5586 15388
rect 5528 15379 5586 15385
rect 7469 15385 7481 15388
rect 7515 15385 7527 15419
rect 7668 15416 7696 15444
rect 8294 15416 8300 15428
rect 7668 15388 8300 15416
rect 7469 15379 7527 15385
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 1394 15348 1400 15360
rect 1355 15320 1400 15348
rect 1394 15308 1400 15320
rect 1452 15308 1458 15360
rect 17589 15351 17647 15357
rect 17589 15317 17601 15351
rect 17635 15348 17647 15351
rect 17862 15348 17868 15360
rect 17635 15320 17868 15348
rect 17635 15317 17647 15320
rect 17589 15311 17647 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 18598 15144 18604 15156
rect 18559 15116 18604 15144
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 8294 15076 8300 15088
rect 8207 15048 8300 15076
rect 8294 15036 8300 15048
rect 8352 15076 8358 15088
rect 10870 15076 10876 15088
rect 8352 15048 10876 15076
rect 8352 15036 8358 15048
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 15008 1455 15011
rect 2038 15008 2044 15020
rect 1443 14980 2044 15008
rect 1443 14977 1455 14980
rect 1397 14971 1455 14977
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 2372 14980 2421 15008
rect 2372 14968 2378 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 7742 15008 7748 15020
rect 7156 14980 7748 15008
rect 7156 14968 7162 14980
rect 7742 14968 7748 14980
rect 7800 15008 7806 15020
rect 10060 15017 10088 15048
rect 10870 15036 10876 15048
rect 10928 15036 10934 15088
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7800 14980 8125 15008
rect 7800 14968 7806 14980
rect 8113 14977 8125 14980
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 10229 15011 10287 15017
rect 10229 14977 10241 15011
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 12158 15008 12164 15020
rect 10367 14980 12164 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10244 14940 10272 14971
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 17494 15017 17500 15020
rect 17488 14971 17500 15017
rect 17552 15008 17558 15020
rect 17552 14980 17588 15008
rect 17494 14968 17500 14971
rect 17552 14968 17558 14980
rect 11238 14940 11244 14952
rect 10244 14912 11244 14940
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 13906 14940 13912 14952
rect 13867 14912 13912 14940
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14940 14243 14943
rect 14274 14940 14280 14952
rect 14231 14912 14280 14940
rect 14231 14909 14243 14912
rect 14185 14903 14243 14909
rect 14274 14900 14280 14912
rect 14332 14900 14338 14952
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 17221 14943 17279 14949
rect 17221 14940 17233 14943
rect 16816 14912 17233 14940
rect 16816 14900 16822 14912
rect 17221 14909 17233 14912
rect 17267 14909 17279 14943
rect 17221 14903 17279 14909
rect 1578 14872 1584 14884
rect 1539 14844 1584 14872
rect 1578 14832 1584 14844
rect 1636 14832 1642 14884
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 10318 14872 10324 14884
rect 5776 14844 10324 14872
rect 5776 14832 5782 14844
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 2222 14804 2228 14816
rect 2183 14776 2228 14804
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 9214 14764 9220 14816
rect 9272 14804 9278 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9272 14776 9873 14804
rect 9272 14764 9278 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 9861 14767 9919 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1397 14603 1455 14609
rect 1397 14569 1409 14603
rect 1443 14569 1455 14603
rect 2314 14600 2320 14612
rect 2275 14572 2320 14600
rect 1397 14563 1455 14569
rect 1412 14532 1440 14563
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 4341 14603 4399 14609
rect 4341 14600 4353 14603
rect 2740 14572 4353 14600
rect 2740 14560 2746 14572
rect 4341 14569 4353 14572
rect 4387 14569 4399 14603
rect 10318 14600 10324 14612
rect 10279 14572 10324 14600
rect 4341 14563 4399 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 10560 14572 10885 14600
rect 10560 14560 10566 14572
rect 10873 14569 10885 14572
rect 10919 14569 10931 14603
rect 11238 14600 11244 14612
rect 11199 14572 11244 14600
rect 10873 14563 10931 14569
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 14332 14572 16865 14600
rect 14332 14560 14338 14572
rect 16853 14569 16865 14572
rect 16899 14600 16911 14603
rect 17310 14600 17316 14612
rect 16899 14572 17316 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 17494 14600 17500 14612
rect 17455 14572 17500 14600
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 4614 14532 4620 14544
rect 1412 14504 4620 14532
rect 4614 14492 4620 14504
rect 4672 14492 4678 14544
rect 1394 14424 1400 14476
rect 1452 14464 1458 14476
rect 2777 14467 2835 14473
rect 2777 14464 2789 14467
rect 1452 14436 2789 14464
rect 1452 14424 1458 14436
rect 2777 14433 2789 14436
rect 2823 14433 2835 14467
rect 2777 14427 2835 14433
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 5810 14464 5816 14476
rect 3007 14436 3041 14464
rect 5771 14436 5816 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 2682 14356 2688 14408
rect 2740 14396 2746 14408
rect 2976 14396 3004 14427
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 10336 14464 10364 14560
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 14918 14532 14924 14544
rect 13587 14504 14924 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 14918 14492 14924 14504
rect 14976 14492 14982 14544
rect 16546 14504 16896 14532
rect 10965 14467 11023 14473
rect 10965 14464 10977 14467
rect 5960 14436 6005 14464
rect 10336 14436 10977 14464
rect 5960 14424 5966 14436
rect 10965 14433 10977 14436
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 16546 14464 16574 14504
rect 11112 14436 16574 14464
rect 11112 14424 11118 14436
rect 5920 14396 5948 14424
rect 16868 14408 16896 14504
rect 2740 14368 5948 14396
rect 2740 14356 2746 14368
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 9214 14405 9220 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8812 14368 8953 14396
rect 8812 14356 8818 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 9208 14396 9220 14405
rect 9175 14368 9220 14396
rect 8941 14359 8999 14365
rect 9208 14359 9220 14368
rect 9214 14356 9220 14359
rect 9272 14356 9278 14408
rect 10870 14396 10876 14408
rect 10831 14368 10876 14396
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 13722 14396 13728 14408
rect 12952 14368 13728 14396
rect 12952 14356 12958 14368
rect 13722 14356 13728 14368
rect 13780 14396 13786 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13780 14368 14105 14396
rect 13780 14356 13786 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 14458 14396 14464 14408
rect 14415 14368 14464 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14458 14356 14464 14368
rect 14516 14396 14522 14408
rect 16669 14399 16727 14405
rect 16669 14396 16681 14399
rect 14516 14368 16681 14396
rect 14516 14356 14522 14368
rect 16669 14365 16681 14368
rect 16715 14365 16727 14399
rect 16850 14396 16856 14408
rect 16811 14368 16856 14396
rect 16669 14359 16727 14365
rect 4246 14328 4252 14340
rect 4207 14300 4252 14328
rect 4246 14288 4252 14300
rect 4304 14288 4310 14340
rect 7742 14328 7748 14340
rect 4356 14300 7748 14328
rect 2685 14263 2743 14269
rect 2685 14229 2697 14263
rect 2731 14260 2743 14263
rect 3326 14260 3332 14272
rect 2731 14232 3332 14260
rect 2731 14229 2743 14232
rect 2685 14223 2743 14229
rect 3326 14220 3332 14232
rect 3384 14260 3390 14272
rect 4356 14260 4384 14300
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13630 14328 13636 14340
rect 13403 14300 13636 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 16684 14328 16712 14359
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17644 14368 17693 14396
rect 17644 14356 17650 14368
rect 17681 14365 17693 14368
rect 17727 14365 17739 14399
rect 17862 14396 17868 14408
rect 17823 14368 17868 14396
rect 17681 14359 17739 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 17957 14399 18015 14405
rect 17957 14365 17969 14399
rect 18003 14396 18015 14399
rect 19334 14396 19340 14408
rect 18003 14368 19340 14396
rect 18003 14365 18015 14368
rect 17957 14359 18015 14365
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 17126 14328 17132 14340
rect 16684 14300 17132 14328
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 5350 14260 5356 14272
rect 3384 14232 4384 14260
rect 5311 14232 5356 14260
rect 3384 14220 3390 14232
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 5718 14260 5724 14272
rect 5679 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 17037 14263 17095 14269
rect 17037 14229 17049 14263
rect 17083 14260 17095 14263
rect 17218 14260 17224 14272
rect 17083 14232 17224 14260
rect 17083 14229 17095 14232
rect 17037 14223 17095 14229
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 2746 14028 14105 14056
rect 2222 13997 2228 14000
rect 2216 13988 2228 13997
rect 2183 13960 2228 13988
rect 2216 13951 2228 13960
rect 2222 13948 2228 13951
rect 2280 13948 2286 14000
rect 1854 13880 1860 13932
rect 1912 13920 1918 13932
rect 2746 13920 2774 14028
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 14108 13988 14136 14019
rect 16850 14016 16856 14068
rect 16908 14056 16914 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 16908 14028 18061 14056
rect 16908 14016 16914 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 14108 13960 14780 13988
rect 1912 13892 2774 13920
rect 1912 13880 1918 13892
rect 3142 13880 3148 13932
rect 3200 13920 3206 13932
rect 3510 13920 3516 13932
rect 3200 13892 3516 13920
rect 3200 13880 3206 13892
rect 3510 13880 3516 13892
rect 3568 13920 3574 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3568 13892 3801 13920
rect 3568 13880 3574 13892
rect 3789 13889 3801 13892
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5408 13892 5733 13920
rect 5408 13880 5414 13892
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 12980 13923 13038 13929
rect 12980 13889 12992 13923
rect 13026 13920 13038 13923
rect 14090 13920 14096 13932
rect 13026 13892 14096 13920
rect 13026 13889 13038 13892
rect 12980 13883 13038 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 14752 13929 14780 13960
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 16758 13920 16764 13932
rect 16715 13892 16764 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 10137 13855 10195 13861
rect 10137 13852 10149 13855
rect 9824 13824 10149 13852
rect 9824 13812 9830 13824
rect 10137 13821 10149 13824
rect 10183 13852 10195 13855
rect 10226 13852 10232 13864
rect 10183 13824 10232 13852
rect 10183 13821 10195 13824
rect 10137 13815 10195 13821
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 10502 13852 10508 13864
rect 10459 13824 10508 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 12526 13852 12532 13864
rect 11756 13824 12532 13852
rect 11756 13812 11762 13824
rect 12526 13812 12532 13824
rect 12584 13852 12590 13864
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12584 13824 12725 13852
rect 12584 13812 12590 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 12713 13815 12771 13821
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 14660 13852 14688 13883
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 16942 13929 16948 13932
rect 16936 13883 16948 13929
rect 17000 13920 17006 13932
rect 17000 13892 17036 13920
rect 16942 13880 16948 13883
rect 17000 13880 17006 13892
rect 13780 13824 14688 13852
rect 13780 13812 13786 13824
rect 3326 13784 3332 13796
rect 3287 13756 3332 13784
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 4246 13744 4252 13796
rect 4304 13744 4310 13796
rect 3973 13719 4031 13725
rect 3973 13685 3985 13719
rect 4019 13716 4031 13719
rect 4264 13716 4292 13744
rect 4798 13716 4804 13728
rect 4019 13688 4804 13716
rect 4019 13685 4031 13688
rect 3973 13679 4031 13685
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 10778 13716 10784 13728
rect 7156 13688 10784 13716
rect 7156 13676 7162 13688
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 14645 13719 14703 13725
rect 14645 13716 14657 13719
rect 13964 13688 14657 13716
rect 13964 13676 13970 13688
rect 14645 13685 14657 13688
rect 14691 13685 14703 13719
rect 15010 13716 15016 13728
rect 14971 13688 15016 13716
rect 14645 13679 14703 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 5626 13512 5632 13524
rect 5460 13484 5632 13512
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5460 13385 5488 13484
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 6822 13512 6828 13524
rect 5776 13484 6828 13512
rect 5776 13472 5782 13484
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 10502 13512 10508 13524
rect 9539 13484 10508 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 14090 13512 14096 13524
rect 14051 13484 14096 13512
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 16853 13515 16911 13521
rect 16853 13481 16865 13515
rect 16899 13512 16911 13515
rect 16942 13512 16948 13524
rect 16899 13484 16948 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 13078 13444 13084 13456
rect 7668 13416 13084 13444
rect 5445 13379 5503 13385
rect 5445 13376 5457 13379
rect 5316 13348 5457 13376
rect 5316 13336 5322 13348
rect 5445 13345 5457 13348
rect 5491 13345 5503 13379
rect 5445 13339 5503 13345
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 1443 13280 5396 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 4249 13243 4307 13249
rect 4249 13209 4261 13243
rect 4295 13240 4307 13243
rect 4798 13240 4804 13252
rect 4295 13212 4804 13240
rect 4295 13209 4307 13212
rect 4249 13203 4307 13209
rect 4798 13200 4804 13212
rect 4856 13240 4862 13252
rect 5368 13240 5396 13280
rect 5534 13268 5540 13320
rect 5592 13308 5598 13320
rect 5701 13311 5759 13317
rect 5701 13308 5713 13311
rect 5592 13280 5713 13308
rect 5592 13268 5598 13280
rect 5701 13277 5713 13280
rect 5747 13277 5759 13311
rect 5701 13271 5759 13277
rect 7558 13240 7564 13252
rect 4856 13212 5304 13240
rect 5368 13212 7564 13240
rect 4856 13200 4862 13212
rect 4338 13172 4344 13184
rect 4299 13144 4344 13172
rect 4338 13132 4344 13144
rect 4396 13132 4402 13184
rect 5276 13172 5304 13212
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 7668 13172 7696 13416
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 10042 13376 10048 13388
rect 9732 13348 10048 13376
rect 9732 13336 9738 13348
rect 10042 13336 10048 13348
rect 10100 13376 10106 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 10100 13348 10149 13376
rect 10100 13336 10106 13348
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 10560 13348 12725 13376
rect 10560 13336 10566 13348
rect 12713 13345 12725 13348
rect 12759 13376 12771 13379
rect 13906 13376 13912 13388
rect 12759 13348 13912 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9490 13308 9496 13320
rect 9451 13280 9496 13308
rect 9309 13271 9367 13277
rect 9324 13240 9352 13271
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 10870 13308 10876 13320
rect 10459 13280 10876 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 10428 13240 10456 13271
rect 10870 13268 10876 13280
rect 10928 13308 10934 13320
rect 12894 13308 12900 13320
rect 10928 13280 12900 13308
rect 10928 13268 10934 13280
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13630 13308 13636 13320
rect 13035 13280 13636 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13780 13280 14289 13308
rect 13780 13268 13786 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 15562 13308 15568 13320
rect 14599 13280 15568 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13277 17095 13311
rect 17218 13308 17224 13320
rect 17179 13280 17224 13308
rect 17037 13271 17095 13277
rect 9324 13212 10456 13240
rect 14461 13243 14519 13249
rect 14461 13209 14473 13243
rect 14507 13240 14519 13243
rect 15010 13240 15016 13252
rect 14507 13212 15016 13240
rect 14507 13209 14519 13212
rect 14461 13203 14519 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 17052 13240 17080 13271
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13308 17371 13311
rect 17494 13308 17500 13320
rect 17359 13280 17500 13308
rect 17359 13277 17371 13280
rect 17313 13271 17371 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 17126 13240 17132 13252
rect 17052 13212 17132 13240
rect 17126 13200 17132 13212
rect 17184 13200 17190 13252
rect 5276 13144 7696 13172
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 10502 13172 10508 13184
rect 9723 13144 10508 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 5810 12968 5816 12980
rect 4571 12940 5816 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 6270 12928 6276 12980
rect 6328 12928 6334 12980
rect 6365 12971 6423 12977
rect 6365 12937 6377 12971
rect 6411 12968 6423 12971
rect 6411 12940 6500 12968
rect 6411 12937 6423 12940
rect 6365 12931 6423 12937
rect 4614 12900 4620 12912
rect 1412 12872 4476 12900
rect 4575 12872 4620 12900
rect 1412 12841 1440 12872
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 2406 12832 2412 12844
rect 2367 12804 2412 12832
rect 1397 12795 1455 12801
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 3050 12832 3056 12844
rect 3011 12804 3056 12832
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 4448 12832 4476 12872
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 6288 12900 6316 12928
rect 4724 12872 6316 12900
rect 4724 12832 4752 12872
rect 4448 12804 4752 12832
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6472 12832 6500 12940
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6788 12940 6837 12968
rect 6788 12928 6794 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 9490 12928 9496 12980
rect 9548 12968 9554 12980
rect 10137 12971 10195 12977
rect 10137 12968 10149 12971
rect 9548 12940 10149 12968
rect 9548 12928 9554 12940
rect 10137 12937 10149 12940
rect 10183 12937 10195 12971
rect 14550 12968 14556 12980
rect 14463 12940 14556 12968
rect 10137 12931 10195 12937
rect 14550 12928 14556 12940
rect 14608 12968 14614 12980
rect 17126 12968 17132 12980
rect 14608 12940 17132 12968
rect 14608 12928 14614 12940
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 18417 12971 18475 12977
rect 18417 12937 18429 12971
rect 18463 12937 18475 12971
rect 18417 12931 18475 12937
rect 7558 12860 7564 12912
rect 7616 12900 7622 12912
rect 18432 12900 18460 12931
rect 7616 12872 18460 12900
rect 7616 12860 7622 12872
rect 5859 12804 6500 12832
rect 6733 12835 6791 12841
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6733 12801 6745 12835
rect 6779 12832 6791 12835
rect 8754 12832 8760 12844
rect 6779 12804 7420 12832
rect 8715 12804 8760 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 4801 12767 4859 12773
rect 4801 12764 4813 12767
rect 4396 12736 4813 12764
rect 4396 12724 4402 12736
rect 4801 12733 4813 12736
rect 4847 12764 4859 12767
rect 5902 12764 5908 12776
rect 4847 12736 5908 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 5902 12724 5908 12736
rect 5960 12764 5966 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 5960 12736 6929 12764
rect 5960 12724 5966 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 7392 12764 7420 12804
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9024 12835 9082 12841
rect 9024 12801 9036 12835
rect 9070 12832 9082 12835
rect 10134 12832 10140 12844
rect 9070 12804 10140 12832
rect 9070 12801 9082 12804
rect 9024 12795 9082 12801
rect 10134 12792 10140 12804
rect 10192 12792 10198 12844
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12952 12804 13093 12832
rect 12952 12792 12958 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 7650 12764 7656 12776
rect 7392 12736 7656 12764
rect 6917 12727 6975 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 13354 12764 13360 12776
rect 13315 12736 13360 12764
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 2869 12699 2927 12705
rect 2869 12665 2881 12699
rect 2915 12696 2927 12699
rect 6730 12696 6736 12708
rect 2915 12668 6736 12696
rect 2915 12665 2927 12668
rect 2869 12659 2927 12665
rect 6730 12656 6736 12668
rect 6788 12656 6794 12708
rect 12342 12696 12348 12708
rect 9692 12668 12348 12696
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4614 12628 4620 12640
rect 4203 12600 4620 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5629 12631 5687 12637
rect 5629 12597 5641 12631
rect 5675 12628 5687 12631
rect 6362 12628 6368 12640
rect 5675 12600 6368 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 9692 12628 9720 12668
rect 12342 12656 12348 12668
rect 12400 12656 12406 12708
rect 10870 12628 10876 12640
rect 6512 12600 9720 12628
rect 10831 12600 10876 12628
rect 6512 12588 6518 12600
rect 10870 12588 10876 12600
rect 10928 12628 10934 12640
rect 13722 12628 13728 12640
rect 10928 12600 13728 12628
rect 10928 12588 10934 12600
rect 13722 12588 13728 12600
rect 13780 12628 13786 12640
rect 14476 12628 14504 12795
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15856 12841 15884 12872
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 15344 12804 15761 12832
rect 15344 12792 15350 12804
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17293 12835 17351 12841
rect 17293 12832 17305 12835
rect 17000 12804 17305 12832
rect 17000 12792 17006 12804
rect 17293 12801 17305 12804
rect 17339 12801 17351 12835
rect 17293 12795 17351 12801
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 16816 12736 17049 12764
rect 16816 12724 16822 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 13780 12600 14504 12628
rect 13780 12588 13786 12600
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15528 12600 15761 12628
rect 15528 12588 15534 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 16117 12631 16175 12637
rect 16117 12597 16129 12631
rect 16163 12628 16175 12631
rect 17310 12628 17316 12640
rect 16163 12600 17316 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2406 12424 2412 12436
rect 2271 12396 2412 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 8754 12424 8760 12436
rect 5684 12396 8760 12424
rect 5684 12384 5690 12396
rect 2682 12248 2688 12300
rect 2740 12288 2746 12300
rect 6288 12297 6316 12396
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 10134 12424 10140 12436
rect 10095 12396 10140 12424
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12400 12396 13093 12424
rect 12400 12384 12406 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 2740 12260 2789 12288
rect 2740 12248 2746 12260
rect 2777 12257 2789 12260
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 13096 12288 13124 12387
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13688 12396 14289 12424
rect 13688 12384 13694 12396
rect 14277 12393 14289 12396
rect 14323 12424 14335 12427
rect 15470 12424 15476 12436
rect 14323 12396 15476 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 16942 12424 16948 12436
rect 16903 12396 16948 12424
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 6273 12251 6331 12257
rect 10612 12260 11836 12288
rect 13096 12260 14197 12288
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 4614 12220 4620 12232
rect 4571 12192 4620 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 6529 12223 6587 12229
rect 6529 12220 6541 12223
rect 6420 12192 6541 12220
rect 6420 12180 6426 12192
rect 6529 12189 6541 12192
rect 6575 12189 6587 12223
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 6529 12183 6587 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10612 12229 10640 12260
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12189 10655 12223
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 10597 12183 10655 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 11808 12220 11836 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 12526 12220 12532 12232
rect 11808 12192 12532 12220
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13354 12220 13360 12232
rect 12768 12192 13360 12220
rect 12768 12180 12774 12192
rect 13354 12180 13360 12192
rect 13412 12220 13418 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13412 12192 14105 12220
rect 13412 12180 13418 12192
rect 14093 12189 14105 12192
rect 14139 12220 14151 12223
rect 15286 12220 15292 12232
rect 14139 12192 15292 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 17126 12220 17132 12232
rect 17087 12192 17132 12220
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17460 12192 17505 12220
rect 17460 12180 17466 12192
rect 2685 12155 2743 12161
rect 2685 12152 2697 12155
rect 1412 12124 2697 12152
rect 1412 12093 1440 12124
rect 2685 12121 2697 12124
rect 2731 12121 2743 12155
rect 2685 12115 2743 12121
rect 11968 12155 12026 12161
rect 11968 12121 11980 12155
rect 12014 12152 12026 12155
rect 13262 12152 13268 12164
rect 12014 12124 13268 12152
rect 12014 12121 12026 12124
rect 11968 12115 12026 12121
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 13722 12152 13728 12164
rect 13556 12124 13728 12152
rect 1397 12087 1455 12093
rect 1397 12053 1409 12087
rect 1443 12053 1455 12087
rect 2590 12084 2596 12096
rect 2551 12056 2596 12084
rect 1397 12047 1455 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 4338 12084 4344 12096
rect 4299 12056 4344 12084
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 7650 12084 7656 12096
rect 7563 12056 7656 12084
rect 7650 12044 7656 12056
rect 7708 12084 7714 12096
rect 8018 12084 8024 12096
rect 7708 12056 8024 12084
rect 7708 12044 7714 12056
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 13556 12084 13584 12124
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 12492 12056 13584 12084
rect 12492 12044 12498 12056
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 13688 12056 14473 12084
rect 13688 12044 13694 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 13262 11880 13268 11892
rect 2096 11852 12434 11880
rect 13223 11852 13268 11880
rect 2096 11840 2102 11852
rect 2124 11815 2182 11821
rect 2124 11781 2136 11815
rect 2170 11812 2182 11815
rect 2222 11812 2228 11824
rect 2170 11784 2228 11812
rect 2170 11781 2182 11784
rect 2124 11775 2182 11781
rect 2222 11772 2228 11784
rect 2280 11772 2286 11824
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 4678 11815 4736 11821
rect 4678 11812 4690 11815
rect 4396 11784 4690 11812
rect 4396 11772 4402 11784
rect 4678 11781 4690 11784
rect 4724 11781 4736 11815
rect 4678 11775 4736 11781
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 10870 11812 10876 11824
rect 10376 11784 10876 11812
rect 10376 11772 10382 11784
rect 10870 11772 10876 11784
rect 10928 11812 10934 11824
rect 11977 11815 12035 11821
rect 11977 11812 11989 11815
rect 10928 11784 11989 11812
rect 10928 11772 10934 11784
rect 11977 11781 11989 11784
rect 12023 11781 12035 11815
rect 11977 11775 12035 11781
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 1946 11744 1952 11756
rect 1903 11716 1952 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11744 4491 11747
rect 5626 11744 5632 11756
rect 4479 11716 5632 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7800 11716 8493 11744
rect 7800 11704 7806 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8680 11676 8708 11707
rect 8260 11648 8708 11676
rect 12406 11676 12434 11852
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13630 11880 13636 11892
rect 13591 11852 13636 11880
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13780 11852 16988 11880
rect 13780 11840 13786 11852
rect 14550 11812 14556 11824
rect 13464 11784 14556 11812
rect 13464 11753 13492 11784
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 16298 11812 16304 11824
rect 15120 11784 16304 11812
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 13449 11707 13507 11713
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 15120 11744 15148 11784
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 16960 11812 16988 11852
rect 16960 11784 17080 11812
rect 15286 11744 15292 11756
rect 13771 11716 15148 11744
rect 15247 11716 15292 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 15286 11704 15292 11716
rect 15344 11744 15350 11756
rect 17052 11753 17080 11784
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 15344 11716 16957 11744
rect 15344 11704 15350 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 18690 11744 18696 11756
rect 17083 11716 18696 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 12406 11648 15393 11676
rect 8260 11636 8266 11648
rect 15381 11645 15393 11648
rect 15427 11676 15439 11679
rect 15930 11676 15936 11688
rect 15427 11648 15936 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 8938 11608 8944 11620
rect 5368 11580 8944 11608
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 3237 11543 3295 11549
rect 3237 11540 3249 11543
rect 2648 11512 3249 11540
rect 2648 11500 2654 11512
rect 3237 11509 3249 11512
rect 3283 11540 3295 11543
rect 5368 11540 5396 11580
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 12161 11611 12219 11617
rect 12161 11577 12173 11611
rect 12207 11608 12219 11611
rect 12250 11608 12256 11620
rect 12207 11580 12256 11608
rect 12207 11577 12219 11580
rect 12161 11571 12219 11577
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 15470 11608 15476 11620
rect 15383 11580 15476 11608
rect 5810 11540 5816 11552
rect 3283 11512 5396 11540
rect 5771 11512 5816 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 8849 11543 8907 11549
rect 8849 11509 8861 11543
rect 8895 11540 8907 11543
rect 9582 11540 9588 11552
rect 8895 11512 9588 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 15396 11549 15424 11580
rect 15470 11568 15476 11580
rect 15528 11608 15534 11620
rect 15528 11580 16988 11608
rect 15528 11568 15534 11580
rect 15381 11543 15439 11549
rect 15381 11509 15393 11543
rect 15427 11509 15439 11543
rect 15654 11540 15660 11552
rect 15615 11512 15660 11540
rect 15381 11503 15439 11509
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16960 11549 16988 11580
rect 16945 11543 17003 11549
rect 16945 11509 16957 11543
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 17313 11543 17371 11549
rect 17313 11509 17325 11543
rect 17359 11540 17371 11543
rect 17862 11540 17868 11552
rect 17359 11512 17868 11540
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 12805 11339 12863 11345
rect 2746 11308 12434 11336
rect 1578 11268 1584 11280
rect 1539 11240 1584 11268
rect 1578 11228 1584 11240
rect 1636 11228 1642 11280
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 2746 11132 2774 11308
rect 6822 11228 6828 11280
rect 6880 11268 6886 11280
rect 6880 11240 9812 11268
rect 6880 11228 6886 11240
rect 8018 11200 8024 11212
rect 7979 11172 8024 11200
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 1443 11104 2774 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8938 11132 8944 11144
rect 8260 11104 8800 11132
rect 8899 11104 8944 11132
rect 8260 11092 8266 11104
rect 8386 11064 8392 11076
rect 8347 11036 8392 11064
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 8772 11064 8800 11104
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 9784 11141 9812 11240
rect 12406 11200 12434 11308
rect 12805 11305 12817 11339
rect 12851 11336 12863 11339
rect 13538 11336 13544 11348
rect 12851 11308 13544 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 15930 11336 15936 11348
rect 15891 11308 15936 11336
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 12526 11228 12532 11280
rect 12584 11268 12590 11280
rect 12584 11240 14596 11268
rect 12584 11228 12590 11240
rect 14568 11200 14596 11240
rect 12406 11172 12848 11200
rect 14568 11172 14688 11200
rect 12820 11144 12848 11172
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9769 11135 9827 11141
rect 9171 11104 9720 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9140 11064 9168 11095
rect 9306 11064 9312 11076
rect 8772 11036 9168 11064
rect 9267 11036 9312 11064
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 9692 11064 9720 11104
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 12618 11132 12624 11144
rect 12579 11104 12624 11132
rect 9953 11095 10011 11101
rect 9968 11064 9996 11095
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 12802 11132 12808 11144
rect 12763 11104 12808 11132
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 14660 11132 14688 11172
rect 16666 11132 16672 11144
rect 14660 11104 16672 11132
rect 14553 11095 14611 11101
rect 9692 11036 9996 11064
rect 10137 11067 10195 11073
rect 10137 11033 10149 11067
rect 10183 11064 10195 11067
rect 10870 11064 10876 11076
rect 10183 11036 10876 11064
rect 10183 11033 10195 11036
rect 10137 11027 10195 11033
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 14568 11064 14596 11095
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 17034 11132 17040 11144
rect 16816 11104 17040 11132
rect 16816 11092 16822 11104
rect 17034 11092 17040 11104
rect 17092 11132 17098 11144
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 17092 11104 17325 11132
rect 17092 11092 17098 11104
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 14820 11067 14878 11073
rect 13688 11036 14780 11064
rect 13688 11024 13694 11036
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12989 10999 13047 11005
rect 12989 10996 13001 10999
rect 12492 10968 13001 10996
rect 12492 10956 12498 10968
rect 12989 10965 13001 10968
rect 13035 10965 13047 10999
rect 14752 10996 14780 11036
rect 14820 11033 14832 11067
rect 14866 11064 14878 11067
rect 15286 11064 15292 11076
rect 14866 11036 15292 11064
rect 14866 11033 14878 11036
rect 14820 11027 14878 11033
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 16776 11064 16804 11092
rect 17586 11073 17592 11076
rect 15396 11036 16804 11064
rect 15396 10996 15424 11036
rect 17580 11027 17592 11073
rect 17644 11064 17650 11076
rect 17644 11036 17680 11064
rect 17586 11024 17592 11027
rect 17644 11024 17650 11036
rect 14752 10968 15424 10996
rect 12989 10959 13047 10965
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 1443 10764 3065 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 12897 10755 12955 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15654 10792 15660 10804
rect 15615 10764 15660 10792
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 17497 10795 17555 10801
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 17586 10792 17592 10804
rect 17543 10764 17592 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 17862 10792 17868 10804
rect 17823 10764 17868 10792
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 11698 10724 11704 10736
rect 11532 10696 11704 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3878 10656 3884 10668
rect 3007 10628 3884 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8202 10656 8208 10668
rect 7984 10628 8208 10656
rect 7984 10616 7990 10628
rect 8202 10616 8208 10628
rect 8260 10656 8266 10668
rect 11532 10665 11560 10696
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 17126 10724 17132 10736
rect 15488 10696 17132 10724
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8260 10628 8677 10656
rect 8260 10616 8266 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11784 10659 11842 10665
rect 11784 10625 11796 10659
rect 11830 10656 11842 10659
rect 12066 10656 12072 10668
rect 11830 10628 12072 10656
rect 11830 10625 11842 10628
rect 11784 10619 11842 10625
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 15488 10665 15516 10696
rect 17126 10684 17132 10696
rect 17184 10724 17190 10736
rect 17184 10696 17724 10724
rect 17184 10684 17190 10696
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 16574 10656 16580 10668
rect 15795 10628 16580 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 17696 10665 17724 10696
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17957 10659 18015 10665
rect 17957 10625 17969 10659
rect 18003 10656 18015 10659
rect 18414 10656 18420 10668
rect 18003 10628 18420 10656
rect 18003 10625 18015 10628
rect 17957 10619 18015 10625
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 3142 10588 3148 10600
rect 3103 10560 3148 10588
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 5868 10560 8493 10588
rect 5868 10548 5874 10560
rect 8481 10557 8493 10560
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 2593 10455 2651 10461
rect 2593 10421 2605 10455
rect 2639 10452 2651 10455
rect 2866 10452 2872 10464
rect 2639 10424 2872 10452
rect 2639 10421 2651 10424
rect 2593 10415 2651 10421
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10452 8907 10455
rect 15930 10452 15936 10464
rect 8895 10424 15936 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10217 5319 10251
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5261 10211 5319 10217
rect 5276 10180 5304 10211
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 12066 10248 12072 10260
rect 12027 10220 12072 10248
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 5626 10180 5632 10192
rect 5276 10152 5632 10180
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 3292 10016 4997 10044
rect 3292 10004 3298 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 4985 10007 5043 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5810 10044 5816 10056
rect 5307 10016 5816 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10044 6147 10047
rect 6730 10044 6736 10056
rect 6135 10016 6736 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10044 8171 10047
rect 8202 10044 8208 10056
rect 8159 10016 8208 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 12250 10044 12256 10056
rect 12211 10016 12256 10044
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 14366 10044 14372 10056
rect 12575 10016 14372 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 6362 9985 6368 9988
rect 6356 9939 6368 9985
rect 6420 9976 6426 9988
rect 6420 9948 6456 9976
rect 6362 9936 6368 9939
rect 6420 9936 6426 9948
rect 2685 9911 2743 9917
rect 2685 9877 2697 9911
rect 2731 9908 2743 9911
rect 2866 9908 2872 9920
rect 2731 9880 2872 9908
rect 2731 9877 2743 9880
rect 2685 9871 2743 9877
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 8846 9908 8852 9920
rect 7515 9880 8852 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12492 9880 12537 9908
rect 12492 9868 12498 9880
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 2866 9704 2872 9716
rect 2792 9676 2872 9704
rect 2792 9645 2820 9676
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 6362 9704 6368 9716
rect 6323 9676 6368 9704
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 2768 9639 2826 9645
rect 2768 9605 2780 9639
rect 2814 9605 2826 9639
rect 2768 9599 2826 9605
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 15841 9639 15899 9645
rect 15841 9636 15853 9639
rect 3016 9608 15853 9636
rect 3016 9596 3022 9608
rect 15841 9605 15853 9608
rect 15887 9605 15899 9639
rect 15841 9599 15899 9605
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9568 1455 9571
rect 1443 9540 6132 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2406 9500 2412 9512
rect 2004 9472 2412 9500
rect 2004 9460 2010 9472
rect 2406 9460 2412 9472
rect 2464 9500 2470 9512
rect 2501 9503 2559 9509
rect 2501 9500 2513 9503
rect 2464 9472 2513 9500
rect 2464 9460 2470 9472
rect 2501 9469 2513 9472
rect 2547 9469 2559 9503
rect 2501 9463 2559 9469
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3878 9364 3884 9376
rect 3839 9336 3884 9364
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 6104 9364 6132 9540
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6236 9540 6561 9568
rect 6236 9528 6242 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 10042 9568 10048 9580
rect 6549 9531 6607 9537
rect 8956 9540 10048 9568
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8956 9509 8984 9540
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 15746 9568 15752 9580
rect 15707 9540 15752 9568
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 16022 9528 16028 9580
rect 16080 9568 16086 9580
rect 16925 9571 16983 9577
rect 16925 9568 16937 9571
rect 16080 9540 16937 9568
rect 16080 9528 16086 9540
rect 16925 9537 16937 9540
rect 16971 9537 16983 9571
rect 16925 9531 16983 9537
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 7892 9472 8493 9500
rect 7892 9460 7898 9472
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9500 10379 9503
rect 10778 9500 10784 9512
rect 10367 9472 10784 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 13078 9460 13084 9512
rect 13136 9500 13142 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 13136 9472 15945 9500
rect 13136 9460 13142 9472
rect 15933 9469 15945 9472
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 8846 9432 8852 9444
rect 8807 9404 8852 9432
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 10594 9392 10600 9444
rect 10652 9432 10658 9444
rect 11698 9432 11704 9444
rect 10652 9404 11704 9432
rect 10652 9392 10658 9404
rect 11698 9392 11704 9404
rect 11756 9392 11762 9444
rect 10962 9364 10968 9376
rect 6104 9336 10968 9364
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 15381 9367 15439 9373
rect 15381 9333 15393 9367
rect 15427 9364 15439 9367
rect 16114 9364 16120 9376
rect 15427 9336 16120 9364
rect 15427 9333 15439 9336
rect 15381 9327 15439 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16684 9364 16712 9463
rect 17034 9364 17040 9376
rect 16684 9336 17040 9364
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 18046 9364 18052 9376
rect 18007 9336 18052 9364
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 5994 9160 6000 9172
rect 5955 9132 6000 9160
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6178 9160 6184 9172
rect 6139 9132 6184 9160
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11020 9132 11989 9160
rect 11020 9120 11026 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 11977 9123 12035 9129
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16022 9160 16028 9172
rect 15979 9132 16028 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 1397 9095 1455 9101
rect 1397 9061 1409 9095
rect 1443 9092 1455 9095
rect 2958 9092 2964 9104
rect 1443 9064 2964 9092
rect 1443 9061 1455 9064
rect 1397 9055 1455 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 5626 9092 5632 9104
rect 5587 9064 5632 9092
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 19245 9095 19303 9101
rect 19245 9092 19257 9095
rect 11624 9064 19257 9092
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2774 8956 2780 8968
rect 2271 8928 2780 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 5644 8956 5672 9052
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 7742 9024 7748 9036
rect 7607 8996 7748 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 7742 8984 7748 8996
rect 7800 9024 7806 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 7800 8996 9137 9024
rect 7800 8984 7806 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10226 9024 10232 9036
rect 10091 8996 10232 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10594 9024 10600 9036
rect 10555 8996 10600 9024
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 7834 8956 7840 8968
rect 5644 8928 7840 8956
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8720 8928 9229 8956
rect 8720 8916 8726 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 11624 8956 11652 9064
rect 19245 9061 19257 9064
rect 19291 9061 19303 9095
rect 19245 9055 19303 9061
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 17681 9027 17739 9033
rect 17681 9024 17693 9027
rect 12216 8996 17693 9024
rect 12216 8984 12222 8996
rect 17681 8993 17693 8996
rect 17727 8993 17739 9027
rect 17681 8987 17739 8993
rect 13354 8956 13360 8968
rect 9217 8919 9275 8925
rect 10704 8928 11652 8956
rect 13315 8928 13360 8956
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 10704 8888 10732 8928
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 16114 8956 16120 8968
rect 16075 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 17862 8956 17868 8968
rect 17823 8928 17868 8956
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 19150 8956 19156 8968
rect 18187 8928 19156 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 19150 8916 19156 8928
rect 19208 8916 19214 8968
rect 19426 8956 19432 8968
rect 19387 8928 19432 8956
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20530 8956 20536 8968
rect 19751 8928 20536 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 8168 8860 10732 8888
rect 10864 8891 10922 8897
rect 8168 8848 8174 8860
rect 10864 8857 10876 8891
rect 10910 8888 10922 8891
rect 11514 8888 11520 8900
rect 10910 8860 11520 8888
rect 10910 8857 10922 8860
rect 10864 8851 10922 8857
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 20346 8888 20352 8900
rect 12406 8860 20352 8888
rect 2038 8820 2044 8832
rect 1999 8792 2044 8820
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5960 8792 6009 8820
rect 5960 8780 5966 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 12406 8820 12434 8860
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 13170 8820 13176 8832
rect 8076 8792 12434 8820
rect 13131 8792 13176 8820
rect 8076 8780 8082 8792
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19300 8792 19625 8820
rect 19300 8780 19306 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19613 8783 19671 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8585 1823 8619
rect 1765 8579 1823 8585
rect 1780 8548 1808 8579
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 11054 8616 11060 8628
rect 2096 8588 11060 8616
rect 2096 8576 2102 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11514 8616 11520 8628
rect 11475 8588 11520 8616
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 11756 8588 12434 8616
rect 11756 8576 11762 8588
rect 2654 8551 2712 8557
rect 2654 8548 2666 8551
rect 1780 8520 2666 8548
rect 2654 8517 2666 8520
rect 2700 8517 2712 8551
rect 2654 8511 2712 8517
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 5868 8520 6469 8548
rect 5868 8508 5874 8520
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 6914 8548 6920 8560
rect 6503 8520 6920 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7742 8548 7748 8560
rect 7703 8520 7748 8548
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 8113 8551 8171 8557
rect 8113 8517 8125 8551
rect 8159 8548 8171 8551
rect 8202 8548 8208 8560
rect 8159 8520 8208 8548
rect 8159 8517 8171 8520
rect 8113 8511 8171 8517
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 12250 8548 12256 8560
rect 11716 8520 12256 8548
rect 11716 8492 11744 8520
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 12406 8548 12434 8588
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15804 8588 16037 8616
rect 15804 8576 15810 8588
rect 16025 8585 16037 8588
rect 16071 8616 16083 8619
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16071 8588 17049 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 20346 8616 20352 8628
rect 20307 8588 20352 8616
rect 17037 8579 17095 8585
rect 12406 8520 13124 8548
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2406 8480 2412 8492
rect 2367 8452 2412 8480
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5960 8452 6377 8480
rect 5960 8440 5966 8452
rect 6365 8449 6377 8452
rect 6411 8480 6423 8483
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 6411 8452 7941 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 7929 8449 7941 8452
rect 7975 8480 7987 8483
rect 8662 8480 8668 8492
rect 7975 8452 8668 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10226 8480 10232 8492
rect 10183 8452 10232 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 11698 8480 11704 8492
rect 11611 8452 11704 8480
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12526 8480 12532 8492
rect 12023 8452 12532 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 13096 8489 13124 8520
rect 13170 8508 13176 8560
rect 13228 8548 13234 8560
rect 13326 8551 13384 8557
rect 13326 8548 13338 8551
rect 13228 8520 13338 8548
rect 13228 8508 13234 8520
rect 13326 8517 13338 8520
rect 13372 8517 13384 8551
rect 16666 8548 16672 8560
rect 16627 8520 16672 8548
rect 13326 8511 13384 8517
rect 16666 8508 16672 8520
rect 16724 8508 16730 8560
rect 17052 8548 17080 8579
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 18046 8548 18052 8560
rect 17052 8520 18052 8548
rect 18046 8508 18052 8520
rect 18104 8548 18110 8560
rect 18104 8520 18184 8548
rect 18104 8508 18110 8520
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13630 8480 13636 8492
rect 13127 8452 13636 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 15930 8480 15936 8492
rect 15887 8452 15936 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 16114 8480 16120 8492
rect 16075 8452 16120 8480
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17678 8480 17684 8492
rect 17175 8452 17684 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 10502 8412 10508 8424
rect 10459 8384 10508 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 15948 8412 15976 8440
rect 16868 8412 16896 8443
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 18156 8489 18184 8520
rect 19242 8508 19248 8560
rect 19300 8548 19306 8560
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 19300 8520 19809 8548
rect 19300 8508 19306 8520
rect 19797 8517 19809 8520
rect 19843 8548 19855 8551
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 19843 8520 20729 8548
rect 19843 8517 19855 8520
rect 19797 8511 19855 8517
rect 20717 8517 20729 8520
rect 20763 8517 20775 8551
rect 20717 8511 20775 8517
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8480 18475 8483
rect 19260 8480 19288 8508
rect 18463 8452 19288 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 19484 8452 19625 8480
rect 19484 8440 19490 8452
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20438 8480 20444 8492
rect 19935 8452 20444 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 15948 8384 16896 8412
rect 19628 8412 19656 8443
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 20548 8412 20576 8443
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 20864 8452 20909 8480
rect 20864 8440 20870 8452
rect 19628 8384 20576 8412
rect 15194 8304 15200 8356
rect 15252 8344 15258 8356
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 15252 8316 19441 8344
rect 15252 8304 15258 8316
rect 19429 8313 19441 8316
rect 19475 8313 19487 8347
rect 19429 8307 19487 8313
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 14458 8276 14464 8288
rect 14419 8248 14464 8276
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 19628 8276 19656 8384
rect 17920 8248 19656 8276
rect 17920 8236 17926 8248
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2501 8075 2559 8081
rect 2501 8072 2513 8075
rect 2004 8044 2513 8072
rect 2004 8032 2010 8044
rect 2501 8041 2513 8044
rect 2547 8041 2559 8075
rect 2501 8035 2559 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7524 8044 7696 8072
rect 7524 8032 7530 8044
rect 7668 8004 7696 8044
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7800 8044 8125 8072
rect 7800 8032 7806 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 10560 8044 10793 8072
rect 10560 8032 10566 8044
rect 10781 8041 10793 8044
rect 10827 8041 10839 8075
rect 10781 8035 10839 8041
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 11882 8072 11888 8084
rect 11195 8044 11888 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8072 12863 8075
rect 13354 8072 13360 8084
rect 12851 8044 13360 8072
rect 12851 8041 12863 8044
rect 12805 8035 12863 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 11238 8004 11244 8016
rect 7668 7976 11244 8004
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 19245 8007 19303 8013
rect 19245 8004 19257 8007
rect 12032 7976 19257 8004
rect 12032 7964 12038 7976
rect 19245 7973 19257 7976
rect 19291 7973 19303 8007
rect 19245 7967 19303 7973
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 3142 7936 3148 7948
rect 3103 7908 3148 7936
rect 3142 7896 3148 7908
rect 3200 7936 3206 7948
rect 3602 7936 3608 7948
rect 3200 7908 3608 7936
rect 3200 7896 3206 7908
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 11112 7908 13277 7936
rect 11112 7896 11118 7908
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7905 13415 7939
rect 17862 7936 17868 7948
rect 17823 7908 17868 7936
rect 13357 7899 13415 7905
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 6730 7868 6736 7880
rect 1443 7840 2774 7868
rect 6691 7840 6736 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 2746 7800 2774 7840
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10962 7868 10968 7880
rect 10923 7840 10968 7868
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 13372 7868 13400 7899
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 14274 7868 14280 7880
rect 13136 7840 13400 7868
rect 14235 7840 14280 7868
rect 13136 7828 13142 7840
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 14826 7868 14832 7880
rect 14599 7840 14832 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 17184 7840 17601 7868
rect 17184 7828 17190 7840
rect 17589 7837 17601 7840
rect 17635 7837 17647 7871
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 17589 7831 17647 7837
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 20622 7868 20628 7880
rect 19751 7840 20628 7868
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 7000 7803 7058 7809
rect 2746 7772 6960 7800
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 3786 7732 3792 7744
rect 2915 7704 3792 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 6932 7732 6960 7772
rect 7000 7769 7012 7803
rect 7046 7800 7058 7803
rect 7098 7800 7104 7812
rect 7046 7772 7104 7800
rect 7046 7769 7058 7772
rect 7000 7763 7058 7769
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 8478 7760 8484 7812
rect 8536 7800 8542 7812
rect 14093 7803 14151 7809
rect 14093 7800 14105 7803
rect 8536 7772 14105 7800
rect 8536 7760 8542 7772
rect 14093 7769 14105 7772
rect 14139 7769 14151 7803
rect 14093 7763 14151 7769
rect 19242 7760 19248 7812
rect 19300 7800 19306 7812
rect 19613 7803 19671 7809
rect 19613 7800 19625 7803
rect 19300 7772 19625 7800
rect 19300 7760 19306 7772
rect 19613 7769 19625 7772
rect 19659 7769 19671 7803
rect 19613 7763 19671 7769
rect 10594 7732 10600 7744
rect 6932 7704 10600 7732
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 13173 7735 13231 7741
rect 13173 7701 13185 7735
rect 13219 7732 13231 7735
rect 13814 7732 13820 7744
rect 13219 7704 13820 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 13814 7692 13820 7704
rect 13872 7732 13878 7744
rect 14458 7732 14464 7744
rect 13872 7704 14464 7732
rect 13872 7692 13878 7704
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 3050 7528 3056 7540
rect 2179 7500 3056 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5902 7528 5908 7540
rect 5215 7500 5908 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 7098 7528 7104 7540
rect 7059 7500 7104 7528
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 13173 7531 13231 7537
rect 13173 7528 13185 7531
rect 7984 7500 13185 7528
rect 7984 7488 7990 7500
rect 13173 7497 13185 7500
rect 13219 7497 13231 7531
rect 13173 7491 13231 7497
rect 13541 7531 13599 7537
rect 13541 7497 13553 7531
rect 13587 7528 13599 7531
rect 13814 7528 13820 7540
rect 13587 7500 13820 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13814 7488 13820 7500
rect 13872 7488 13878 7540
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 14056 7500 14105 7528
rect 14056 7488 14062 7500
rect 14093 7497 14105 7500
rect 14139 7497 14151 7531
rect 14093 7491 14151 7497
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 15381 7531 15439 7537
rect 15381 7528 15393 7531
rect 14516 7500 15393 7528
rect 14516 7488 14522 7500
rect 15381 7497 15393 7500
rect 15427 7497 15439 7531
rect 15381 7491 15439 7497
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7528 18843 7531
rect 19242 7528 19248 7540
rect 18831 7500 19248 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 2685 7463 2743 7469
rect 2685 7429 2697 7463
rect 2731 7460 2743 7463
rect 4706 7460 4712 7472
rect 2731 7432 4712 7460
rect 2731 7429 2743 7432
rect 2685 7423 2743 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 7558 7420 7564 7472
rect 7616 7460 7622 7472
rect 15013 7463 15071 7469
rect 15013 7460 15025 7463
rect 7616 7432 15025 7460
rect 7616 7420 7622 7432
rect 15013 7429 15025 7432
rect 15059 7429 15071 7463
rect 15013 7423 15071 7429
rect 15212 7432 17448 7460
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 2648 7364 2693 7392
rect 2648 7352 2654 7364
rect 3326 7352 3332 7404
rect 3384 7392 3390 7404
rect 4045 7395 4103 7401
rect 4045 7392 4057 7395
rect 3384 7364 4057 7392
rect 3384 7352 3390 7364
rect 4045 7361 4057 7364
rect 4091 7361 4103 7395
rect 4045 7355 4103 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6052 7364 6377 7392
rect 6052 7352 6058 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6549 7355 6607 7361
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 3789 7327 3847 7333
rect 3789 7324 3801 7327
rect 2832 7296 3801 7324
rect 2832 7284 2838 7296
rect 3789 7293 3801 7296
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 3804 7188 3832 7287
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 6564 7324 6592 7355
rect 6914 7352 6920 7364
rect 6972 7392 6978 7404
rect 7466 7392 7472 7404
rect 6972 7364 7472 7392
rect 6972 7352 6978 7364
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 7892 7364 8585 7392
rect 7892 7352 7898 7364
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 8846 7392 8852 7404
rect 8720 7364 8765 7392
rect 8807 7364 8852 7392
rect 8720 7352 8726 7364
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 4856 7296 6592 7324
rect 6641 7327 6699 7333
rect 4856 7284 4862 7296
rect 6641 7293 6653 7327
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 9766 7324 9772 7336
rect 6779 7296 9772 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 6656 7256 6684 7287
rect 9766 7284 9772 7296
rect 9824 7324 9830 7336
rect 10520 7324 10548 7355
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 13357 7395 13415 7401
rect 10652 7364 10697 7392
rect 10652 7352 10658 7364
rect 13357 7361 13369 7395
rect 13403 7361 13415 7395
rect 13630 7392 13636 7404
rect 13591 7364 13636 7392
rect 13357 7355 13415 7361
rect 10778 7324 10784 7336
rect 9824 7296 10784 7324
rect 9824 7284 9830 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 13372 7324 13400 7355
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 14274 7392 14280 7404
rect 14187 7364 14280 7392
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 15212 7401 15240 7432
rect 15197 7395 15255 7401
rect 14608 7364 14653 7392
rect 14608 7352 14614 7364
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 14292 7324 14320 7352
rect 15212 7324 15240 7355
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 17420 7401 17448 7432
rect 17405 7395 17463 7401
rect 15528 7364 15573 7392
rect 15528 7352 15534 7364
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17451 7364 18613 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 18966 7392 18972 7404
rect 18923 7364 18972 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 17126 7324 17132 7336
rect 13372 7296 15240 7324
rect 17087 7296 17132 7324
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 5500 7228 6684 7256
rect 9217 7259 9275 7265
rect 5500 7216 5506 7228
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 11054 7256 11060 7268
rect 9263 7228 11060 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 11296 7228 18429 7256
rect 11296 7216 11302 7228
rect 18417 7225 18429 7228
rect 18463 7225 18475 7259
rect 18417 7219 18475 7225
rect 6730 7188 6736 7200
rect 3804 7160 6736 7188
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 10502 7188 10508 7200
rect 10463 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10870 7188 10876 7200
rect 10831 7160 10876 7188
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 2869 6987 2927 6993
rect 2869 6984 2881 6987
rect 2648 6956 2881 6984
rect 2648 6944 2654 6956
rect 2869 6953 2881 6956
rect 2915 6984 2927 6987
rect 4614 6984 4620 6996
rect 2915 6956 4620 6984
rect 2915 6953 2927 6956
rect 2869 6947 2927 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 6052 6956 6101 6984
rect 6052 6944 6058 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 7377 6987 7435 6993
rect 7377 6953 7389 6987
rect 7423 6984 7435 6987
rect 7834 6984 7840 6996
rect 7423 6956 7840 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 4522 6876 4528 6928
rect 4580 6916 4586 6928
rect 4706 6916 4712 6928
rect 4580 6888 4712 6916
rect 4580 6876 4586 6888
rect 4706 6876 4712 6888
rect 4764 6916 4770 6928
rect 8202 6916 8208 6928
rect 4764 6888 8208 6916
rect 4764 6876 4770 6888
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 11054 6876 11060 6928
rect 11112 6916 11118 6928
rect 11112 6888 15884 6916
rect 11112 6876 11118 6888
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 7193 6851 7251 6857
rect 2004 6820 6040 6848
rect 2004 6808 2010 6820
rect 6012 6792 6040 6820
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 8846 6848 8852 6860
rect 7239 6820 8852 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 9232 6820 9536 6848
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 4522 6780 4528 6792
rect 4483 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 5442 6780 5448 6792
rect 4847 6752 5448 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5994 6780 6000 6792
rect 5907 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6104 6752 7113 6780
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2648 6684 2697 6712
rect 2648 6672 2654 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 3510 6672 3516 6724
rect 3568 6712 3574 6724
rect 6104 6712 6132 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7282 6780 7288 6792
rect 7243 6752 7288 6780
rect 7101 6743 7159 6749
rect 3568 6684 6132 6712
rect 3568 6672 3574 6684
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 2885 6647 2943 6653
rect 2885 6644 2897 6647
rect 2832 6616 2897 6644
rect 2832 6604 2838 6616
rect 2885 6613 2897 6616
rect 2931 6613 2943 6647
rect 2885 6607 2943 6613
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 4798 6644 4804 6656
rect 3099 6616 4804 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 6822 6644 6828 6656
rect 6783 6616 6828 6644
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7116 6644 7144 6743
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7524 6752 7573 6780
rect 7524 6740 7530 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 9232 6780 9260 6820
rect 9508 6789 9536 6820
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 13872 6820 14289 6848
rect 13872 6808 13878 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 14516 6820 14565 6848
rect 14516 6808 14522 6820
rect 14553 6817 14565 6820
rect 14599 6848 14611 6851
rect 14734 6848 14740 6860
rect 14599 6820 14740 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 15856 6857 15884 6888
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6848 15899 6851
rect 17126 6848 17132 6860
rect 15887 6820 17132 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 8260 6752 9260 6780
rect 9309 6783 9367 6789
rect 8260 6740 8266 6752
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 10042 6780 10048 6792
rect 9955 6752 10048 6780
rect 9493 6743 9551 6749
rect 9324 6712 9352 6743
rect 10042 6740 10048 6752
rect 10100 6780 10106 6792
rect 10686 6780 10692 6792
rect 10100 6752 10692 6780
rect 10100 6740 10106 6752
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16117 6783 16175 6789
rect 16117 6780 16129 6783
rect 15988 6752 16129 6780
rect 15988 6740 15994 6752
rect 16117 6749 16129 6752
rect 16163 6780 16175 6783
rect 16482 6780 16488 6792
rect 16163 6752 16488 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6780 17463 6783
rect 17862 6780 17868 6792
rect 17451 6752 17868 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 10312 6715 10370 6721
rect 9324 6684 9536 6712
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 7116 6616 9413 6644
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9508 6644 9536 6684
rect 10312 6681 10324 6715
rect 10358 6712 10370 6715
rect 10410 6712 10416 6724
rect 10358 6684 10416 6712
rect 10358 6681 10370 6684
rect 10312 6675 10370 6681
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 10502 6644 10508 6656
rect 9508 6616 10508 6644
rect 9401 6607 9459 6613
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10652 6616 11437 6644
rect 10652 6604 10658 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 3326 6440 3332 6452
rect 3287 6412 3332 6440
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 7190 6440 7196 6452
rect 7151 6412 7196 6440
rect 7190 6400 7196 6412
rect 7248 6440 7254 6452
rect 8202 6440 8208 6452
rect 7248 6412 8208 6440
rect 7248 6400 7254 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 10781 6443 10839 6449
rect 10781 6409 10793 6443
rect 10827 6440 10839 6443
rect 10870 6440 10876 6452
rect 10827 6412 10876 6440
rect 10827 6409 10839 6412
rect 10781 6403 10839 6409
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 11848 6412 14473 6440
rect 11848 6400 11854 6412
rect 14461 6409 14473 6412
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 14642 6400 14648 6452
rect 14700 6400 14706 6452
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14792 6412 14841 6440
rect 14792 6400 14798 6412
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6409 16911 6443
rect 43806 6440 43812 6452
rect 16853 6403 16911 6409
rect 18340 6412 43812 6440
rect 2777 6375 2835 6381
rect 2777 6341 2789 6375
rect 2823 6372 2835 6375
rect 3697 6375 3755 6381
rect 3697 6372 3709 6375
rect 2823 6344 3709 6372
rect 2823 6341 2835 6344
rect 2777 6335 2835 6341
rect 3697 6341 3709 6344
rect 3743 6341 3755 6375
rect 3697 6335 3755 6341
rect 5994 6332 6000 6384
rect 6052 6372 6058 6384
rect 7101 6375 7159 6381
rect 7101 6372 7113 6375
rect 6052 6344 7113 6372
rect 6052 6332 6058 6344
rect 7101 6341 7113 6344
rect 7147 6341 7159 6375
rect 11330 6372 11336 6384
rect 7101 6335 7159 6341
rect 10612 6344 11336 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6273 1455 6307
rect 2682 6304 2688 6316
rect 2643 6276 2688 6304
rect 1397 6267 1455 6273
rect 1412 6168 1440 6267
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 3602 6264 3608 6316
rect 3660 6304 3666 6316
rect 3789 6307 3847 6313
rect 3789 6304 3801 6307
rect 3660 6276 3801 6304
rect 3660 6264 3666 6276
rect 3789 6273 3801 6276
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 10042 6304 10048 6316
rect 6788 6276 10048 6304
rect 6788 6264 6794 6276
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 10612 6313 10640 6344
rect 11330 6332 11336 6344
rect 11388 6372 11394 6384
rect 11698 6372 11704 6384
rect 11388 6344 11704 6372
rect 11388 6332 11394 6344
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 14185 6375 14243 6381
rect 14185 6341 14197 6375
rect 14231 6372 14243 6375
rect 14660 6372 14688 6400
rect 16868 6372 16896 6403
rect 17742 6375 17800 6381
rect 17742 6372 17754 6375
rect 14231 6344 14964 6372
rect 16868 6344 17754 6372
rect 14231 6341 14243 6344
rect 14185 6335 14243 6341
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10870 6304 10876 6316
rect 10831 6276 10876 6304
rect 10597 6267 10655 6273
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 14936 6313 14964 6344
rect 17742 6341 17754 6344
rect 17788 6341 17800 6375
rect 17742 6335 17800 6341
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14516 6276 14657 6304
rect 14516 6264 14522 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16448 6276 17049 6304
rect 16448 6264 16454 6276
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 18340 6304 18368 6412
rect 43806 6400 43812 6412
rect 43864 6400 43870 6452
rect 45278 6372 45284 6384
rect 17037 6267 17095 6273
rect 17420 6276 18368 6304
rect 18524 6344 45284 6372
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 7558 6236 7564 6248
rect 1728 6208 7564 6236
rect 1728 6196 1734 6208
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 17420 6236 17448 6276
rect 14608 6208 17448 6236
rect 17497 6239 17555 6245
rect 14608 6196 14614 6208
rect 17497 6205 17509 6239
rect 17543 6205 17555 6239
rect 17497 6199 17555 6205
rect 10686 6168 10692 6180
rect 1412 6140 10692 6168
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 13078 6128 13084 6180
rect 13136 6168 13142 6180
rect 16942 6168 16948 6180
rect 13136 6140 16948 6168
rect 13136 6128 13142 6140
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 17034 6128 17040 6180
rect 17092 6168 17098 6180
rect 17512 6168 17540 6199
rect 17092 6140 17540 6168
rect 17092 6128 17098 6140
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 5350 6100 5356 6112
rect 2740 6072 5356 6100
rect 2740 6060 2746 6072
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 18524 6100 18552 6344
rect 45278 6332 45284 6344
rect 45336 6332 45342 6384
rect 18874 6100 18880 6112
rect 13688 6072 18552 6100
rect 18835 6072 18880 6100
rect 13688 6060 13694 6072
rect 18874 6060 18880 6072
rect 18932 6060 18938 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 13504 5868 14289 5896
rect 13504 5856 13510 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 15197 5899 15255 5905
rect 15197 5896 15209 5899
rect 15160 5868 15209 5896
rect 15160 5856 15166 5868
rect 15197 5865 15209 5868
rect 15243 5865 15255 5899
rect 16390 5896 16396 5908
rect 16351 5868 16396 5896
rect 15197 5859 15255 5865
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 15654 5788 15660 5840
rect 15712 5828 15718 5840
rect 17589 5831 17647 5837
rect 17589 5828 17601 5831
rect 15712 5800 17601 5828
rect 15712 5788 15718 5800
rect 17589 5797 17601 5800
rect 17635 5797 17647 5831
rect 17589 5791 17647 5797
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3418 5760 3424 5772
rect 3099 5732 3424 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3418 5720 3424 5732
rect 3476 5760 3482 5772
rect 3602 5760 3608 5772
rect 3476 5732 3608 5760
rect 3476 5720 3482 5732
rect 3602 5720 3608 5732
rect 3660 5720 3666 5772
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 7616 5732 16865 5760
rect 7616 5720 7622 5732
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17000 5732 17045 5760
rect 17000 5720 17006 5732
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1544 5664 1593 5692
rect 1544 5652 1550 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 6638 5692 6644 5704
rect 6595 5664 6644 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 6822 5701 6828 5704
rect 6816 5692 6828 5701
rect 6783 5664 6828 5692
rect 6816 5655 6828 5664
rect 6822 5652 6828 5655
rect 6880 5652 6886 5704
rect 14458 5692 14464 5704
rect 14371 5664 14464 5692
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15010 5692 15016 5704
rect 14783 5664 15016 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5692 15715 5695
rect 16022 5692 16028 5704
rect 15703 5664 16028 5692
rect 15703 5661 15715 5664
rect 15657 5655 15715 5661
rect 2869 5627 2927 5633
rect 2869 5624 2881 5627
rect 1412 5596 2881 5624
rect 1412 5565 1440 5596
rect 2869 5593 2881 5596
rect 2915 5593 2927 5627
rect 14476 5624 14504 5652
rect 15396 5624 15424 5655
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 16132 5664 17785 5692
rect 16132 5624 16160 5664
rect 17773 5661 17785 5664
rect 17819 5692 17831 5695
rect 17862 5692 17868 5704
rect 17819 5664 17868 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 19058 5692 19064 5704
rect 18095 5664 19064 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 19058 5652 19064 5664
rect 19116 5652 19122 5704
rect 17957 5627 18015 5633
rect 17957 5624 17969 5627
rect 14476 5596 16160 5624
rect 17052 5596 17969 5624
rect 2869 5587 2927 5593
rect 17052 5568 17080 5596
rect 17957 5593 17969 5596
rect 18003 5624 18015 5627
rect 18874 5624 18880 5636
rect 18003 5596 18880 5624
rect 18003 5593 18015 5596
rect 17957 5587 18015 5593
rect 18874 5584 18880 5596
rect 18932 5584 18938 5636
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5525 1455 5559
rect 1397 5519 1455 5525
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 2590 5556 2596 5568
rect 2455 5528 2596 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 3602 5556 3608 5568
rect 2823 5528 3608 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 7834 5556 7840 5568
rect 7340 5528 7840 5556
rect 7340 5516 7346 5528
rect 7834 5516 7840 5528
rect 7892 5556 7898 5568
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 7892 5528 7941 5556
rect 7892 5516 7898 5528
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 7929 5519 7987 5525
rect 14645 5559 14703 5565
rect 14645 5525 14657 5559
rect 14691 5556 14703 5559
rect 14734 5556 14740 5568
rect 14691 5528 14740 5556
rect 14691 5525 14703 5528
rect 14645 5519 14703 5525
rect 14734 5516 14740 5528
rect 14792 5556 14798 5568
rect 15565 5559 15623 5565
rect 15565 5556 15577 5559
rect 14792 5528 15577 5556
rect 14792 5516 14798 5528
rect 15565 5525 15577 5528
rect 15611 5525 15623 5559
rect 15565 5519 15623 5525
rect 16761 5559 16819 5565
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 17034 5556 17040 5568
rect 16807 5528 17040 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 3602 5352 3608 5364
rect 3563 5324 3608 5352
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 10744 5324 12909 5352
rect 10744 5312 10750 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 14461 5355 14519 5361
rect 14461 5352 14473 5355
rect 13320 5324 14473 5352
rect 13320 5312 13326 5324
rect 14461 5321 14473 5324
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14792 5324 14841 5352
rect 14792 5312 14798 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 14829 5315 14887 5321
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 15896 5324 16681 5352
rect 15896 5312 15902 5324
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 18601 5355 18659 5361
rect 18601 5352 18613 5355
rect 17644 5324 18613 5352
rect 17644 5312 17650 5324
rect 18601 5321 18613 5324
rect 18647 5321 18659 5355
rect 18601 5315 18659 5321
rect 3234 5284 3240 5296
rect 2240 5256 3240 5284
rect 2240 5225 2268 5256
rect 3234 5244 3240 5256
rect 3292 5244 3298 5296
rect 18969 5287 19027 5293
rect 18969 5253 18981 5287
rect 19015 5284 19027 5287
rect 19426 5284 19432 5296
rect 19015 5256 19432 5284
rect 19015 5253 19027 5256
rect 18969 5247 19027 5253
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 2498 5225 2504 5228
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2492 5179 2504 5225
rect 2556 5216 2562 5228
rect 2556 5188 2592 5216
rect 2498 5176 2504 5179
rect 2556 5176 2562 5188
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 3568 5188 4261 5216
rect 3568 5176 3574 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5442 5216 5448 5228
rect 4939 5188 5448 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 5442 5176 5448 5188
rect 5500 5216 5506 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 5500 5188 6561 5216
rect 5500 5176 5506 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 6549 5179 6607 5185
rect 9766 5176 9772 5188
rect 9824 5216 9830 5228
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 9824 5188 10609 5216
rect 9824 5176 9830 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10744 5188 10789 5216
rect 10744 5176 10750 5188
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11773 5219 11831 5225
rect 11773 5216 11785 5219
rect 11204 5188 11785 5216
rect 11204 5176 11210 5188
rect 11773 5185 11785 5188
rect 11819 5185 11831 5219
rect 11773 5179 11831 5185
rect 14458 5176 14464 5228
rect 14516 5216 14522 5228
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 14516 5188 14657 5216
rect 14516 5176 14522 5188
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15102 5216 15108 5228
rect 14967 5188 15108 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 17034 5216 17040 5228
rect 16995 5188 17040 5216
rect 16853 5179 16911 5185
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 4709 5151 4767 5157
rect 4709 5148 4721 5151
rect 3844 5120 4721 5148
rect 3844 5108 3850 5120
rect 4709 5117 4721 5120
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5224 5120 6377 5148
rect 5224 5108 5230 5120
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 9950 5148 9956 5160
rect 9907 5120 9956 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 10836 5120 11529 5148
rect 10836 5108 10842 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 16868 5148 16896 5179
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 17184 5188 17229 5216
rect 17184 5176 17190 5188
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18564 5188 18797 5216
rect 18564 5176 18570 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 19061 5219 19119 5225
rect 19061 5185 19073 5219
rect 19107 5216 19119 5219
rect 30282 5216 30288 5228
rect 19107 5188 30288 5216
rect 19107 5185 19119 5188
rect 19061 5179 19119 5185
rect 30282 5176 30288 5188
rect 30340 5176 30346 5228
rect 18524 5148 18552 5176
rect 16868 5120 18552 5148
rect 11517 5111 11575 5117
rect 4065 5083 4123 5089
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 6822 5080 6828 5092
rect 4111 5052 6828 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 10502 5080 10508 5092
rect 9968 5052 10508 5080
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 3142 5012 3148 5024
rect 1627 4984 3148 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5718 5012 5724 5024
rect 5123 4984 5724 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6730 5012 6736 5024
rect 6691 4984 6736 5012
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 9968 5021 9996 5052
rect 10502 5040 10508 5052
rect 10560 5080 10566 5092
rect 10560 5052 10640 5080
rect 10560 5040 10566 5052
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 4981 10011 5015
rect 10134 5012 10140 5024
rect 10095 4984 10140 5012
rect 9953 4975 10011 4981
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10612 5021 10640 5052
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 4981 10655 5015
rect 10597 4975 10655 4981
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 11514 5012 11520 5024
rect 11011 4984 11520 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2498 4808 2504 4820
rect 2455 4780 2504 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 4614 4808 4620 4820
rect 4575 4780 4620 4808
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 6730 4768 6736 4820
rect 6788 4808 6794 4820
rect 11146 4808 11152 4820
rect 6788 4780 9904 4808
rect 11107 4780 11152 4808
rect 6788 4768 6794 4780
rect 9876 4740 9904 4780
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 15381 4811 15439 4817
rect 15381 4808 15393 4811
rect 14240 4780 15393 4808
rect 14240 4768 14246 4780
rect 15381 4777 15393 4780
rect 15427 4777 15439 4811
rect 15381 4771 15439 4777
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 18233 4811 18291 4817
rect 18233 4808 18245 4811
rect 17828 4780 18245 4808
rect 17828 4768 17834 4780
rect 18233 4777 18245 4780
rect 18279 4777 18291 4811
rect 18233 4771 18291 4777
rect 9876 4712 24624 4740
rect 3602 4632 3608 4684
rect 3660 4672 3666 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3660 4644 3801 4672
rect 3660 4632 3666 4644
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 5442 4672 5448 4684
rect 3789 4635 3847 4641
rect 3988 4644 5448 4672
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 2590 4604 2596 4616
rect 2551 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3234 4604 3240 4616
rect 3147 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4604 3298 4616
rect 3510 4604 3516 4616
rect 3292 4576 3516 4604
rect 3292 4564 3298 4576
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 3988 4613 4016 4644
rect 5442 4632 5448 4644
rect 5500 4672 5506 4684
rect 5500 4644 6408 4672
rect 5500 4632 5506 4644
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 6380 4613 6408 4644
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 17092 4644 19257 4672
rect 17092 4632 17098 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4764 4576 4813 4604
rect 4764 4564 4770 4576
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 10778 4604 10784 4616
rect 8987 4576 10784 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 3878 4496 3884 4548
rect 3936 4536 3942 4548
rect 6196 4536 6224 4567
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 11330 4604 11336 4616
rect 11291 4576 11336 4604
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 15565 4607 15623 4613
rect 15565 4573 15577 4607
rect 15611 4573 15623 4607
rect 15838 4604 15844 4616
rect 15799 4576 15844 4604
rect 15565 4567 15623 4573
rect 3936 4508 6224 4536
rect 9208 4539 9266 4545
rect 3936 4496 3942 4508
rect 9208 4505 9220 4539
rect 9254 4536 9266 4539
rect 9766 4536 9772 4548
rect 9254 4508 9772 4536
rect 9254 4505 9266 4508
rect 9208 4499 9266 4505
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 11514 4536 11520 4548
rect 11475 4508 11520 4536
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 15580 4536 15608 4567
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 16482 4604 16488 4616
rect 16347 4576 16488 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4604 16635 4607
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 16623 4576 18429 4604
rect 16623 4573 16635 4576
rect 16577 4567 16635 4573
rect 18417 4573 18429 4576
rect 18463 4604 18475 4607
rect 18506 4604 18512 4616
rect 18463 4576 18512 4604
rect 18463 4573 18475 4576
rect 18417 4567 18475 4573
rect 16592 4536 16620 4567
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 24596 4613 24624 4712
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4573 18751 4607
rect 18693 4567 18751 4573
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 15580 4508 16620 4536
rect 18708 4536 18736 4567
rect 28810 4536 28816 4548
rect 18708 4508 28816 4536
rect 28810 4496 28816 4508
rect 28868 4496 28874 4548
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 4154 4468 4160 4480
rect 4115 4440 4160 4468
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4468 6607 4471
rect 8202 4468 8208 4480
rect 6595 4440 8208 4468
rect 6595 4437 6607 4440
rect 6549 4431 6607 4437
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10321 4471 10379 4477
rect 10321 4468 10333 4471
rect 10008 4440 10333 4468
rect 10008 4428 10014 4440
rect 10321 4437 10333 4440
rect 10367 4437 10379 4471
rect 10321 4431 10379 4437
rect 15749 4471 15807 4477
rect 15749 4437 15761 4471
rect 15795 4468 15807 4471
rect 17034 4468 17040 4480
rect 15795 4440 17040 4468
rect 15795 4437 15807 4440
rect 15749 4431 15807 4437
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 18690 4468 18696 4480
rect 18647 4440 18696 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 18690 4428 18696 4440
rect 18748 4468 18754 4480
rect 19426 4468 19432 4480
rect 18748 4440 19432 4468
rect 18748 4428 18754 4440
rect 19426 4428 19432 4440
rect 19484 4477 19490 4480
rect 19484 4471 19533 4477
rect 19484 4437 19487 4471
rect 19521 4437 19533 4471
rect 19484 4431 19533 4437
rect 24397 4471 24455 4477
rect 24397 4437 24409 4471
rect 24443 4468 24455 4471
rect 24670 4468 24676 4480
rect 24443 4440 24676 4468
rect 24443 4437 24455 4440
rect 24397 4431 24455 4437
rect 19484 4428 19490 4431
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 9950 4264 9956 4276
rect 1452 4236 9956 4264
rect 1452 4224 1458 4236
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10134 4264 10140 4276
rect 10095 4236 10140 4264
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 19426 4264 19432 4276
rect 18564 4236 19432 4264
rect 18564 4224 18570 4236
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 2130 4156 2136 4208
rect 2188 4196 2194 4208
rect 2225 4199 2283 4205
rect 2225 4196 2237 4199
rect 2188 4168 2237 4196
rect 2188 4156 2194 4168
rect 2225 4165 2237 4168
rect 2271 4165 2283 4199
rect 2225 4159 2283 4165
rect 3510 4156 3516 4208
rect 3568 4196 3574 4208
rect 3568 4168 3924 4196
rect 3568 4156 3574 4168
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 3418 4128 3424 4140
rect 1443 4100 2774 4128
rect 3379 4100 3424 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 2746 3992 2774 4100
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 3620 4060 3648 4091
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 3896 4128 3924 4168
rect 4540 4168 5120 4196
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 3752 4100 3797 4128
rect 3896 4100 4353 4128
rect 3752 4088 3758 4100
rect 4341 4097 4353 4100
rect 4387 4128 4399 4131
rect 4540 4128 4568 4168
rect 4387 4100 4568 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4614 4088 4620 4140
rect 4672 4128 4678 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4672 4100 4997 4128
rect 4672 4088 4678 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 5092 4128 5120 4168
rect 5258 4156 5264 4208
rect 5316 4196 5322 4208
rect 6733 4199 6791 4205
rect 5316 4168 5856 4196
rect 5316 4156 5322 4168
rect 5442 4128 5448 4140
rect 5092 4100 5448 4128
rect 4985 4091 5043 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5166 4060 5172 4072
rect 2924 4032 5172 4060
rect 2924 4020 2930 4032
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 5828 4060 5856 4168
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 8018 4196 8024 4208
rect 6779 4168 8024 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 8018 4156 8024 4168
rect 8076 4156 8082 4208
rect 19705 4199 19763 4205
rect 19705 4196 19717 4199
rect 18800 4168 19717 4196
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 9766 4128 9772 4140
rect 6880 4100 6925 4128
rect 9727 4100 9772 4128
rect 6880 4088 6886 4100
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4128 10287 4131
rect 10410 4128 10416 4140
rect 10275 4100 10416 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 5408 4032 5488 4060
rect 5828 4032 6929 4060
rect 5408 4020 5414 4032
rect 3694 3992 3700 4004
rect 2746 3964 3700 3992
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 5460 4001 5488 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 9968 4060 9996 4091
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16206 4128 16212 4140
rect 16163 4100 16212 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 16206 4088 16212 4100
rect 16264 4088 16270 4140
rect 18414 4128 18420 4140
rect 18375 4100 18420 4128
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 18598 4128 18604 4140
rect 18559 4100 18604 4128
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 18800 4137 18828 4168
rect 19705 4165 19717 4168
rect 19751 4165 19763 4199
rect 19705 4159 19763 4165
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18748 4100 18797 4128
rect 18748 4088 18754 4100
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4097 18935 4131
rect 19334 4128 19340 4140
rect 19295 4100 19340 4128
rect 18877 4091 18935 4097
rect 11330 4060 11336 4072
rect 9968 4032 11336 4060
rect 6917 4023 6975 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16540 4032 16681 4060
rect 16540 4020 16546 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 16945 4063 17003 4069
rect 16945 4029 16957 4063
rect 16991 4060 17003 4063
rect 18616 4060 18644 4088
rect 16991 4032 18644 4060
rect 18892 4060 18920 4091
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 19484 4100 19533 4128
rect 19484 4088 19490 4100
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 19521 4091 19579 4097
rect 19797 4131 19855 4137
rect 19797 4097 19809 4131
rect 19843 4128 19855 4131
rect 23014 4128 23020 4140
rect 19843 4100 23020 4128
rect 19843 4097 19855 4100
rect 19797 4091 19855 4097
rect 23014 4088 23020 4100
rect 23072 4088 23078 4140
rect 26050 4060 26056 4072
rect 18892 4032 26056 4060
rect 16991 4029 17003 4032
rect 16945 4023 17003 4029
rect 26050 4020 26056 4032
rect 26108 4020 26114 4072
rect 5445 3995 5503 4001
rect 5445 3961 5457 3995
rect 5491 3961 5503 3995
rect 5445 3955 5503 3961
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 11020 3964 16896 3992
rect 11020 3952 11026 3964
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2958 3924 2964 3936
rect 1627 3896 2964 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3878 3924 3884 3936
rect 3283 3896 3884 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4028 3896 4169 3924
rect 4028 3884 4034 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4798 3924 4804 3936
rect 4759 3896 4804 3924
rect 4157 3887 4215 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 6365 3927 6423 3933
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 6454 3924 6460 3936
rect 6411 3896 6460 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 14918 3884 14924 3936
rect 14976 3924 14982 3936
rect 15933 3927 15991 3933
rect 15933 3924 15945 3927
rect 14976 3896 15945 3924
rect 14976 3884 14982 3896
rect 15933 3893 15945 3896
rect 15979 3893 15991 3927
rect 16868 3924 16896 3964
rect 17126 3952 17132 4004
rect 17184 3992 17190 4004
rect 33686 3992 33692 4004
rect 17184 3964 33692 3992
rect 17184 3952 17190 3964
rect 33686 3952 33692 3964
rect 33744 3952 33750 4004
rect 21266 3924 21272 3936
rect 16868 3896 21272 3924
rect 15933 3887 15991 3893
rect 21266 3884 21272 3896
rect 21324 3884 21330 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 2682 3680 2688 3732
rect 2740 3720 2746 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 2740 3692 5641 3720
rect 2740 3680 2746 3692
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 5629 3683 5687 3689
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 10870 3720 10876 3732
rect 10735 3692 10876 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 16574 3720 16580 3732
rect 16535 3692 16580 3720
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 17494 3680 17500 3732
rect 17552 3720 17558 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 17552 3692 18245 3720
rect 17552 3680 17558 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 19150 3680 19156 3732
rect 19208 3720 19214 3732
rect 23750 3720 23756 3732
rect 19208 3692 23756 3720
rect 19208 3680 19214 3692
rect 23750 3680 23756 3692
rect 23808 3680 23814 3732
rect 5166 3652 5172 3664
rect 5127 3624 5172 3652
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 6638 3652 6644 3664
rect 5500 3624 6644 3652
rect 5500 3612 5506 3624
rect 6638 3612 6644 3624
rect 6696 3612 6702 3664
rect 10778 3652 10784 3664
rect 9508 3624 10784 3652
rect 3050 3584 3056 3596
rect 1412 3556 3056 3584
rect 1412 3525 1440 3556
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3568 3556 3801 3584
rect 3568 3544 3574 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 9508 3584 9536 3624
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 15562 3652 15568 3664
rect 14384 3624 15568 3652
rect 4856 3556 9536 3584
rect 4856 3544 4862 3556
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 14384 3584 14412 3624
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 16114 3612 16120 3664
rect 16172 3652 16178 3664
rect 57977 3655 58035 3661
rect 57977 3652 57989 3655
rect 16172 3624 57989 3652
rect 16172 3612 16178 3624
rect 57977 3621 57989 3624
rect 58023 3621 58035 3655
rect 57977 3615 58035 3621
rect 9640 3556 14412 3584
rect 14645 3587 14703 3593
rect 9640 3544 9646 3556
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 16482 3584 16488 3596
rect 14691 3556 16488 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 23658 3584 23664 3596
rect 17052 3556 23664 3584
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 2179 3488 2774 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 2746 3448 2774 3488
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 2924 3488 2969 3516
rect 2924 3476 2930 3488
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4045 3519 4103 3525
rect 4045 3516 4057 3519
rect 3936 3488 4057 3516
rect 3936 3476 3942 3488
rect 4045 3485 4057 3488
rect 4091 3485 4103 3519
rect 4045 3479 4103 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 5813 3479 5871 3485
rect 2746 3420 3188 3448
rect 198 3340 204 3392
rect 256 3380 262 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 256 3352 1593 3380
rect 256 3340 262 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 2317 3383 2375 3389
rect 2317 3380 2329 3383
rect 1728 3352 2329 3380
rect 1728 3340 1734 3352
rect 2317 3349 2329 3352
rect 2363 3349 2375 3383
rect 2317 3343 2375 3349
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 2832 3352 3065 3380
rect 2832 3340 2838 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3160 3380 3188 3420
rect 3234 3408 3240 3460
rect 3292 3448 3298 3460
rect 5828 3448 5856 3479
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6604 3488 7113 3516
rect 6604 3476 6610 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7524 3488 7757 3516
rect 7524 3476 7530 3488
rect 7745 3485 7757 3488
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10318 3516 10324 3528
rect 10275 3488 10324 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3516 10931 3519
rect 10962 3516 10968 3528
rect 10919 3488 10968 3516
rect 10919 3485 10931 3488
rect 10873 3479 10931 3485
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 7834 3448 7840 3460
rect 3292 3420 5856 3448
rect 6104 3420 7840 3448
rect 3292 3408 3298 3420
rect 3602 3380 3608 3392
rect 3160 3352 3608 3380
rect 3053 3343 3111 3349
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 6104 3380 6132 3420
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 11164 3448 11192 3479
rect 11330 3476 11336 3528
rect 11388 3516 11394 3528
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 11388 3488 11805 3516
rect 11388 3476 11394 3488
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13412 3488 13553 3516
rect 13412 3476 13418 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14792 3488 14933 3516
rect 14792 3476 14798 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 17052 3525 17080 3556
rect 23658 3544 23664 3556
rect 23716 3544 23722 3596
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15344 3488 16129 3516
rect 15344 3476 15350 3488
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 10060 3420 11192 3448
rect 6270 3380 6276 3392
rect 3752 3352 6132 3380
rect 6231 3352 6276 3380
rect 3752 3340 3758 3352
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 7558 3380 7564 3392
rect 7519 3352 7564 3380
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 10060 3389 10088 3420
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 14752 3448 14780 3476
rect 16776 3448 16804 3479
rect 17678 3476 17684 3528
rect 17736 3516 17742 3528
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17736 3488 17785 3516
rect 17736 3476 17742 3488
rect 17773 3485 17785 3488
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18598 3516 18604 3528
rect 18463 3488 18604 3516
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 16850 3448 16856 3460
rect 12768 3420 14780 3448
rect 16763 3420 16856 3448
rect 12768 3408 12774 3420
rect 16850 3408 16856 3420
rect 16908 3448 16914 3460
rect 17954 3448 17960 3460
rect 16908 3420 17960 3448
rect 16908 3408 16914 3420
rect 17954 3408 17960 3420
rect 18012 3448 18018 3460
rect 18432 3448 18460 3479
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 18012 3420 18460 3448
rect 18708 3448 18736 3479
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18840 3488 19441 3516
rect 18840 3476 18846 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21361 3519 21419 3525
rect 21361 3516 21373 3519
rect 21140 3488 21373 3516
rect 21140 3476 21146 3488
rect 21361 3485 21373 3488
rect 21407 3485 21419 3519
rect 21361 3479 21419 3485
rect 22462 3448 22468 3460
rect 18708 3420 22468 3448
rect 18012 3408 18018 3420
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 57793 3451 57851 3457
rect 57793 3417 57805 3451
rect 57839 3448 57851 3451
rect 59630 3448 59636 3460
rect 57839 3420 59636 3448
rect 57839 3417 57851 3420
rect 57793 3411 57851 3417
rect 59630 3408 59636 3420
rect 59688 3408 59694 3460
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3349 10103 3383
rect 10045 3343 10103 3349
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10836 3352 11069 3380
rect 10836 3340 10842 3352
rect 11057 3349 11069 3352
rect 11103 3380 11115 3383
rect 12434 3380 12440 3392
rect 11103 3352 12440 3380
rect 11103 3349 11115 3352
rect 11057 3343 11115 3349
rect 12434 3340 12440 3352
rect 12492 3340 12498 3392
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 13044 3352 13369 3380
rect 13044 3340 13050 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 16942 3380 16948 3392
rect 16903 3352 16948 3380
rect 13357 3343 13415 3349
rect 16942 3340 16948 3352
rect 17000 3380 17006 3392
rect 18046 3380 18052 3392
rect 17000 3352 18052 3380
rect 17000 3340 17006 3352
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18601 3383 18659 3389
rect 18601 3349 18613 3383
rect 18647 3380 18659 3383
rect 18690 3380 18696 3392
rect 18647 3352 18696 3380
rect 18647 3349 18659 3352
rect 18601 3343 18659 3349
rect 18690 3340 18696 3352
rect 18748 3340 18754 3392
rect 19242 3380 19248 3392
rect 19203 3352 19248 3380
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 21174 3380 21180 3392
rect 21135 3352 21180 3380
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 3602 3136 3608 3188
rect 3660 3176 3666 3188
rect 4890 3176 4896 3188
rect 3660 3148 4896 3176
rect 3660 3136 3666 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8018 3176 8024 3188
rect 7975 3148 8024 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 10410 3176 10416 3188
rect 10371 3148 10416 3176
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 10778 3176 10784 3188
rect 10739 3148 10784 3176
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 11606 3176 11612 3188
rect 11563 3148 11612 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12434 3176 12440 3188
rect 11931 3148 12440 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12434 3136 12440 3148
rect 12492 3176 12498 3188
rect 13446 3176 13452 3188
rect 12492 3148 13452 3176
rect 12492 3136 12498 3148
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14424 3148 14473 3176
rect 14424 3136 14430 3148
rect 14461 3145 14473 3148
rect 14507 3145 14519 3179
rect 16942 3176 16948 3188
rect 14461 3139 14519 3145
rect 15028 3148 16948 3176
rect 3970 3108 3976 3120
rect 2700 3080 3976 3108
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 1946 3040 1952 3052
rect 1719 3012 1952 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2700 3049 2728 3080
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 5626 3108 5632 3120
rect 4120 3080 5632 3108
rect 4120 3068 4126 3080
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 6270 3068 6276 3120
rect 6328 3108 6334 3120
rect 6794 3111 6852 3117
rect 6794 3108 6806 3111
rect 6328 3080 6806 3108
rect 6328 3068 6334 3080
rect 6794 3077 6806 3080
rect 6840 3077 6852 3111
rect 6794 3071 6852 3077
rect 7558 3068 7564 3120
rect 7616 3108 7622 3120
rect 15028 3108 15056 3148
rect 16942 3136 16948 3148
rect 17000 3176 17006 3188
rect 17129 3179 17187 3185
rect 17129 3176 17141 3179
rect 17000 3148 17141 3176
rect 17000 3136 17006 3148
rect 17129 3145 17141 3148
rect 17175 3145 17187 3179
rect 19242 3176 19248 3188
rect 17129 3139 17187 3145
rect 17308 3148 19248 3176
rect 7616 3080 12020 3108
rect 7616 3068 7622 3080
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 4154 3040 4160 3052
rect 3743 3012 4160 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 5718 3040 5724 3052
rect 5679 3012 5724 3040
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6638 3040 6644 3052
rect 6595 3012 6644 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8573 3043 8631 3049
rect 8573 3040 8585 3043
rect 8260 3012 8585 3040
rect 8260 3000 8266 3012
rect 8573 3009 8585 3012
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9364 3012 9965 3040
rect 9364 3000 9370 3012
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 10597 3003 10655 3009
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 2648 2944 4353 2972
rect 2648 2932 2654 2944
rect 4341 2941 4353 2944
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 10612 2972 10640 3003
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11992 3049 12020 3080
rect 13188 3080 15056 3108
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 10962 2972 10968 2984
rect 8076 2944 9168 2972
rect 10612 2944 10968 2972
rect 8076 2932 8082 2944
rect 3602 2864 3608 2916
rect 3660 2904 3666 2916
rect 4985 2907 5043 2913
rect 4985 2904 4997 2907
rect 3660 2876 4997 2904
rect 3660 2864 3666 2876
rect 4985 2873 4997 2876
rect 5031 2873 5043 2907
rect 4985 2867 5043 2873
rect 8389 2907 8447 2913
rect 8389 2873 8401 2907
rect 8435 2904 8447 2907
rect 9030 2904 9036 2916
rect 8435 2876 9036 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 9140 2904 9168 2944
rect 10962 2932 10968 2944
rect 11020 2972 11026 2984
rect 11716 2972 11744 3003
rect 12710 2972 12716 2984
rect 11020 2944 12716 2972
rect 11020 2932 11026 2944
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 13188 2981 13216 3080
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 16761 3111 16819 3117
rect 16761 3108 16773 3111
rect 16356 3080 16773 3108
rect 16356 3068 16362 3080
rect 16761 3077 16773 3080
rect 16807 3077 16819 3111
rect 16761 3071 16819 3077
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14734 3040 14740 3052
rect 14691 3012 14740 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13446 2972 13452 2984
rect 13359 2944 13452 2972
rect 13173 2935 13231 2941
rect 13188 2904 13216 2935
rect 13446 2932 13452 2944
rect 13504 2972 13510 2984
rect 14844 2972 14872 3003
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 14976 3012 15021 3040
rect 14976 3000 14982 3012
rect 15930 3000 15936 3052
rect 15988 3040 15994 3052
rect 16117 3043 16175 3049
rect 16117 3040 16129 3043
rect 15988 3012 16129 3040
rect 15988 3000 15994 3012
rect 16117 3009 16129 3012
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 16850 3000 16856 3052
rect 16908 3040 16914 3052
rect 16945 3043 17003 3049
rect 16945 3040 16957 3043
rect 16908 3012 16957 3040
rect 16908 3000 16914 3012
rect 16945 3009 16957 3012
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 17221 3044 17279 3049
rect 17308 3044 17336 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 23658 3176 23664 3188
rect 23619 3148 23664 3176
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 56965 3179 57023 3185
rect 56965 3176 56977 3179
rect 23808 3148 56977 3176
rect 23808 3136 23814 3148
rect 56965 3145 56977 3148
rect 57011 3145 57023 3179
rect 56965 3139 57023 3145
rect 17402 3068 17408 3120
rect 17460 3108 17466 3120
rect 17681 3111 17739 3117
rect 17681 3108 17693 3111
rect 17460 3080 17693 3108
rect 17460 3068 17466 3080
rect 17681 3077 17693 3080
rect 17727 3077 17739 3111
rect 18046 3108 18052 3120
rect 18007 3080 18052 3108
rect 17681 3071 17739 3077
rect 18046 3068 18052 3080
rect 18104 3068 18110 3120
rect 21174 3108 21180 3120
rect 18156 3080 21180 3108
rect 17221 3043 17336 3044
rect 17221 3009 17233 3043
rect 17267 3016 17336 3043
rect 17865 3043 17923 3049
rect 17267 3009 17279 3016
rect 17221 3003 17279 3009
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 17954 3040 17960 3052
rect 17911 3012 17960 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 18156 3049 18184 3080
rect 21174 3068 21180 3080
rect 21232 3068 21238 3120
rect 23014 3068 23020 3120
rect 23072 3108 23078 3120
rect 32398 3108 32404 3120
rect 23072 3080 32404 3108
rect 23072 3068 23078 3080
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 19061 3043 19119 3049
rect 19061 3009 19073 3043
rect 19107 3009 19119 3043
rect 21266 3040 21272 3052
rect 21227 3012 21272 3040
rect 19061 3003 19119 3009
rect 13504 2944 14872 2972
rect 13504 2932 13510 2944
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 19076 2972 19104 3003
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 23566 3000 23572 3052
rect 23624 3040 23630 3052
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23624 3012 23857 3040
rect 23624 3000 23630 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 27430 3000 27436 3052
rect 27488 3040 27494 3052
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 27488 3012 27721 3040
rect 27488 3000 27494 3012
rect 27709 3009 27721 3012
rect 27755 3009 27767 3043
rect 33686 3040 33692 3052
rect 33647 3012 33692 3040
rect 27709 3003 27767 3009
rect 33686 3000 33692 3012
rect 33744 3000 33750 3052
rect 56686 3000 56692 3052
rect 56744 3040 56750 3052
rect 56781 3043 56839 3049
rect 56781 3040 56793 3043
rect 56744 3012 56793 3040
rect 56744 3000 56750 3012
rect 56781 3009 56793 3012
rect 56827 3009 56839 3043
rect 56781 3003 56839 3009
rect 15620 2944 19104 2972
rect 15620 2932 15626 2944
rect 22462 2932 22468 2984
rect 22520 2972 22526 2984
rect 22520 2944 26234 2972
rect 22520 2932 22526 2944
rect 9140 2876 13216 2904
rect 15933 2907 15991 2913
rect 15933 2873 15945 2907
rect 15979 2904 15991 2907
rect 17310 2904 17316 2916
rect 15979 2876 17316 2904
rect 15979 2873 15991 2876
rect 15933 2867 15991 2873
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 18877 2907 18935 2913
rect 18877 2873 18889 2907
rect 18923 2904 18935 2907
rect 19610 2904 19616 2916
rect 18923 2876 19616 2904
rect 18923 2873 18935 2876
rect 18877 2867 18935 2873
rect 19610 2864 19616 2876
rect 19668 2864 19674 2916
rect 21085 2907 21143 2913
rect 21085 2873 21097 2907
rect 21131 2904 21143 2907
rect 22186 2904 22192 2916
rect 21131 2876 22192 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 26206 2904 26234 2944
rect 33318 2932 33324 2984
rect 33376 2972 33382 2984
rect 33413 2975 33471 2981
rect 33413 2972 33425 2975
rect 33376 2944 33425 2972
rect 33376 2932 33382 2944
rect 33413 2941 33425 2944
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 27525 2907 27583 2913
rect 27525 2904 27537 2907
rect 26206 2876 27537 2904
rect 27525 2873 27537 2876
rect 27571 2873 27583 2907
rect 27525 2867 27583 2873
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 2869 2839 2927 2845
rect 2869 2836 2881 2839
rect 716 2808 2881 2836
rect 716 2796 722 2808
rect 2869 2805 2881 2808
rect 2915 2805 2927 2839
rect 2869 2799 2927 2805
rect 3513 2839 3571 2845
rect 3513 2805 3525 2839
rect 3559 2836 3571 2839
rect 3786 2836 3792 2848
rect 3559 2808 3792 2836
rect 3559 2805 3571 2808
rect 3513 2799 3571 2805
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 6362 2836 6368 2848
rect 5583 2808 6368 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 9217 2839 9275 2845
rect 9217 2836 9229 2839
rect 8536 2808 9229 2836
rect 8536 2796 8542 2808
rect 9217 2805 9229 2808
rect 9263 2805 9275 2839
rect 9217 2799 9275 2805
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 11790 2836 11796 2848
rect 9815 2808 11796 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 12621 2839 12679 2845
rect 12621 2836 12633 2839
rect 12400 2808 12633 2836
rect 12400 2796 12406 2808
rect 12621 2805 12633 2808
rect 12667 2805 12679 2839
rect 12621 2799 12679 2805
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19705 2839 19763 2845
rect 19705 2836 19717 2839
rect 19208 2808 19717 2836
rect 19208 2796 19214 2808
rect 19705 2805 19717 2808
rect 19751 2805 19763 2839
rect 19705 2799 19763 2805
rect 21634 2796 21640 2848
rect 21692 2836 21698 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21692 2808 22017 2836
rect 21692 2796 21698 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 32306 2796 32312 2848
rect 32364 2836 32370 2848
rect 32585 2839 32643 2845
rect 32585 2836 32597 2839
rect 32364 2808 32597 2836
rect 32364 2796 32370 2808
rect 32585 2805 32597 2808
rect 32631 2805 32643 2839
rect 32585 2799 32643 2805
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35529 2839 35587 2845
rect 35529 2836 35541 2839
rect 35400 2808 35541 2836
rect 35400 2796 35406 2808
rect 35529 2805 35541 2808
rect 35575 2805 35587 2839
rect 35529 2799 35587 2805
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36780 2808 37473 2836
rect 36780 2796 36786 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 39666 2796 39672 2848
rect 39724 2836 39730 2848
rect 39945 2839 40003 2845
rect 39945 2836 39957 2839
rect 39724 2808 39957 2836
rect 39724 2796 39730 2808
rect 39945 2805 39957 2808
rect 39991 2805 40003 2839
rect 39945 2799 40003 2805
rect 42610 2796 42616 2848
rect 42668 2836 42674 2848
rect 42889 2839 42947 2845
rect 42889 2836 42901 2839
rect 42668 2808 42901 2836
rect 42668 2796 42674 2808
rect 42889 2805 42901 2808
rect 42935 2805 42947 2839
rect 42889 2799 42947 2805
rect 44082 2796 44088 2848
rect 44140 2836 44146 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 44140 2808 44373 2836
rect 44140 2796 44146 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 46934 2796 46940 2848
rect 46992 2836 46998 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 46992 2808 47777 2836
rect 46992 2796 46998 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 47765 2799 47823 2805
rect 49878 2796 49884 2848
rect 49936 2836 49942 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49936 2808 50169 2836
rect 49936 2796 49942 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 52822 2796 52828 2848
rect 52880 2836 52886 2848
rect 53101 2839 53159 2845
rect 53101 2836 53113 2839
rect 52880 2808 53113 2836
rect 52880 2796 52886 2808
rect 53101 2805 53113 2808
rect 53147 2805 53159 2839
rect 53101 2799 53159 2805
rect 54294 2796 54300 2848
rect 54352 2836 54358 2848
rect 54573 2839 54631 2845
rect 54573 2836 54585 2839
rect 54352 2808 54585 2836
rect 54352 2796 54358 2808
rect 54573 2805 54585 2808
rect 54619 2805 54631 2839
rect 54573 2799 54631 2805
rect 58161 2839 58219 2845
rect 58161 2805 58173 2839
rect 58207 2836 58219 2839
rect 58710 2836 58716 2848
rect 58207 2808 58716 2836
rect 58207 2805 58219 2808
rect 58161 2799 58219 2805
rect 58710 2796 58716 2808
rect 58768 2796 58774 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 4706 2632 4712 2644
rect 2924 2604 4712 2632
rect 2924 2592 2930 2604
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 12526 2632 12532 2644
rect 12487 2604 12532 2632
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 19794 2632 19800 2644
rect 15528 2604 19800 2632
rect 15528 2592 15534 2604
rect 19794 2592 19800 2604
rect 19852 2592 19858 2644
rect 24946 2632 24952 2644
rect 19996 2604 24952 2632
rect 14093 2567 14151 2573
rect 14093 2533 14105 2567
rect 14139 2533 14151 2567
rect 14093 2527 14151 2533
rect 1118 2456 1124 2508
rect 1176 2496 1182 2508
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 1176 2468 4537 2496
rect 1176 2456 1182 2468
rect 4525 2465 4537 2468
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 5592 2468 7297 2496
rect 5592 2456 5598 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 8386 2456 8392 2508
rect 8444 2496 8450 2508
rect 14108 2496 14136 2527
rect 14274 2524 14280 2576
rect 14332 2564 14338 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 14332 2536 16865 2564
rect 14332 2524 14338 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 19996 2564 20024 2604
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 26050 2632 26056 2644
rect 26011 2604 26056 2632
rect 26050 2592 26056 2604
rect 26108 2592 26114 2644
rect 28810 2632 28816 2644
rect 28771 2604 28816 2632
rect 28810 2592 28816 2604
rect 28868 2592 28874 2644
rect 30282 2632 30288 2644
rect 30243 2604 30288 2632
rect 30282 2592 30288 2604
rect 30340 2592 30346 2644
rect 31018 2592 31024 2644
rect 31076 2632 31082 2644
rect 51169 2635 51227 2641
rect 51169 2632 51181 2635
rect 31076 2604 51181 2632
rect 31076 2592 31082 2604
rect 51169 2601 51181 2604
rect 51215 2601 51227 2635
rect 51169 2595 51227 2601
rect 17828 2536 20024 2564
rect 17828 2524 17834 2536
rect 20070 2524 20076 2576
rect 20128 2564 20134 2576
rect 48225 2567 48283 2573
rect 48225 2564 48237 2567
rect 20128 2536 48237 2564
rect 20128 2524 20134 2536
rect 48225 2533 48237 2536
rect 48271 2533 48283 2567
rect 48225 2527 48283 2533
rect 8444 2468 13124 2496
rect 14108 2468 14964 2496
rect 8444 2456 8450 2468
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 1397 2391 1455 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 6362 2428 6368 2440
rect 6323 2400 6368 2428
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 9030 2428 9036 2440
rect 8991 2400 9036 2428
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9398 2388 9404 2440
rect 9456 2428 9462 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9456 2400 9965 2428
rect 9456 2388 9462 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 11790 2428 11796 2440
rect 11751 2400 11796 2428
rect 9953 2391 10011 2397
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 12710 2428 12716 2440
rect 12671 2400 12716 2428
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 12986 2428 12992 2440
rect 12947 2400 12992 2428
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13096 2428 13124 2468
rect 14936 2437 14964 2468
rect 16758 2456 16764 2508
rect 16816 2496 16822 2508
rect 18233 2499 18291 2505
rect 18233 2496 18245 2499
rect 16816 2468 18245 2496
rect 16816 2456 16822 2468
rect 18233 2465 18245 2468
rect 18279 2465 18291 2499
rect 18233 2459 18291 2465
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 32398 2496 32404 2508
rect 19116 2468 32260 2496
rect 32359 2468 32404 2496
rect 19116 2456 19122 2468
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13096 2400 14289 2428
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2397 14979 2431
rect 17310 2428 17316 2440
rect 17271 2400 17316 2428
rect 14921 2391 14979 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 19610 2388 19616 2440
rect 19668 2428 19674 2440
rect 19797 2431 19855 2437
rect 19797 2428 19809 2431
rect 19668 2400 19809 2428
rect 19668 2388 19674 2400
rect 19797 2397 19809 2400
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 20162 2388 20168 2440
rect 20220 2428 20226 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20220 2400 20729 2428
rect 20220 2388 20226 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 22186 2428 22192 2440
rect 22147 2400 22192 2428
rect 20717 2391 20775 2397
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 23109 2431 23167 2437
rect 23109 2428 23121 2431
rect 22612 2400 23121 2428
rect 22612 2388 22618 2400
rect 23109 2397 23121 2400
rect 23155 2397 23167 2431
rect 23109 2391 23167 2397
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 24026 2428 24032 2440
rect 23891 2400 24032 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 24670 2428 24676 2440
rect 24631 2400 24676 2428
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 25038 2388 25044 2440
rect 25096 2428 25102 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 25096 2400 25605 2428
rect 25096 2388 25102 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 25958 2388 25964 2440
rect 26016 2428 26022 2440
rect 26237 2431 26295 2437
rect 26237 2428 26249 2431
rect 26016 2400 26249 2428
rect 26016 2388 26022 2400
rect 26237 2397 26249 2400
rect 26283 2397 26295 2431
rect 26237 2391 26295 2397
rect 26510 2388 26516 2440
rect 26568 2428 26574 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26568 2400 27169 2428
rect 26568 2388 26574 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27982 2388 27988 2440
rect 28040 2428 28046 2440
rect 28261 2431 28319 2437
rect 28261 2428 28273 2431
rect 28040 2400 28273 2428
rect 28040 2388 28046 2400
rect 28261 2397 28273 2400
rect 28307 2397 28319 2431
rect 28261 2391 28319 2397
rect 28902 2388 28908 2440
rect 28960 2428 28966 2440
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 28960 2400 29009 2428
rect 28960 2388 28966 2400
rect 28997 2397 29009 2400
rect 29043 2397 29055 2431
rect 28997 2391 29055 2397
rect 29454 2388 29460 2440
rect 29512 2428 29518 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29512 2400 29745 2428
rect 29512 2388 29518 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30469 2431 30527 2437
rect 30469 2428 30481 2431
rect 30432 2400 30481 2428
rect 30432 2388 30438 2400
rect 30469 2397 30481 2400
rect 30515 2397 30527 2431
rect 30469 2391 30527 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30892 2400 31125 2428
rect 30892 2388 30898 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 31846 2388 31852 2440
rect 31904 2428 31910 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31904 2400 32137 2428
rect 31904 2388 31910 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32232 2428 32260 2468
rect 32398 2456 32404 2468
rect 32456 2456 32462 2508
rect 38105 2499 38163 2505
rect 38105 2496 38117 2499
rect 32600 2468 38117 2496
rect 32232 2424 32444 2428
rect 32490 2424 32496 2440
rect 32232 2400 32496 2424
rect 32125 2391 32183 2397
rect 32416 2396 32496 2400
rect 32490 2388 32496 2396
rect 32548 2388 32554 2440
rect 2593 2363 2651 2369
rect 2593 2329 2605 2363
rect 2639 2360 2651 2363
rect 3694 2360 3700 2372
rect 2639 2332 3700 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 12897 2363 12955 2369
rect 12897 2329 12909 2363
rect 12943 2360 12955 2363
rect 13446 2360 13452 2372
rect 12943 2332 13452 2360
rect 12943 2329 12955 2332
rect 12897 2323 12955 2329
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 13872 2332 15669 2360
rect 13872 2320 13878 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 16022 2320 16028 2372
rect 16080 2360 16086 2372
rect 32600 2360 32628 2468
rect 38105 2465 38117 2468
rect 38151 2465 38163 2499
rect 38105 2459 38163 2465
rect 38856 2468 50384 2496
rect 16080 2332 32628 2360
rect 32692 2400 32904 2428
rect 16080 2320 16086 2332
rect 3050 2252 3056 2304
rect 3108 2292 3114 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3108 2264 3985 2292
rect 3108 2252 3114 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 5074 2252 5080 2304
rect 5132 2292 5138 2304
rect 5169 2295 5227 2301
rect 5169 2292 5181 2295
rect 5132 2264 5181 2292
rect 5132 2252 5138 2264
rect 5169 2261 5181 2264
rect 5215 2261 5227 2295
rect 5169 2255 5227 2261
rect 5994 2252 6000 2304
rect 6052 2292 6058 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6052 2264 6561 2292
rect 6052 2252 6058 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7984 2264 8033 2292
rect 7984 2252 7990 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8996 2264 9229 2292
rect 8996 2252 9002 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 10781 2295 10839 2301
rect 10781 2261 10793 2295
rect 10827 2292 10839 2295
rect 10870 2292 10876 2304
rect 10827 2264 10876 2292
rect 10827 2261 10839 2264
rect 10781 2255 10839 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 11977 2295 12035 2301
rect 11977 2292 11989 2295
rect 11940 2264 11989 2292
rect 11940 2252 11946 2264
rect 11977 2261 11989 2264
rect 12023 2261 12035 2295
rect 11977 2255 12035 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17497 2295 17555 2301
rect 17497 2292 17509 2295
rect 17276 2264 17509 2292
rect 17276 2252 17282 2264
rect 17497 2261 17509 2264
rect 17543 2261 17555 2295
rect 19978 2292 19984 2304
rect 19939 2264 19984 2292
rect 17497 2255 17555 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 22094 2252 22100 2304
rect 22152 2292 22158 2304
rect 22373 2295 22431 2301
rect 22373 2292 22385 2295
rect 22152 2264 22385 2292
rect 22152 2252 22158 2264
rect 22373 2261 22385 2264
rect 22419 2261 22431 2295
rect 22373 2255 22431 2261
rect 24578 2252 24584 2304
rect 24636 2292 24642 2304
rect 24857 2295 24915 2301
rect 24857 2292 24869 2295
rect 24636 2264 24869 2292
rect 24636 2252 24642 2264
rect 24857 2261 24869 2264
rect 24903 2261 24915 2295
rect 24857 2255 24915 2261
rect 24946 2252 24952 2304
rect 25004 2292 25010 2304
rect 32692 2292 32720 2400
rect 32876 2360 32904 2400
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34057 2431 34115 2437
rect 34057 2428 34069 2431
rect 33836 2400 34069 2428
rect 33836 2388 33842 2400
rect 34057 2397 34069 2400
rect 34103 2397 34115 2431
rect 34057 2391 34115 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 35158 2428 35164 2440
rect 35119 2400 35164 2428
rect 34885 2391 34943 2397
rect 35158 2388 35164 2400
rect 35216 2388 35222 2440
rect 35866 2400 38148 2428
rect 35866 2360 35894 2400
rect 32876 2332 35894 2360
rect 36262 2320 36268 2372
rect 36320 2360 36326 2372
rect 36449 2363 36507 2369
rect 36449 2360 36461 2363
rect 36320 2332 36461 2360
rect 36320 2320 36326 2332
rect 36449 2329 36461 2332
rect 36495 2329 36507 2363
rect 36449 2323 36507 2329
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 37921 2363 37979 2369
rect 37921 2360 37933 2363
rect 37792 2332 37933 2360
rect 37792 2320 37798 2332
rect 37921 2329 37933 2332
rect 37967 2329 37979 2363
rect 38120 2360 38148 2400
rect 38194 2388 38200 2440
rect 38252 2428 38258 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38252 2400 38761 2428
rect 38252 2388 38258 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 38856 2360 38884 2468
rect 41138 2388 41144 2440
rect 41196 2428 41202 2440
rect 41601 2431 41659 2437
rect 41601 2428 41613 2431
rect 41196 2400 41613 2428
rect 41196 2388 41202 2400
rect 41601 2397 41613 2400
rect 41647 2397 41659 2431
rect 41601 2391 41659 2397
rect 43530 2388 43536 2440
rect 43588 2428 43594 2440
rect 43625 2431 43683 2437
rect 43625 2428 43637 2431
rect 43588 2400 43637 2428
rect 43588 2388 43594 2400
rect 43625 2397 43637 2400
rect 43671 2397 43683 2431
rect 43625 2391 43683 2397
rect 45002 2388 45008 2440
rect 45060 2428 45066 2440
rect 45097 2431 45155 2437
rect 45097 2428 45109 2431
rect 45060 2400 45109 2428
rect 45060 2388 45066 2400
rect 45097 2397 45109 2400
rect 45143 2397 45155 2431
rect 45097 2391 45155 2397
rect 45462 2388 45468 2440
rect 45520 2428 45526 2440
rect 46017 2431 46075 2437
rect 46017 2428 46029 2431
rect 45520 2400 46029 2428
rect 45520 2388 45526 2400
rect 46017 2397 46029 2400
rect 46063 2397 46075 2431
rect 46017 2391 46075 2397
rect 46474 2388 46480 2440
rect 46532 2428 46538 2440
rect 46569 2431 46627 2437
rect 46569 2428 46581 2431
rect 46532 2400 46581 2428
rect 46532 2388 46538 2400
rect 46569 2397 46581 2400
rect 46615 2397 46627 2431
rect 46569 2391 46627 2397
rect 47946 2388 47952 2440
rect 48004 2428 48010 2440
rect 48041 2431 48099 2437
rect 48041 2428 48053 2431
rect 48004 2400 48053 2428
rect 48004 2388 48010 2400
rect 48041 2397 48053 2400
rect 48087 2397 48099 2431
rect 48041 2391 48099 2397
rect 48406 2388 48412 2440
rect 48464 2428 48470 2440
rect 48961 2431 49019 2437
rect 48961 2428 48973 2431
rect 48464 2400 48973 2428
rect 48464 2388 48470 2400
rect 48961 2397 48973 2400
rect 49007 2397 49019 2431
rect 48961 2391 49019 2397
rect 49418 2388 49424 2440
rect 49476 2428 49482 2440
rect 50157 2431 50215 2437
rect 50157 2428 50169 2431
rect 49476 2400 50169 2428
rect 49476 2388 49482 2400
rect 50157 2397 50169 2400
rect 50203 2397 50215 2431
rect 50157 2391 50215 2397
rect 38120 2332 38884 2360
rect 37921 2323 37979 2329
rect 39206 2320 39212 2372
rect 39264 2360 39270 2372
rect 39945 2363 40003 2369
rect 39945 2360 39957 2363
rect 39264 2332 39957 2360
rect 39264 2320 39270 2332
rect 39945 2329 39957 2332
rect 39991 2329 40003 2363
rect 39945 2323 40003 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 40773 2363 40831 2369
rect 40773 2360 40785 2363
rect 40644 2332 40785 2360
rect 40644 2320 40650 2332
rect 40773 2329 40785 2332
rect 40819 2329 40831 2363
rect 40773 2323 40831 2329
rect 42058 2320 42064 2372
rect 42116 2360 42122 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 42116 2332 42901 2360
rect 42116 2320 42122 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 50356 2360 50384 2468
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 50985 2431 51043 2437
rect 50985 2428 50997 2431
rect 50948 2400 50997 2428
rect 50948 2388 50954 2400
rect 50985 2397 50997 2400
rect 51031 2397 51043 2431
rect 50985 2391 51043 2397
rect 51350 2388 51356 2440
rect 51408 2428 51414 2440
rect 51905 2431 51963 2437
rect 51905 2428 51917 2431
rect 51408 2400 51917 2428
rect 51408 2388 51414 2400
rect 51905 2397 51917 2400
rect 51951 2397 51963 2431
rect 51905 2391 51963 2397
rect 52362 2388 52368 2440
rect 52420 2428 52426 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52420 2400 52745 2428
rect 52420 2388 52426 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 53834 2388 53840 2440
rect 53892 2428 53898 2440
rect 53929 2431 53987 2437
rect 53929 2428 53941 2431
rect 53892 2400 53941 2428
rect 53892 2388 53898 2400
rect 53929 2397 53941 2400
rect 53975 2397 53987 2431
rect 53929 2391 53987 2397
rect 55214 2388 55220 2440
rect 55272 2428 55278 2440
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 55272 2400 55321 2428
rect 55272 2388 55278 2400
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 55309 2391 55367 2397
rect 55766 2388 55772 2440
rect 55824 2428 55830 2440
rect 56229 2431 56287 2437
rect 56229 2428 56241 2431
rect 55824 2400 56241 2428
rect 55824 2388 55830 2400
rect 56229 2397 56241 2400
rect 56275 2397 56287 2431
rect 56229 2391 56287 2397
rect 57238 2388 57244 2440
rect 57296 2428 57302 2440
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 57296 2400 58081 2428
rect 57296 2388 57302 2400
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 58069 2391 58127 2397
rect 56965 2363 57023 2369
rect 50356 2332 56180 2360
rect 42889 2323 42947 2329
rect 25004 2264 32720 2292
rect 25004 2252 25010 2264
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 36541 2295 36599 2301
rect 36541 2292 36553 2295
rect 32916 2264 36553 2292
rect 32916 2252 32922 2264
rect 36541 2261 36553 2264
rect 36587 2261 36599 2295
rect 40034 2292 40040 2304
rect 39995 2264 40040 2292
rect 36541 2255 36599 2261
rect 40034 2252 40040 2264
rect 40092 2252 40098 2304
rect 40862 2292 40868 2304
rect 40823 2264 40868 2292
rect 40862 2252 40868 2264
rect 40920 2252 40926 2304
rect 42978 2292 42984 2304
rect 42939 2264 42984 2292
rect 42978 2252 42984 2264
rect 43036 2252 43042 2304
rect 43806 2292 43812 2304
rect 43767 2264 43812 2292
rect 43806 2252 43812 2264
rect 43864 2252 43870 2304
rect 45278 2292 45284 2304
rect 45239 2264 45284 2292
rect 45278 2252 45284 2264
rect 45336 2252 45342 2304
rect 46750 2292 46756 2304
rect 46711 2264 46756 2292
rect 46750 2252 46756 2264
rect 46808 2252 46814 2304
rect 48314 2252 48320 2304
rect 48372 2292 48378 2304
rect 50341 2295 50399 2301
rect 50341 2292 50353 2295
rect 48372 2264 50353 2292
rect 48372 2252 48378 2264
rect 50341 2261 50353 2264
rect 50387 2261 50399 2295
rect 52914 2292 52920 2304
rect 52875 2264 52920 2292
rect 50341 2255 50399 2261
rect 52914 2252 52920 2264
rect 52972 2252 52978 2304
rect 54110 2292 54116 2304
rect 54071 2264 54116 2292
rect 54110 2252 54116 2264
rect 54168 2252 54174 2304
rect 55490 2292 55496 2304
rect 55451 2264 55496 2292
rect 55490 2252 55496 2264
rect 55548 2252 55554 2304
rect 56152 2292 56180 2332
rect 56965 2329 56977 2363
rect 57011 2360 57023 2363
rect 58158 2360 58164 2372
rect 57011 2332 58164 2360
rect 57011 2329 57023 2332
rect 56965 2323 57023 2329
rect 58158 2320 58164 2332
rect 58216 2320 58222 2372
rect 57057 2295 57115 2301
rect 57057 2292 57069 2295
rect 56152 2264 57069 2292
rect 57057 2261 57069 2264
rect 57103 2261 57115 2295
rect 57057 2255 57115 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 14918 2048 14924 2100
rect 14976 2088 14982 2100
rect 46750 2088 46756 2100
rect 14976 2060 46756 2088
rect 14976 2048 14982 2060
rect 46750 2048 46756 2060
rect 46808 2048 46814 2100
rect 18966 1980 18972 2032
rect 19024 2020 19030 2032
rect 48314 2020 48320 2032
rect 19024 1992 48320 2020
rect 19024 1980 19030 1992
rect 48314 1980 48320 1992
rect 48372 1980 48378 2032
rect 14642 1912 14648 1964
rect 14700 1952 14706 1964
rect 42978 1952 42984 1964
rect 14700 1924 42984 1952
rect 14700 1912 14706 1924
rect 42978 1912 42984 1924
rect 43036 1912 43042 1964
rect 15010 1844 15016 1896
rect 15068 1884 15074 1896
rect 40034 1884 40040 1896
rect 15068 1856 40040 1884
rect 15068 1844 15074 1856
rect 40034 1844 40040 1856
rect 40092 1844 40098 1896
rect 20438 1776 20444 1828
rect 20496 1816 20502 1828
rect 31018 1816 31024 1828
rect 20496 1788 31024 1816
rect 20496 1776 20502 1788
rect 31018 1776 31024 1788
rect 31076 1776 31082 1828
rect 15102 1708 15108 1760
rect 15160 1748 15166 1760
rect 40862 1748 40868 1760
rect 15160 1720 40868 1748
rect 15160 1708 15166 1720
rect 40862 1708 40868 1720
rect 40920 1708 40926 1760
rect 15838 1640 15844 1692
rect 15896 1680 15902 1692
rect 35158 1680 35164 1692
rect 15896 1652 35164 1680
rect 15896 1640 15902 1652
rect 35158 1640 35164 1652
rect 35216 1640 35222 1692
rect 20806 1572 20812 1624
rect 20864 1612 20870 1624
rect 55490 1612 55496 1624
rect 20864 1584 55496 1612
rect 20864 1572 20870 1584
rect 55490 1572 55496 1584
rect 55548 1572 55554 1624
rect 20622 1504 20628 1556
rect 20680 1544 20686 1556
rect 52914 1544 52920 1556
rect 20680 1516 52920 1544
rect 20680 1504 20686 1516
rect 52914 1504 52920 1516
rect 52972 1504 52978 1556
rect 20530 1436 20536 1488
rect 20588 1476 20594 1488
rect 54110 1476 54116 1488
rect 20588 1448 54116 1476
rect 20588 1436 20594 1448
rect 54110 1436 54116 1448
rect 54168 1436 54174 1488
<< via1 >>
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 2780 39584 2832 39636
rect 3056 39627 3108 39636
rect 3056 39593 3065 39627
rect 3065 39593 3099 39627
rect 3099 39593 3108 39627
rect 3056 39584 3108 39593
rect 3700 39584 3752 39636
rect 26240 39584 26292 39636
rect 41420 39627 41472 39636
rect 41420 39593 41429 39627
rect 41429 39593 41463 39627
rect 41463 39593 41472 39627
rect 41420 39584 41472 39593
rect 48688 39584 48740 39636
rect 56140 39584 56192 39636
rect 18696 39448 18748 39500
rect 2136 39423 2188 39432
rect 2136 39389 2145 39423
rect 2145 39389 2179 39423
rect 2179 39389 2188 39423
rect 2136 39380 2188 39389
rect 9496 39380 9548 39432
rect 6644 39312 6696 39364
rect 1584 39287 1636 39296
rect 1584 39253 1593 39287
rect 1593 39253 1627 39287
rect 1627 39253 1636 39287
rect 1584 39244 1636 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 2596 38904 2648 38956
rect 1584 38743 1636 38752
rect 1584 38709 1593 38743
rect 1593 38709 1627 38743
rect 1627 38709 1636 38743
rect 1584 38700 1636 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 2872 38496 2924 38548
rect 1492 38292 1544 38344
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 1400 37859 1452 37868
rect 1400 37825 1409 37859
rect 1409 37825 1443 37859
rect 1443 37825 1452 37859
rect 1400 37816 1452 37825
rect 1584 37655 1636 37664
rect 1584 37621 1593 37655
rect 1593 37621 1627 37655
rect 1627 37621 1636 37655
rect 1584 37612 1636 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 1768 36728 1820 36780
rect 1584 36635 1636 36644
rect 1584 36601 1593 36635
rect 1593 36601 1627 36635
rect 1627 36601 1636 36635
rect 1584 36592 1636 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1676 36116 1728 36168
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5448 35028 5500 35080
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 2872 34688 2924 34740
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2044 33940 2096 33992
rect 1584 33847 1636 33856
rect 1584 33813 1593 33847
rect 1593 33813 1627 33847
rect 1627 33813 1636 33847
rect 1584 33804 1636 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 1584 33507 1636 33516
rect 1584 33473 1593 33507
rect 1593 33473 1627 33507
rect 1627 33473 1636 33507
rect 1584 33464 1636 33473
rect 2412 33507 2464 33516
rect 2412 33473 2421 33507
rect 2421 33473 2455 33507
rect 2455 33473 2464 33507
rect 2412 33464 2464 33473
rect 4988 33328 5040 33380
rect 2228 33303 2280 33312
rect 2228 33269 2237 33303
rect 2237 33269 2271 33303
rect 2271 33269 2280 33303
rect 2228 33260 2280 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4620 32988 4672 33040
rect 4988 32963 5040 32972
rect 4988 32929 4997 32963
rect 4997 32929 5031 32963
rect 5031 32929 5040 32963
rect 4988 32920 5040 32929
rect 5080 32963 5132 32972
rect 5080 32929 5089 32963
rect 5089 32929 5123 32963
rect 5123 32929 5132 32963
rect 5080 32920 5132 32929
rect 2228 32784 2280 32836
rect 2780 32784 2832 32836
rect 4804 32716 4856 32768
rect 4896 32759 4948 32768
rect 4896 32725 4905 32759
rect 4905 32725 4939 32759
rect 4939 32725 4948 32759
rect 4896 32716 4948 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 1584 32555 1636 32564
rect 1584 32521 1593 32555
rect 1593 32521 1627 32555
rect 1627 32521 1636 32555
rect 1584 32512 1636 32521
rect 2412 32555 2464 32564
rect 2412 32521 2421 32555
rect 2421 32521 2455 32555
rect 2455 32521 2464 32555
rect 2412 32512 2464 32521
rect 2872 32555 2924 32564
rect 2872 32521 2881 32555
rect 2881 32521 2915 32555
rect 2915 32521 2924 32555
rect 2872 32512 2924 32521
rect 4896 32512 4948 32564
rect 4620 32444 4672 32496
rect 3332 32376 3384 32428
rect 4712 32419 4764 32428
rect 4712 32385 4746 32419
rect 4746 32385 4764 32419
rect 4712 32376 4764 32385
rect 3148 32308 3200 32360
rect 2780 32240 2832 32292
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4712 31968 4764 32020
rect 2964 31900 3016 31952
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 3056 31807 3108 31816
rect 3056 31773 3065 31807
rect 3065 31773 3099 31807
rect 3099 31773 3108 31807
rect 3056 31764 3108 31773
rect 4804 31764 4856 31816
rect 2872 31671 2924 31680
rect 2872 31637 2881 31671
rect 2881 31637 2915 31671
rect 2915 31637 2924 31671
rect 2872 31628 2924 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 2872 31356 2924 31408
rect 4620 31356 4672 31408
rect 3700 31288 3752 31340
rect 4896 31331 4948 31340
rect 4896 31297 4905 31331
rect 4905 31297 4939 31331
rect 4939 31297 4948 31331
rect 4896 31288 4948 31297
rect 4988 31331 5040 31340
rect 4988 31297 4997 31331
rect 4997 31297 5031 31331
rect 5031 31297 5040 31331
rect 4988 31288 5040 31297
rect 2780 31220 2832 31272
rect 1584 31195 1636 31204
rect 1584 31161 1593 31195
rect 1593 31161 1627 31195
rect 1627 31161 1636 31195
rect 1584 31152 1636 31161
rect 1400 31084 1452 31136
rect 1860 31084 1912 31136
rect 2872 31084 2924 31136
rect 4804 31084 4856 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3056 30880 3108 30932
rect 2964 30787 3016 30796
rect 2964 30753 2973 30787
rect 2973 30753 3007 30787
rect 3007 30753 3016 30787
rect 2964 30744 3016 30753
rect 3148 30787 3200 30796
rect 3148 30753 3157 30787
rect 3157 30753 3191 30787
rect 3191 30753 3200 30787
rect 3148 30744 3200 30753
rect 4712 30744 4764 30796
rect 5080 30744 5132 30796
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 2872 30719 2924 30728
rect 2872 30685 2881 30719
rect 2881 30685 2915 30719
rect 2915 30685 2924 30719
rect 2872 30676 2924 30685
rect 4620 30540 4672 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4988 30336 5040 30388
rect 7564 30268 7616 30320
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 2780 30064 2832 30116
rect 1584 30039 1636 30048
rect 1584 30005 1593 30039
rect 1593 30005 1627 30039
rect 1627 30005 1636 30039
rect 1584 29996 1636 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2688 29792 2740 29844
rect 4712 29656 4764 29708
rect 1584 29631 1636 29640
rect 1584 29597 1593 29631
rect 1593 29597 1627 29631
rect 1627 29597 1636 29631
rect 1584 29588 1636 29597
rect 4988 29588 5040 29640
rect 4620 29520 4672 29572
rect 2872 29452 2924 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 2872 29291 2924 29300
rect 2872 29257 2881 29291
rect 2881 29257 2915 29291
rect 2915 29257 2924 29291
rect 2872 29248 2924 29257
rect 2412 29112 2464 29164
rect 2780 29155 2832 29164
rect 2780 29121 2789 29155
rect 2789 29121 2823 29155
rect 2823 29121 2832 29155
rect 2780 29112 2832 29121
rect 2228 29044 2280 29096
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 2504 28908 2556 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2688 28500 2740 28552
rect 2320 28432 2372 28484
rect 2780 28364 2832 28416
rect 3792 28364 3844 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 2320 28203 2372 28212
rect 2320 28169 2329 28203
rect 2329 28169 2363 28203
rect 2363 28169 2372 28203
rect 2320 28160 2372 28169
rect 1400 28024 1452 28076
rect 2504 28067 2556 28076
rect 2504 28033 2513 28067
rect 2513 28033 2547 28067
rect 2547 28033 2556 28067
rect 2504 28024 2556 28033
rect 3884 28067 3936 28076
rect 3884 28033 3893 28067
rect 3893 28033 3927 28067
rect 3927 28033 3936 28067
rect 3884 28024 3936 28033
rect 3976 27999 4028 28008
rect 3976 27965 3985 27999
rect 3985 27965 4019 27999
rect 4019 27965 4028 27999
rect 3976 27956 4028 27965
rect 2320 27888 2372 27940
rect 2688 27820 2740 27872
rect 4068 27820 4120 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3976 27616 4028 27668
rect 2412 27455 2464 27464
rect 2412 27421 2421 27455
rect 2421 27421 2455 27455
rect 2455 27421 2464 27455
rect 2412 27412 2464 27421
rect 3056 27455 3108 27464
rect 3056 27421 3065 27455
rect 3065 27421 3099 27455
rect 3099 27421 3108 27455
rect 3056 27412 3108 27421
rect 2780 27344 2832 27396
rect 13084 27412 13136 27464
rect 3976 27344 4028 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 2228 27319 2280 27328
rect 2228 27285 2237 27319
rect 2237 27285 2271 27319
rect 2271 27285 2280 27319
rect 2228 27276 2280 27285
rect 3884 27276 3936 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 1952 27072 2004 27124
rect 3976 27115 4028 27124
rect 3976 27081 3985 27115
rect 3985 27081 4019 27115
rect 4019 27081 4028 27115
rect 3976 27072 4028 27081
rect 2228 27004 2280 27056
rect 2780 26936 2832 26988
rect 4160 26979 4212 26988
rect 4160 26945 4169 26979
rect 4169 26945 4203 26979
rect 4203 26945 4212 26979
rect 4160 26936 4212 26945
rect 3148 26775 3200 26784
rect 3148 26741 3157 26775
rect 3157 26741 3191 26775
rect 3191 26741 3200 26775
rect 3148 26732 3200 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2412 26528 2464 26580
rect 3148 26528 3200 26580
rect 2412 26392 2464 26444
rect 2688 26435 2740 26444
rect 2688 26401 2697 26435
rect 2697 26401 2731 26435
rect 2731 26401 2740 26435
rect 2688 26392 2740 26401
rect 4896 26460 4948 26512
rect 3884 26435 3936 26444
rect 3884 26401 3893 26435
rect 3893 26401 3927 26435
rect 3927 26401 3936 26435
rect 3884 26392 3936 26401
rect 15752 26392 15804 26444
rect 3792 26299 3844 26308
rect 3792 26265 3801 26299
rect 3801 26265 3835 26299
rect 3835 26265 3844 26299
rect 3792 26256 3844 26265
rect 3976 26256 4028 26308
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 3424 25848 3476 25900
rect 3608 25644 3660 25696
rect 3884 25644 3936 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4068 25440 4120 25492
rect 1952 25236 2004 25288
rect 3884 25236 3936 25288
rect 7932 25168 7984 25220
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 3424 24939 3476 24948
rect 3424 24905 3433 24939
rect 3433 24905 3467 24939
rect 3467 24905 3476 24939
rect 3424 24896 3476 24905
rect 4068 24896 4120 24948
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 2228 24760 2280 24812
rect 3608 24760 3660 24812
rect 2688 24624 2740 24676
rect 2136 24556 2188 24608
rect 2412 24556 2464 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1952 24148 2004 24200
rect 2136 24191 2188 24200
rect 2136 24157 2170 24191
rect 2170 24157 2188 24191
rect 2136 24148 2188 24157
rect 1400 24012 1452 24064
rect 1676 24012 1728 24064
rect 3792 24012 3844 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 2228 23851 2280 23860
rect 2228 23817 2237 23851
rect 2237 23817 2271 23851
rect 2271 23817 2280 23851
rect 2228 23808 2280 23817
rect 2688 23851 2740 23860
rect 2688 23817 2697 23851
rect 2697 23817 2731 23851
rect 2731 23817 2740 23851
rect 2688 23808 2740 23817
rect 3792 23740 3844 23792
rect 1676 23672 1728 23724
rect 3516 23715 3568 23724
rect 3516 23681 3525 23715
rect 3525 23681 3559 23715
rect 3559 23681 3568 23715
rect 3516 23672 3568 23681
rect 2412 23604 2464 23656
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1584 23264 1636 23316
rect 1768 23264 1820 23316
rect 1768 23128 1820 23180
rect 1952 23128 2004 23180
rect 1400 23060 1452 23112
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 5540 23060 5592 23112
rect 4620 22992 4672 23044
rect 1952 22924 2004 22976
rect 3884 22924 3936 22976
rect 3976 22924 4028 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 3884 22763 3936 22772
rect 3884 22729 3893 22763
rect 3893 22729 3927 22763
rect 3927 22729 3936 22763
rect 3884 22720 3936 22729
rect 4620 22763 4672 22772
rect 4620 22729 4629 22763
rect 4629 22729 4663 22763
rect 4663 22729 4672 22763
rect 4620 22720 4672 22729
rect 3976 22652 4028 22704
rect 2044 22584 2096 22636
rect 2412 22627 2464 22636
rect 2412 22593 2421 22627
rect 2421 22593 2455 22627
rect 2455 22593 2464 22627
rect 2412 22584 2464 22593
rect 2688 22516 2740 22568
rect 1216 22380 1268 22432
rect 2136 22380 2188 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 3240 22176 3292 22185
rect 5356 22176 5408 22228
rect 1768 22040 1820 22092
rect 3976 22083 4028 22092
rect 3976 22049 3985 22083
rect 3985 22049 4019 22083
rect 4019 22049 4028 22083
rect 3976 22040 4028 22049
rect 2136 22015 2188 22024
rect 2136 21981 2170 22015
rect 2170 21981 2188 22015
rect 2136 21972 2188 21981
rect 3792 22015 3844 22024
rect 3792 21981 3801 22015
rect 3801 21981 3835 22015
rect 3835 21981 3844 22015
rect 3792 21972 3844 21981
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 4804 22083 4856 22092
rect 4804 22049 4813 22083
rect 4813 22049 4847 22083
rect 4847 22049 4856 22083
rect 4804 22040 4856 22049
rect 5540 22040 5592 22092
rect 4896 21972 4948 22024
rect 9680 21972 9732 22024
rect 10876 21972 10928 22024
rect 2228 21836 2280 21888
rect 5264 21836 5316 21888
rect 8024 21904 8076 21956
rect 8116 21836 8168 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 1584 21632 1636 21684
rect 2136 21632 2188 21684
rect 2412 21632 2464 21684
rect 3240 21632 3292 21684
rect 8024 21675 8076 21684
rect 8024 21641 8033 21675
rect 8033 21641 8067 21675
rect 8067 21641 8076 21675
rect 8024 21632 8076 21641
rect 17316 21564 17368 21616
rect 1676 21496 1728 21548
rect 1952 21496 2004 21548
rect 7472 21496 7524 21548
rect 1400 21360 1452 21412
rect 8484 21539 8536 21548
rect 8484 21505 8493 21539
rect 8493 21505 8527 21539
rect 8527 21505 8536 21539
rect 8484 21496 8536 21505
rect 9680 21496 9732 21548
rect 10416 21496 10468 21548
rect 8576 21428 8628 21480
rect 2688 21360 2740 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 10968 21335 11020 21344
rect 10968 21301 10977 21335
rect 10977 21301 11011 21335
rect 11011 21301 11020 21335
rect 10968 21292 11020 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1768 21088 1820 21140
rect 1952 21088 2004 21140
rect 8208 21131 8260 21140
rect 8208 21097 8217 21131
rect 8217 21097 8251 21131
rect 8251 21097 8260 21131
rect 8208 21088 8260 21097
rect 10416 21131 10468 21140
rect 10416 21097 10425 21131
rect 10425 21097 10459 21131
rect 10459 21097 10468 21131
rect 10416 21088 10468 21097
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 1492 21020 1544 21072
rect 1860 21020 1912 21072
rect 7564 21020 7616 21072
rect 2136 20952 2188 21004
rect 5264 20952 5316 21004
rect 5540 20952 5592 21004
rect 8116 20995 8168 21004
rect 8116 20961 8125 20995
rect 8125 20961 8159 20995
rect 8159 20961 8168 20995
rect 8116 20952 8168 20961
rect 10968 21020 11020 21072
rect 1584 20927 1636 20936
rect 1584 20893 1593 20927
rect 1593 20893 1627 20927
rect 1627 20893 1636 20927
rect 1584 20884 1636 20893
rect 1860 20884 1912 20936
rect 2412 20927 2464 20936
rect 2412 20893 2421 20927
rect 2421 20893 2455 20927
rect 2455 20893 2464 20927
rect 2412 20884 2464 20893
rect 4712 20884 4764 20936
rect 8392 20884 8444 20936
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 1308 20816 1360 20868
rect 1768 20816 1820 20868
rect 7288 20816 7340 20868
rect 10968 20884 11020 20936
rect 11612 20816 11664 20868
rect 2044 20748 2096 20800
rect 2228 20791 2280 20800
rect 2228 20757 2237 20791
rect 2237 20757 2271 20791
rect 2271 20757 2280 20791
rect 2228 20748 2280 20757
rect 3332 20748 3384 20800
rect 8300 20748 8352 20800
rect 8576 20748 8628 20800
rect 12532 20884 12584 20936
rect 12440 20816 12492 20868
rect 14648 20859 14700 20868
rect 14648 20825 14682 20859
rect 14682 20825 14700 20859
rect 14648 20816 14700 20825
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 3332 20587 3384 20596
rect 3332 20553 3341 20587
rect 3341 20553 3375 20587
rect 3375 20553 3384 20587
rect 3332 20544 3384 20553
rect 4068 20544 4120 20596
rect 7288 20587 7340 20596
rect 7288 20553 7297 20587
rect 7297 20553 7331 20587
rect 7331 20553 7340 20587
rect 7288 20544 7340 20553
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 14648 20587 14700 20596
rect 14648 20553 14657 20587
rect 14657 20553 14691 20587
rect 14691 20553 14700 20587
rect 14648 20544 14700 20553
rect 2228 20519 2280 20528
rect 2228 20485 2262 20519
rect 2262 20485 2280 20519
rect 2228 20476 2280 20485
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 7472 20451 7524 20460
rect 7472 20417 7481 20451
rect 7481 20417 7515 20451
rect 7515 20417 7524 20451
rect 7472 20408 7524 20417
rect 7932 20408 7984 20460
rect 8392 20408 8444 20460
rect 9036 20408 9088 20460
rect 12532 20408 12584 20460
rect 12716 20408 12768 20460
rect 13452 20408 13504 20460
rect 15016 20451 15068 20460
rect 15016 20417 15025 20451
rect 15025 20417 15059 20451
rect 15059 20417 15068 20451
rect 15016 20408 15068 20417
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 8300 20383 8352 20392
rect 8300 20349 8309 20383
rect 8309 20349 8343 20383
rect 8343 20349 8352 20383
rect 8300 20340 8352 20349
rect 7380 20204 7432 20256
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2412 20000 2464 20052
rect 2688 20000 2740 20052
rect 7380 20043 7432 20052
rect 7380 20009 7389 20043
rect 7389 20009 7423 20043
rect 7423 20009 7432 20043
rect 7380 20000 7432 20009
rect 12716 20043 12768 20052
rect 1584 19975 1636 19984
rect 1584 19941 1593 19975
rect 1593 19941 1627 19975
rect 1627 19941 1636 19975
rect 1584 19932 1636 19941
rect 2504 19932 2556 19984
rect 12716 20009 12725 20043
rect 12725 20009 12759 20043
rect 12759 20009 12768 20043
rect 12716 20000 12768 20009
rect 15016 20043 15068 20052
rect 2044 19864 2096 19916
rect 12808 19932 12860 19984
rect 15016 20009 15025 20043
rect 15025 20009 15059 20043
rect 15059 20009 15068 20043
rect 15016 20000 15068 20009
rect 2412 19796 2464 19848
rect 3332 19796 3384 19848
rect 6552 19796 6604 19848
rect 8392 19864 8444 19916
rect 12348 19839 12400 19848
rect 7288 19728 7340 19780
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 13084 19796 13136 19848
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 15752 19796 15804 19848
rect 7748 19703 7800 19712
rect 7748 19669 7757 19703
rect 7757 19669 7791 19703
rect 7791 19669 7800 19703
rect 7748 19660 7800 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 3700 19456 3752 19508
rect 7288 19456 7340 19508
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 1584 19363 1636 19372
rect 1584 19329 1593 19363
rect 1593 19329 1627 19363
rect 1627 19329 1636 19363
rect 1584 19320 1636 19329
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 5448 19252 5500 19304
rect 7472 19320 7524 19372
rect 14004 19456 14056 19508
rect 12532 19388 12584 19440
rect 8208 19320 8260 19372
rect 12348 19320 12400 19372
rect 14280 19320 14332 19372
rect 14648 19320 14700 19372
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 7748 19184 7800 19236
rect 9680 19252 9732 19304
rect 12900 19295 12952 19304
rect 12900 19261 12909 19295
rect 12909 19261 12943 19295
rect 12943 19261 12952 19295
rect 12900 19252 12952 19261
rect 9772 19184 9824 19236
rect 2688 19116 2740 19168
rect 7380 19116 7432 19168
rect 8024 19116 8076 19168
rect 16856 19184 16908 19236
rect 12808 19159 12860 19168
rect 12808 19125 12817 19159
rect 12817 19125 12851 19159
rect 12851 19125 12860 19159
rect 12808 19116 12860 19125
rect 13176 19159 13228 19168
rect 13176 19125 13185 19159
rect 13185 19125 13219 19159
rect 13219 19125 13228 19159
rect 13176 19116 13228 19125
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 15568 19116 15620 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2228 18912 2280 18964
rect 5448 18955 5500 18964
rect 5448 18921 5457 18955
rect 5457 18921 5491 18955
rect 5491 18921 5500 18955
rect 5448 18912 5500 18921
rect 9036 18955 9088 18964
rect 9036 18921 9045 18955
rect 9045 18921 9079 18955
rect 9079 18921 9088 18955
rect 9036 18912 9088 18921
rect 12900 18912 12952 18964
rect 12808 18844 12860 18896
rect 14464 18912 14516 18964
rect 16856 18955 16908 18964
rect 16856 18921 16865 18955
rect 16865 18921 16899 18955
rect 16899 18921 16908 18955
rect 16856 18912 16908 18921
rect 1952 18776 2004 18828
rect 3976 18776 4028 18828
rect 7472 18776 7524 18828
rect 10968 18819 11020 18828
rect 10968 18785 10977 18819
rect 10977 18785 11011 18819
rect 11011 18785 11020 18819
rect 10968 18776 11020 18785
rect 2228 18708 2280 18760
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 7748 18751 7800 18760
rect 7748 18717 7757 18751
rect 7757 18717 7791 18751
rect 7791 18717 7800 18751
rect 7748 18708 7800 18717
rect 4160 18640 4212 18692
rect 7472 18640 7524 18692
rect 9680 18708 9732 18760
rect 12532 18708 12584 18760
rect 13176 18751 13228 18760
rect 13176 18717 13185 18751
rect 13185 18717 13219 18751
rect 13219 18717 13228 18751
rect 13176 18708 13228 18717
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 14280 18751 14332 18760
rect 13268 18708 13320 18717
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 13544 18640 13596 18692
rect 15568 18708 15620 18760
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 2136 18572 2188 18624
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2688 18368 2740 18377
rect 4160 18368 4212 18420
rect 15200 18368 15252 18420
rect 1400 18300 1452 18352
rect 14464 18300 14516 18352
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 3240 18232 3292 18284
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 7564 18232 7616 18284
rect 2504 18164 2556 18216
rect 7748 18207 7800 18216
rect 7748 18173 7757 18207
rect 7757 18173 7791 18207
rect 7791 18173 7800 18207
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 10968 18232 11020 18284
rect 7748 18164 7800 18173
rect 9772 18164 9824 18216
rect 12808 18232 12860 18284
rect 14372 18232 14424 18284
rect 13544 18207 13596 18216
rect 13544 18173 13553 18207
rect 13553 18173 13587 18207
rect 13587 18173 13596 18207
rect 13544 18164 13596 18173
rect 2688 18028 2740 18080
rect 4620 18028 4672 18080
rect 5172 18028 5224 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1768 17824 1820 17876
rect 7380 17824 7432 17876
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 7196 17688 7248 17740
rect 1952 17620 2004 17672
rect 2136 17663 2188 17672
rect 2136 17629 2170 17663
rect 2170 17629 2188 17663
rect 2136 17620 2188 17629
rect 7564 17620 7616 17672
rect 14372 17620 14424 17672
rect 14648 17620 14700 17672
rect 14188 17552 14240 17604
rect 16764 17620 16816 17672
rect 17224 17552 17276 17604
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 7656 17484 7708 17536
rect 18052 17527 18104 17536
rect 18052 17493 18061 17527
rect 18061 17493 18095 17527
rect 18095 17493 18104 17527
rect 18052 17484 18104 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 2412 17212 2464 17264
rect 18052 17212 18104 17264
rect 2320 17144 2372 17196
rect 5724 17144 5776 17196
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 9772 17187 9824 17196
rect 7380 17144 7432 17153
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 17132 17187 17184 17196
rect 17132 17153 17166 17187
rect 17166 17153 17184 17187
rect 17132 17144 17184 17153
rect 1860 17076 1912 17128
rect 11520 17076 11572 17128
rect 16764 17076 16816 17128
rect 11060 17008 11112 17060
rect 7380 16940 7432 16992
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 12348 16940 12400 16992
rect 15200 16940 15252 16992
rect 16396 16940 16448 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7380 16779 7432 16788
rect 7380 16745 7389 16779
rect 7389 16745 7423 16779
rect 7423 16745 7432 16779
rect 7380 16736 7432 16745
rect 11520 16779 11572 16788
rect 11520 16745 11529 16779
rect 11529 16745 11563 16779
rect 11563 16745 11572 16779
rect 11520 16736 11572 16745
rect 2412 16668 2464 16720
rect 2688 16668 2740 16720
rect 17132 16736 17184 16788
rect 17408 16668 17460 16720
rect 1952 16600 2004 16652
rect 2136 16532 2188 16584
rect 6644 16532 6696 16584
rect 7288 16575 7340 16584
rect 7288 16541 7297 16575
rect 7297 16541 7331 16575
rect 7331 16541 7340 16575
rect 7288 16532 7340 16541
rect 4068 16464 4120 16516
rect 5356 16464 5408 16516
rect 16396 16600 16448 16652
rect 18052 16600 18104 16652
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 10968 16532 11020 16584
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 2228 16439 2280 16448
rect 2228 16405 2237 16439
rect 2237 16405 2271 16439
rect 2271 16405 2280 16439
rect 2228 16396 2280 16405
rect 2504 16396 2556 16448
rect 7288 16396 7340 16448
rect 7840 16396 7892 16448
rect 10232 16464 10284 16516
rect 10876 16396 10928 16448
rect 12348 16532 12400 16584
rect 15200 16532 15252 16584
rect 17592 16532 17644 16584
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 17132 16464 17184 16516
rect 18604 16439 18656 16448
rect 18604 16405 18613 16439
rect 18613 16405 18647 16439
rect 18647 16405 18656 16439
rect 18604 16396 18656 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 2044 16192 2096 16244
rect 1492 16124 1544 16176
rect 1400 16056 1452 16108
rect 2228 16124 2280 16176
rect 5356 16192 5408 16244
rect 7840 16235 7892 16244
rect 7840 16201 7849 16235
rect 7849 16201 7883 16235
rect 7883 16201 7892 16235
rect 7840 16192 7892 16201
rect 17224 16235 17276 16244
rect 14556 16124 14608 16176
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 18604 16192 18656 16244
rect 6644 16099 6696 16108
rect 1952 15988 2004 16040
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 6736 16099 6788 16108
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 7656 16099 7708 16108
rect 6736 16056 6788 16065
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 8208 16056 8260 16108
rect 10232 16056 10284 16108
rect 10784 16056 10836 16108
rect 13544 16056 13596 16108
rect 15660 16099 15712 16108
rect 5816 15920 5868 15972
rect 3424 15895 3476 15904
rect 3424 15861 3433 15895
rect 3433 15861 3467 15895
rect 3467 15861 3476 15895
rect 3424 15852 3476 15861
rect 5080 15852 5132 15904
rect 7380 15920 7432 15972
rect 10968 15988 11020 16040
rect 12532 15988 12584 16040
rect 14464 15988 14516 16040
rect 14924 15988 14976 16040
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 15844 16056 15896 16108
rect 17684 16099 17736 16108
rect 17684 16065 17693 16099
rect 17693 16065 17727 16099
rect 17727 16065 17736 16099
rect 17684 16056 17736 16065
rect 17592 15988 17644 16040
rect 7012 15895 7064 15904
rect 7012 15861 7021 15895
rect 7021 15861 7055 15895
rect 7055 15861 7064 15895
rect 7012 15852 7064 15861
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11152 15852 11204 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 4068 15648 4120 15700
rect 1952 15580 2004 15632
rect 6736 15648 6788 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 10968 15648 11020 15700
rect 12532 15648 12584 15700
rect 14280 15648 14332 15700
rect 15660 15648 15712 15700
rect 17408 15691 17460 15700
rect 17408 15657 17417 15691
rect 17417 15657 17451 15691
rect 17451 15657 17460 15691
rect 17408 15648 17460 15657
rect 12440 15580 12492 15632
rect 2596 15555 2648 15564
rect 2596 15521 2605 15555
rect 2605 15521 2639 15555
rect 2639 15521 2648 15555
rect 2596 15512 2648 15521
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 5264 15555 5316 15564
rect 2688 15512 2740 15521
rect 5264 15521 5273 15555
rect 5273 15521 5307 15555
rect 5307 15521 5316 15555
rect 5264 15512 5316 15521
rect 7012 15512 7064 15564
rect 14556 15555 14608 15564
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 3424 15444 3476 15496
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 17316 15512 17368 15564
rect 8024 15444 8076 15496
rect 10876 15444 10928 15496
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 11980 15444 12032 15496
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 17132 15444 17184 15496
rect 18604 15444 18656 15496
rect 8300 15376 8352 15428
rect 1400 15351 1452 15360
rect 1400 15317 1409 15351
rect 1409 15317 1443 15351
rect 1443 15317 1452 15351
rect 1400 15308 1452 15317
rect 17868 15308 17920 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 18604 15147 18656 15156
rect 18604 15113 18613 15147
rect 18613 15113 18647 15147
rect 18647 15113 18656 15147
rect 18604 15104 18656 15113
rect 8300 15079 8352 15088
rect 8300 15045 8309 15079
rect 8309 15045 8343 15079
rect 8343 15045 8352 15079
rect 8300 15036 8352 15045
rect 2044 14968 2096 15020
rect 2320 14968 2372 15020
rect 7104 14968 7156 15020
rect 7748 14968 7800 15020
rect 10876 15036 10928 15088
rect 12164 14968 12216 15020
rect 17500 15011 17552 15020
rect 17500 14977 17534 15011
rect 17534 14977 17552 15011
rect 17500 14968 17552 14977
rect 11244 14900 11296 14952
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 14280 14900 14332 14952
rect 16764 14900 16816 14952
rect 1584 14875 1636 14884
rect 1584 14841 1593 14875
rect 1593 14841 1627 14875
rect 1627 14841 1636 14875
rect 1584 14832 1636 14841
rect 5724 14832 5776 14884
rect 10324 14832 10376 14884
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 9220 14764 9272 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 2688 14560 2740 14612
rect 10324 14603 10376 14612
rect 10324 14569 10333 14603
rect 10333 14569 10367 14603
rect 10367 14569 10376 14603
rect 10324 14560 10376 14569
rect 10508 14560 10560 14612
rect 11244 14603 11296 14612
rect 11244 14569 11253 14603
rect 11253 14569 11287 14603
rect 11287 14569 11296 14603
rect 11244 14560 11296 14569
rect 14280 14560 14332 14612
rect 17316 14560 17368 14612
rect 17500 14603 17552 14612
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 4620 14492 4672 14544
rect 1400 14424 1452 14476
rect 5816 14467 5868 14476
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 2688 14356 2740 14408
rect 5816 14433 5825 14467
rect 5825 14433 5859 14467
rect 5859 14433 5868 14467
rect 5816 14424 5868 14433
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 14924 14492 14976 14544
rect 5908 14424 5960 14433
rect 11060 14424 11112 14476
rect 8760 14356 8812 14408
rect 9220 14399 9272 14408
rect 9220 14365 9254 14399
rect 9254 14365 9272 14399
rect 9220 14356 9272 14365
rect 10876 14399 10928 14408
rect 10876 14365 10885 14399
rect 10885 14365 10919 14399
rect 10919 14365 10928 14399
rect 10876 14356 10928 14365
rect 12900 14356 12952 14408
rect 13728 14356 13780 14408
rect 14464 14356 14516 14408
rect 16856 14399 16908 14408
rect 4252 14331 4304 14340
rect 4252 14297 4261 14331
rect 4261 14297 4295 14331
rect 4295 14297 4304 14331
rect 4252 14288 4304 14297
rect 3332 14220 3384 14272
rect 7748 14288 7800 14340
rect 13636 14288 13688 14340
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 17592 14356 17644 14408
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 19340 14356 19392 14408
rect 17132 14288 17184 14340
rect 5356 14263 5408 14272
rect 5356 14229 5365 14263
rect 5365 14229 5399 14263
rect 5399 14229 5408 14263
rect 5356 14220 5408 14229
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 17224 14220 17276 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 2228 13991 2280 14000
rect 2228 13957 2262 13991
rect 2262 13957 2280 13991
rect 2228 13948 2280 13957
rect 1860 13880 1912 13932
rect 16856 14016 16908 14068
rect 3148 13880 3200 13932
rect 3516 13880 3568 13932
rect 5356 13880 5408 13932
rect 14096 13880 14148 13932
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 9772 13812 9824 13864
rect 10232 13812 10284 13864
rect 10508 13812 10560 13864
rect 11704 13812 11756 13864
rect 12532 13812 12584 13864
rect 13728 13812 13780 13864
rect 16764 13880 16816 13932
rect 16948 13923 17000 13932
rect 16948 13889 16982 13923
rect 16982 13889 17000 13923
rect 16948 13880 17000 13889
rect 3332 13787 3384 13796
rect 3332 13753 3341 13787
rect 3341 13753 3375 13787
rect 3375 13753 3384 13787
rect 3332 13744 3384 13753
rect 4252 13744 4304 13796
rect 4804 13676 4856 13728
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 7104 13676 7156 13728
rect 10784 13676 10836 13728
rect 13912 13676 13964 13728
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 5264 13336 5316 13388
rect 5632 13472 5684 13524
rect 5724 13472 5776 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 10508 13472 10560 13524
rect 14096 13515 14148 13524
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 16948 13472 17000 13524
rect 4804 13200 4856 13252
rect 5540 13268 5592 13320
rect 4344 13175 4396 13184
rect 4344 13141 4353 13175
rect 4353 13141 4387 13175
rect 4387 13141 4396 13175
rect 4344 13132 4396 13141
rect 7564 13200 7616 13252
rect 13084 13404 13136 13456
rect 9680 13336 9732 13388
rect 10048 13336 10100 13388
rect 10508 13336 10560 13388
rect 13912 13336 13964 13388
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 10876 13268 10928 13320
rect 12900 13268 12952 13320
rect 13636 13268 13688 13320
rect 13728 13268 13780 13320
rect 15568 13268 15620 13320
rect 17224 13311 17276 13320
rect 15016 13200 15068 13252
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 17500 13268 17552 13320
rect 17132 13200 17184 13252
rect 10508 13132 10560 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 5816 12928 5868 12980
rect 6276 12928 6328 12980
rect 4620 12903 4672 12912
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 4620 12869 4629 12903
rect 4629 12869 4663 12903
rect 4663 12869 4672 12903
rect 4620 12860 4672 12869
rect 6736 12928 6788 12980
rect 9496 12928 9548 12980
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 17132 12928 17184 12980
rect 7564 12860 7616 12912
rect 8760 12835 8812 12844
rect 4344 12724 4396 12776
rect 5908 12724 5960 12776
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 10140 12792 10192 12844
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 12900 12792 12952 12844
rect 7656 12724 7708 12776
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 6736 12656 6788 12708
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 4620 12588 4672 12640
rect 6368 12588 6420 12640
rect 6460 12588 6512 12640
rect 12348 12656 12400 12708
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 13728 12588 13780 12640
rect 15292 12792 15344 12844
rect 16948 12792 17000 12844
rect 16764 12724 16816 12776
rect 15476 12588 15528 12640
rect 17316 12588 17368 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2412 12384 2464 12436
rect 5632 12384 5684 12436
rect 2688 12248 2740 12300
rect 8760 12384 8812 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 12348 12384 12400 12436
rect 13636 12384 13688 12436
rect 15476 12384 15528 12436
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 4620 12180 4672 12232
rect 6368 12180 6420 12232
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 12532 12180 12584 12232
rect 12716 12180 12768 12232
rect 13360 12180 13412 12232
rect 15292 12180 15344 12232
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 13268 12112 13320 12164
rect 2596 12087 2648 12096
rect 2596 12053 2605 12087
rect 2605 12053 2639 12087
rect 2639 12053 2648 12087
rect 2596 12044 2648 12053
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 8024 12044 8076 12096
rect 12440 12044 12492 12096
rect 13728 12112 13780 12164
rect 13636 12044 13688 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2044 11840 2096 11892
rect 13268 11883 13320 11892
rect 2228 11772 2280 11824
rect 4344 11772 4396 11824
rect 10324 11772 10376 11824
rect 10876 11772 10928 11824
rect 1952 11704 2004 11756
rect 5632 11704 5684 11756
rect 7748 11704 7800 11756
rect 8208 11636 8260 11688
rect 13268 11849 13277 11883
rect 13277 11849 13311 11883
rect 13311 11849 13320 11883
rect 13268 11840 13320 11849
rect 13636 11883 13688 11892
rect 13636 11849 13645 11883
rect 13645 11849 13679 11883
rect 13679 11849 13688 11883
rect 13636 11840 13688 11849
rect 13728 11840 13780 11892
rect 14556 11772 14608 11824
rect 16304 11772 16356 11824
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 18696 11704 18748 11756
rect 15936 11636 15988 11688
rect 2596 11500 2648 11552
rect 8944 11568 8996 11620
rect 12256 11568 12308 11620
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 9588 11500 9640 11552
rect 15476 11568 15528 11620
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 17868 11500 17920 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1584 11271 1636 11280
rect 1584 11237 1593 11271
rect 1593 11237 1627 11271
rect 1627 11237 1636 11271
rect 1584 11228 1636 11237
rect 6828 11228 6880 11280
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8944 11135 8996 11144
rect 8208 11092 8260 11101
rect 8392 11067 8444 11076
rect 8392 11033 8401 11067
rect 8401 11033 8435 11067
rect 8435 11033 8444 11067
rect 8392 11024 8444 11033
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 13544 11296 13596 11348
rect 15936 11339 15988 11348
rect 15936 11305 15945 11339
rect 15945 11305 15979 11339
rect 15979 11305 15988 11339
rect 15936 11296 15988 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 12532 11228 12584 11280
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 10876 11024 10928 11076
rect 13636 11024 13688 11076
rect 16672 11092 16724 11144
rect 16764 11092 16816 11144
rect 17040 11092 17092 11144
rect 12440 10956 12492 11008
rect 15292 11024 15344 11076
rect 17592 11067 17644 11076
rect 17592 11033 17626 11067
rect 17626 11033 17644 11067
rect 17592 11024 17644 11033
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 12808 10752 12860 10804
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 15660 10795 15712 10804
rect 15660 10761 15669 10795
rect 15669 10761 15703 10795
rect 15703 10761 15712 10795
rect 15660 10752 15712 10761
rect 17592 10752 17644 10804
rect 17868 10795 17920 10804
rect 17868 10761 17877 10795
rect 17877 10761 17911 10795
rect 17911 10761 17920 10795
rect 17868 10752 17920 10761
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 3884 10616 3936 10668
rect 7932 10616 7984 10668
rect 8208 10616 8260 10668
rect 11704 10684 11756 10736
rect 12072 10616 12124 10668
rect 17132 10684 17184 10736
rect 16580 10616 16632 10668
rect 18420 10616 18472 10668
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 5816 10548 5868 10600
rect 2872 10412 2924 10464
rect 15936 10412 15988 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 5632 10140 5684 10192
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3240 10004 3292 10056
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5816 10004 5868 10056
rect 6736 10004 6788 10056
rect 8208 10004 8260 10056
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 14372 10004 14424 10056
rect 6368 9979 6420 9988
rect 6368 9945 6402 9979
rect 6402 9945 6420 9979
rect 6368 9936 6420 9945
rect 2872 9868 2924 9920
rect 8852 9868 8904 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 2872 9664 2924 9716
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 2964 9596 3016 9648
rect 1952 9460 2004 9512
rect 2412 9460 2464 9512
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 6184 9528 6236 9580
rect 10048 9571 10100 9580
rect 7840 9460 7892 9512
rect 10048 9537 10057 9571
rect 10057 9537 10091 9571
rect 10091 9537 10100 9571
rect 10048 9528 10100 9537
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 16028 9528 16080 9580
rect 10784 9460 10836 9512
rect 13084 9460 13136 9512
rect 8852 9435 8904 9444
rect 8852 9401 8861 9435
rect 8861 9401 8895 9435
rect 8895 9401 8904 9435
rect 8852 9392 8904 9401
rect 10600 9392 10652 9444
rect 11704 9392 11756 9444
rect 10968 9324 11020 9376
rect 16120 9324 16172 9376
rect 17040 9324 17092 9376
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 6000 9163 6052 9172
rect 6000 9129 6009 9163
rect 6009 9129 6043 9163
rect 6043 9129 6052 9163
rect 6000 9120 6052 9129
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 10968 9120 11020 9172
rect 16028 9120 16080 9172
rect 2964 9052 3016 9104
rect 5632 9095 5684 9104
rect 5632 9061 5641 9095
rect 5641 9061 5675 9095
rect 5675 9061 5684 9095
rect 5632 9052 5684 9061
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2780 8916 2832 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 7748 8984 7800 9036
rect 10232 8984 10284 9036
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 8668 8916 8720 8968
rect 12164 8984 12216 9036
rect 13360 8959 13412 8968
rect 8116 8848 8168 8900
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 19156 8916 19208 8968
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 20536 8916 20588 8968
rect 11520 8848 11572 8900
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 5908 8780 5960 8832
rect 8024 8780 8076 8832
rect 20352 8848 20404 8900
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 19248 8780 19300 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 2044 8576 2096 8628
rect 11060 8576 11112 8628
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 11704 8576 11756 8628
rect 5816 8508 5868 8560
rect 6920 8508 6972 8560
rect 7748 8551 7800 8560
rect 7748 8517 7757 8551
rect 7757 8517 7791 8551
rect 7791 8517 7800 8551
rect 7748 8508 7800 8517
rect 8208 8508 8260 8560
rect 12256 8508 12308 8560
rect 15568 8576 15620 8628
rect 15752 8576 15804 8628
rect 20352 8619 20404 8628
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 5908 8440 5960 8492
rect 8668 8440 8720 8492
rect 10232 8440 10284 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12532 8440 12584 8492
rect 13176 8508 13228 8560
rect 16672 8551 16724 8560
rect 16672 8517 16681 8551
rect 16681 8517 16715 8551
rect 16715 8517 16724 8551
rect 16672 8508 16724 8517
rect 20352 8585 20361 8619
rect 20361 8585 20395 8619
rect 20395 8585 20404 8619
rect 20352 8576 20404 8585
rect 18052 8508 18104 8560
rect 13636 8440 13688 8492
rect 15936 8440 15988 8492
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 10508 8372 10560 8424
rect 17684 8440 17736 8492
rect 19248 8508 19300 8560
rect 19432 8440 19484 8492
rect 20444 8440 20496 8492
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 15200 8304 15252 8356
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 14464 8279 14516 8288
rect 14464 8245 14473 8279
rect 14473 8245 14507 8279
rect 14507 8245 14516 8279
rect 14464 8236 14516 8245
rect 17868 8236 17920 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1952 8032 2004 8084
rect 7472 8032 7524 8084
rect 7748 8032 7800 8084
rect 10508 8032 10560 8084
rect 11888 8032 11940 8084
rect 13360 8032 13412 8084
rect 11244 7964 11296 8016
rect 11980 7964 12032 8016
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 3608 7896 3660 7948
rect 11060 7896 11112 7948
rect 17868 7939 17920 7948
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 13084 7828 13136 7880
rect 17868 7905 17877 7939
rect 17877 7905 17911 7939
rect 17911 7905 17920 7939
rect 17868 7896 17920 7905
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 14832 7828 14884 7880
rect 17132 7828 17184 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 20628 7828 20680 7880
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 3792 7692 3844 7744
rect 7104 7760 7156 7812
rect 8484 7760 8536 7812
rect 19248 7760 19300 7812
rect 10600 7692 10652 7744
rect 13820 7692 13872 7744
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 3056 7488 3108 7540
rect 5908 7488 5960 7540
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 7932 7488 7984 7540
rect 13820 7488 13872 7540
rect 14004 7488 14056 7540
rect 14464 7488 14516 7540
rect 19248 7488 19300 7540
rect 4712 7420 4764 7472
rect 7564 7420 7616 7472
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 3332 7352 3384 7404
rect 6000 7352 6052 7404
rect 6920 7395 6972 7404
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 2780 7284 2832 7336
rect 4804 7284 4856 7336
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 7472 7352 7524 7404
rect 7840 7352 7892 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8852 7395 8904 7404
rect 8668 7352 8720 7361
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 5448 7216 5500 7268
rect 9772 7284 9824 7336
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 13636 7395 13688 7404
rect 10784 7284 10836 7336
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 18972 7352 19024 7404
rect 17132 7327 17184 7336
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 11060 7216 11112 7268
rect 11244 7216 11296 7268
rect 6736 7148 6788 7200
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2596 6944 2648 6996
rect 4620 6944 4672 6996
rect 6000 6944 6052 6996
rect 7840 6944 7892 6996
rect 4528 6876 4580 6928
rect 4712 6876 4764 6928
rect 8208 6876 8260 6928
rect 11060 6876 11112 6928
rect 1952 6808 2004 6860
rect 8852 6808 8904 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 5448 6740 5500 6792
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 2596 6672 2648 6724
rect 3516 6672 3568 6724
rect 7288 6783 7340 6792
rect 2780 6604 2832 6656
rect 4804 6604 4856 6656
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 7472 6740 7524 6792
rect 8208 6740 8260 6792
rect 13820 6808 13872 6860
rect 14464 6808 14516 6860
rect 14740 6808 14792 6860
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10692 6740 10744 6792
rect 15936 6740 15988 6792
rect 16488 6740 16540 6792
rect 17868 6740 17920 6792
rect 10416 6672 10468 6724
rect 10508 6604 10560 6656
rect 10600 6604 10652 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 3332 6443 3384 6452
rect 3332 6409 3341 6443
rect 3341 6409 3375 6443
rect 3375 6409 3384 6443
rect 3332 6400 3384 6409
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 8208 6400 8260 6452
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 10876 6400 10928 6452
rect 11796 6400 11848 6452
rect 14648 6400 14700 6452
rect 14740 6400 14792 6452
rect 6000 6332 6052 6384
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3608 6264 3660 6316
rect 6736 6264 6788 6316
rect 10048 6264 10100 6316
rect 11336 6332 11388 6384
rect 11704 6332 11756 6384
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 14464 6264 14516 6316
rect 16396 6264 16448 6316
rect 43812 6400 43864 6452
rect 1676 6196 1728 6248
rect 7564 6196 7616 6248
rect 14556 6196 14608 6248
rect 10692 6128 10744 6180
rect 13084 6128 13136 6180
rect 16948 6128 17000 6180
rect 17040 6128 17092 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 2688 6060 2740 6112
rect 5356 6060 5408 6112
rect 13636 6060 13688 6112
rect 45284 6332 45336 6384
rect 18880 6103 18932 6112
rect 18880 6069 18889 6103
rect 18889 6069 18923 6103
rect 18923 6069 18932 6103
rect 18880 6060 18932 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 13452 5856 13504 5908
rect 15108 5856 15160 5908
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 15660 5788 15712 5840
rect 3424 5720 3476 5772
rect 3608 5720 3660 5772
rect 7564 5720 7616 5772
rect 16948 5763 17000 5772
rect 16948 5729 16957 5763
rect 16957 5729 16991 5763
rect 16991 5729 17000 5763
rect 16948 5720 17000 5729
rect 1492 5652 1544 5704
rect 6644 5652 6696 5704
rect 6828 5695 6880 5704
rect 6828 5661 6862 5695
rect 6862 5661 6880 5695
rect 6828 5652 6880 5661
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 15016 5652 15068 5704
rect 16028 5652 16080 5704
rect 17868 5652 17920 5704
rect 19064 5652 19116 5704
rect 18880 5584 18932 5636
rect 2596 5516 2648 5568
rect 3608 5516 3660 5568
rect 7288 5516 7340 5568
rect 7840 5516 7892 5568
rect 14740 5516 14792 5568
rect 17040 5516 17092 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 10692 5312 10744 5364
rect 13268 5312 13320 5364
rect 14740 5312 14792 5364
rect 15844 5312 15896 5364
rect 17592 5312 17644 5364
rect 3240 5244 3292 5296
rect 19432 5244 19484 5296
rect 2504 5219 2556 5228
rect 2504 5185 2538 5219
rect 2538 5185 2556 5219
rect 2504 5176 2556 5185
rect 3516 5176 3568 5228
rect 5448 5176 5500 5228
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 11152 5176 11204 5228
rect 14464 5176 14516 5228
rect 15108 5176 15160 5228
rect 17040 5219 17092 5228
rect 3792 5108 3844 5160
rect 5172 5108 5224 5160
rect 9956 5108 10008 5160
rect 10784 5108 10836 5160
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 18512 5176 18564 5228
rect 30288 5176 30340 5228
rect 6828 5040 6880 5092
rect 3148 4972 3200 5024
rect 5724 4972 5776 5024
rect 6736 5015 6788 5024
rect 6736 4981 6745 5015
rect 6745 4981 6779 5015
rect 6779 4981 6788 5015
rect 6736 4972 6788 4981
rect 10508 5040 10560 5092
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 11520 4972 11572 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2504 4768 2556 4820
rect 4620 4811 4672 4820
rect 4620 4777 4629 4811
rect 4629 4777 4663 4811
rect 4663 4777 4672 4811
rect 4620 4768 4672 4777
rect 6736 4768 6788 4820
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 14188 4768 14240 4820
rect 17776 4768 17828 4820
rect 3608 4632 3660 4684
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 3516 4564 3568 4616
rect 5448 4632 5500 4684
rect 4712 4564 4764 4616
rect 17040 4632 17092 4684
rect 3884 4496 3936 4548
rect 10784 4564 10836 4616
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 15844 4607 15896 4616
rect 9772 4496 9824 4548
rect 11520 4539 11572 4548
rect 11520 4505 11529 4539
rect 11529 4505 11563 4539
rect 11563 4505 11572 4539
rect 11520 4496 11572 4505
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 16488 4564 16540 4616
rect 18512 4564 18564 4616
rect 28816 4496 28868 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 8208 4428 8260 4480
rect 9956 4428 10008 4480
rect 17040 4428 17092 4480
rect 18696 4428 18748 4480
rect 19432 4428 19484 4480
rect 24676 4428 24728 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 1400 4224 1452 4276
rect 9956 4224 10008 4276
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 18512 4224 18564 4276
rect 19432 4224 19484 4276
rect 2136 4156 2188 4208
rect 3516 4156 3568 4208
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 2872 4020 2924 4072
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 4620 4088 4672 4140
rect 5264 4156 5316 4208
rect 5448 4088 5500 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5172 4020 5224 4072
rect 5356 4020 5408 4072
rect 8024 4156 8076 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 9772 4131 9824 4140
rect 6828 4088 6880 4097
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 3700 3952 3752 4004
rect 10416 4088 10468 4140
rect 16212 4088 16264 4140
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 18696 4088 18748 4140
rect 19340 4131 19392 4140
rect 11336 4020 11388 4072
rect 16488 4020 16540 4072
rect 19340 4097 19349 4131
rect 19349 4097 19383 4131
rect 19383 4097 19392 4131
rect 19340 4088 19392 4097
rect 19432 4088 19484 4140
rect 23020 4088 23072 4140
rect 26056 4020 26108 4072
rect 10968 3952 11020 4004
rect 2964 3884 3016 3936
rect 3884 3884 3936 3936
rect 3976 3884 4028 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 6460 3884 6512 3936
rect 14924 3884 14976 3936
rect 17132 3952 17184 4004
rect 33692 3952 33744 4004
rect 21272 3884 21324 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2688 3680 2740 3732
rect 10876 3680 10928 3732
rect 16580 3723 16632 3732
rect 16580 3689 16589 3723
rect 16589 3689 16623 3723
rect 16623 3689 16632 3723
rect 16580 3680 16632 3689
rect 17500 3680 17552 3732
rect 19156 3680 19208 3732
rect 23756 3680 23808 3732
rect 5172 3655 5224 3664
rect 5172 3621 5181 3655
rect 5181 3621 5215 3655
rect 5215 3621 5224 3655
rect 5172 3612 5224 3621
rect 5448 3612 5500 3664
rect 6644 3612 6696 3664
rect 3056 3544 3108 3596
rect 3516 3544 3568 3596
rect 4804 3544 4856 3596
rect 10784 3612 10836 3664
rect 9588 3544 9640 3596
rect 15568 3612 15620 3664
rect 16120 3612 16172 3664
rect 16488 3544 16540 3596
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3884 3476 3936 3528
rect 6460 3519 6512 3528
rect 204 3340 256 3392
rect 1676 3340 1728 3392
rect 2780 3340 2832 3392
rect 3240 3408 3292 3460
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 6552 3476 6604 3528
rect 7472 3476 7524 3528
rect 10324 3476 10376 3528
rect 10968 3476 11020 3528
rect 3608 3340 3660 3392
rect 3700 3340 3752 3392
rect 7840 3408 7892 3460
rect 11336 3476 11388 3528
rect 13360 3476 13412 3528
rect 14740 3476 14792 3528
rect 15292 3476 15344 3528
rect 23664 3544 23716 3596
rect 6276 3383 6328 3392
rect 6276 3349 6285 3383
rect 6285 3349 6319 3383
rect 6319 3349 6328 3383
rect 6276 3340 6328 3349
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 12716 3408 12768 3460
rect 17684 3476 17736 3528
rect 16856 3408 16908 3460
rect 17960 3408 18012 3460
rect 18604 3476 18656 3528
rect 18788 3476 18840 3528
rect 21088 3476 21140 3528
rect 22468 3408 22520 3460
rect 59636 3408 59688 3460
rect 10784 3340 10836 3392
rect 12440 3340 12492 3392
rect 12992 3340 13044 3392
rect 16948 3383 17000 3392
rect 16948 3349 16957 3383
rect 16957 3349 16991 3383
rect 16991 3349 17000 3383
rect 16948 3340 17000 3349
rect 18052 3340 18104 3392
rect 18696 3340 18748 3392
rect 19248 3383 19300 3392
rect 19248 3349 19257 3383
rect 19257 3349 19291 3383
rect 19291 3349 19300 3383
rect 19248 3340 19300 3349
rect 21180 3383 21232 3392
rect 21180 3349 21189 3383
rect 21189 3349 21223 3383
rect 21223 3349 21232 3383
rect 21180 3340 21232 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 3608 3136 3660 3188
rect 4896 3136 4948 3188
rect 8024 3136 8076 3188
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11612 3136 11664 3188
rect 12440 3136 12492 3188
rect 13452 3136 13504 3188
rect 14372 3136 14424 3188
rect 1952 3000 2004 3052
rect 3976 3068 4028 3120
rect 4068 3068 4120 3120
rect 5632 3068 5684 3120
rect 6276 3068 6328 3120
rect 7564 3068 7616 3120
rect 16948 3136 17000 3188
rect 4160 3000 4212 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6644 3000 6696 3052
rect 8208 3000 8260 3052
rect 9312 3000 9364 3052
rect 10876 3043 10928 3052
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 2596 2932 2648 2984
rect 8024 2932 8076 2984
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 3608 2864 3660 2916
rect 9036 2864 9088 2916
rect 10968 2932 11020 2984
rect 12716 2932 12768 2984
rect 16304 3068 16356 3120
rect 14740 3000 14792 3052
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15936 3000 15988 3052
rect 16856 3000 16908 3052
rect 19248 3136 19300 3188
rect 23664 3179 23716 3188
rect 23664 3145 23673 3179
rect 23673 3145 23707 3179
rect 23707 3145 23716 3179
rect 23664 3136 23716 3145
rect 23756 3136 23808 3188
rect 17408 3068 17460 3120
rect 18052 3111 18104 3120
rect 18052 3077 18061 3111
rect 18061 3077 18095 3111
rect 18095 3077 18104 3111
rect 18052 3068 18104 3077
rect 17960 3000 18012 3052
rect 21180 3068 21232 3120
rect 23020 3068 23072 3120
rect 32404 3068 32456 3120
rect 21272 3043 21324 3052
rect 13452 2932 13504 2941
rect 15568 2932 15620 2984
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 23572 3000 23624 3052
rect 27436 3000 27488 3052
rect 33692 3043 33744 3052
rect 33692 3009 33701 3043
rect 33701 3009 33735 3043
rect 33735 3009 33744 3043
rect 33692 3000 33744 3009
rect 56692 3000 56744 3052
rect 22468 2932 22520 2984
rect 17316 2864 17368 2916
rect 19616 2864 19668 2916
rect 22192 2864 22244 2916
rect 33324 2932 33376 2984
rect 664 2796 716 2848
rect 3792 2796 3844 2848
rect 6368 2796 6420 2848
rect 8484 2796 8536 2848
rect 11796 2796 11848 2848
rect 12348 2796 12400 2848
rect 19156 2796 19208 2848
rect 21640 2796 21692 2848
rect 32312 2796 32364 2848
rect 35348 2796 35400 2848
rect 36728 2796 36780 2848
rect 39672 2796 39724 2848
rect 42616 2796 42668 2848
rect 44088 2796 44140 2848
rect 46940 2796 46992 2848
rect 49884 2796 49936 2848
rect 52828 2796 52880 2848
rect 54300 2796 54352 2848
rect 58716 2796 58768 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2872 2592 2924 2644
rect 4712 2592 4764 2644
rect 12532 2635 12584 2644
rect 12532 2601 12541 2635
rect 12541 2601 12575 2635
rect 12575 2601 12584 2635
rect 12532 2592 12584 2601
rect 15476 2592 15528 2644
rect 19800 2592 19852 2644
rect 1124 2456 1176 2508
rect 5540 2456 5592 2508
rect 8392 2456 8444 2508
rect 14280 2524 14332 2576
rect 17776 2524 17828 2576
rect 24952 2592 25004 2644
rect 26056 2635 26108 2644
rect 26056 2601 26065 2635
rect 26065 2601 26099 2635
rect 26099 2601 26108 2635
rect 26056 2592 26108 2601
rect 28816 2635 28868 2644
rect 28816 2601 28825 2635
rect 28825 2601 28859 2635
rect 28859 2601 28868 2635
rect 28816 2592 28868 2601
rect 30288 2635 30340 2644
rect 30288 2601 30297 2635
rect 30297 2601 30331 2635
rect 30331 2601 30340 2635
rect 30288 2592 30340 2601
rect 31024 2592 31076 2644
rect 20076 2524 20128 2576
rect 1308 2388 1360 2440
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 9404 2388 9456 2440
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 16764 2456 16816 2508
rect 19064 2456 19116 2508
rect 32404 2499 32456 2508
rect 17316 2431 17368 2440
rect 17316 2397 17325 2431
rect 17325 2397 17359 2431
rect 17359 2397 17368 2431
rect 17316 2388 17368 2397
rect 19616 2388 19668 2440
rect 20168 2388 20220 2440
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 22560 2388 22612 2440
rect 24032 2388 24084 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 25044 2388 25096 2440
rect 25964 2388 26016 2440
rect 26516 2388 26568 2440
rect 27988 2388 28040 2440
rect 28908 2388 28960 2440
rect 29460 2388 29512 2440
rect 30380 2388 30432 2440
rect 30840 2388 30892 2440
rect 31852 2388 31904 2440
rect 32404 2465 32413 2499
rect 32413 2465 32447 2499
rect 32447 2465 32456 2499
rect 32404 2456 32456 2465
rect 32496 2388 32548 2440
rect 3700 2320 3752 2372
rect 13452 2320 13504 2372
rect 13820 2320 13872 2372
rect 16028 2320 16080 2372
rect 3056 2252 3108 2304
rect 5080 2252 5132 2304
rect 6000 2252 6052 2304
rect 7932 2252 7984 2304
rect 8944 2252 8996 2304
rect 10876 2252 10928 2304
rect 11888 2252 11940 2304
rect 14832 2252 14884 2304
rect 17224 2252 17276 2304
rect 19984 2295 20036 2304
rect 19984 2261 19993 2295
rect 19993 2261 20027 2295
rect 20027 2261 20036 2295
rect 19984 2252 20036 2261
rect 22100 2252 22152 2304
rect 24584 2252 24636 2304
rect 24952 2252 25004 2304
rect 33784 2388 33836 2440
rect 34796 2388 34848 2440
rect 35164 2431 35216 2440
rect 35164 2397 35173 2431
rect 35173 2397 35207 2431
rect 35207 2397 35216 2431
rect 35164 2388 35216 2397
rect 36268 2320 36320 2372
rect 37740 2320 37792 2372
rect 38200 2388 38252 2440
rect 41144 2388 41196 2440
rect 43536 2388 43588 2440
rect 45008 2388 45060 2440
rect 45468 2388 45520 2440
rect 46480 2388 46532 2440
rect 47952 2388 48004 2440
rect 48412 2388 48464 2440
rect 49424 2388 49476 2440
rect 39212 2320 39264 2372
rect 40592 2320 40644 2372
rect 42064 2320 42116 2372
rect 50896 2388 50948 2440
rect 51356 2388 51408 2440
rect 52368 2388 52420 2440
rect 53840 2388 53892 2440
rect 55220 2388 55272 2440
rect 55772 2388 55824 2440
rect 57244 2388 57296 2440
rect 32864 2252 32916 2304
rect 40040 2295 40092 2304
rect 40040 2261 40049 2295
rect 40049 2261 40083 2295
rect 40083 2261 40092 2295
rect 40040 2252 40092 2261
rect 40868 2295 40920 2304
rect 40868 2261 40877 2295
rect 40877 2261 40911 2295
rect 40911 2261 40920 2295
rect 40868 2252 40920 2261
rect 42984 2295 43036 2304
rect 42984 2261 42993 2295
rect 42993 2261 43027 2295
rect 43027 2261 43036 2295
rect 42984 2252 43036 2261
rect 43812 2295 43864 2304
rect 43812 2261 43821 2295
rect 43821 2261 43855 2295
rect 43855 2261 43864 2295
rect 43812 2252 43864 2261
rect 45284 2295 45336 2304
rect 45284 2261 45293 2295
rect 45293 2261 45327 2295
rect 45327 2261 45336 2295
rect 45284 2252 45336 2261
rect 46756 2295 46808 2304
rect 46756 2261 46765 2295
rect 46765 2261 46799 2295
rect 46799 2261 46808 2295
rect 46756 2252 46808 2261
rect 48320 2252 48372 2304
rect 52920 2295 52972 2304
rect 52920 2261 52929 2295
rect 52929 2261 52963 2295
rect 52963 2261 52972 2295
rect 52920 2252 52972 2261
rect 54116 2295 54168 2304
rect 54116 2261 54125 2295
rect 54125 2261 54159 2295
rect 54159 2261 54168 2295
rect 54116 2252 54168 2261
rect 55496 2295 55548 2304
rect 55496 2261 55505 2295
rect 55505 2261 55539 2295
rect 55539 2261 55548 2295
rect 55496 2252 55548 2261
rect 58164 2320 58216 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 14924 2048 14976 2100
rect 46756 2048 46808 2100
rect 18972 1980 19024 2032
rect 48320 1980 48372 2032
rect 14648 1912 14700 1964
rect 42984 1912 43036 1964
rect 15016 1844 15068 1896
rect 40040 1844 40092 1896
rect 20444 1776 20496 1828
rect 31024 1776 31076 1828
rect 15108 1708 15160 1760
rect 40868 1708 40920 1760
rect 15844 1640 15896 1692
rect 35164 1640 35216 1692
rect 20812 1572 20864 1624
rect 55496 1572 55548 1624
rect 20628 1504 20680 1556
rect 52920 1504 52972 1556
rect 20536 1436 20588 1488
rect 54116 1436 54168 1488
<< metal2 >>
rect 2870 41712 2926 41721
rect 2870 41647 2926 41656
rect 2778 40080 2834 40089
rect 2778 40015 2834 40024
rect 2792 39642 2820 40015
rect 2780 39636 2832 39642
rect 2780 39578 2832 39584
rect 2136 39432 2188 39438
rect 2136 39374 2188 39380
rect 1584 39296 1636 39302
rect 1582 39264 1584 39273
rect 1636 39264 1638 39273
rect 1582 39199 1638 39208
rect 1584 38752 1636 38758
rect 1584 38694 1636 38700
rect 1596 38457 1624 38694
rect 1582 38448 1638 38457
rect 1582 38383 1638 38392
rect 1492 38344 1544 38350
rect 1492 38286 1544 38292
rect 1400 37868 1452 37874
rect 1400 37810 1452 37816
rect 1412 31142 1440 37810
rect 1400 31136 1452 31142
rect 1400 31078 1452 31084
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 26625 1440 28018
rect 1398 26616 1454 26625
rect 1398 26551 1454 26560
rect 1400 24064 1452 24070
rect 1400 24006 1452 24012
rect 1412 23202 1440 24006
rect 1320 23174 1440 23202
rect 1216 22432 1268 22438
rect 1214 22400 1216 22409
rect 1268 22400 1270 22409
rect 1214 22335 1270 22344
rect 1320 20874 1348 23174
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 21593 1440 23054
rect 1398 21584 1454 21593
rect 1398 21519 1454 21528
rect 1504 21434 1532 38286
rect 1584 37664 1636 37670
rect 1582 37632 1584 37641
rect 1636 37632 1638 37641
rect 1582 37567 1638 37576
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1582 36680 1638 36689
rect 1582 36615 1584 36624
rect 1636 36615 1638 36624
rect 1584 36586 1636 36592
rect 1676 36168 1728 36174
rect 1676 36110 1728 36116
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1596 35873 1624 35974
rect 1582 35864 1638 35873
rect 1582 35799 1638 35808
rect 1582 35048 1638 35057
rect 1582 34983 1638 34992
rect 1596 34950 1624 34983
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 34241 1624 34546
rect 1582 34232 1638 34241
rect 1582 34167 1638 34176
rect 1584 33856 1636 33862
rect 1582 33824 1584 33833
rect 1636 33824 1638 33833
rect 1582 33759 1638 33768
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1596 33017 1624 33458
rect 1582 33008 1638 33017
rect 1582 32943 1638 32952
rect 1584 32564 1636 32570
rect 1584 32506 1636 32512
rect 1596 32473 1624 32506
rect 1582 32464 1638 32473
rect 1582 32399 1638 32408
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1596 31657 1624 31758
rect 1582 31648 1638 31657
rect 1582 31583 1638 31592
rect 1582 31240 1638 31249
rect 1582 31175 1584 31184
rect 1636 31175 1638 31184
rect 1584 31146 1636 31152
rect 1584 30728 1636 30734
rect 1584 30670 1636 30676
rect 1596 30433 1624 30670
rect 1582 30424 1638 30433
rect 1582 30359 1638 30368
rect 1584 30048 1636 30054
rect 1582 30016 1584 30025
rect 1636 30016 1638 30025
rect 1582 29951 1638 29960
rect 1584 29640 1636 29646
rect 1584 29582 1636 29588
rect 1596 29209 1624 29582
rect 1582 29200 1638 29209
rect 1582 29135 1638 29144
rect 1584 29028 1636 29034
rect 1584 28970 1636 28976
rect 1596 28801 1624 28970
rect 1582 28792 1638 28801
rect 1582 28727 1638 28736
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 1596 27334 1624 27367
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1584 26240 1636 26246
rect 1582 26208 1584 26217
rect 1636 26208 1638 26217
rect 1582 26143 1638 26152
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1596 25401 1624 25842
rect 1582 25392 1638 25401
rect 1582 25327 1638 25336
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 24993 1624 25094
rect 1582 24984 1638 24993
rect 1582 24919 1638 24928
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1596 24177 1624 24754
rect 1582 24168 1638 24177
rect 1582 24103 1638 24112
rect 1688 24070 1716 36110
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1596 23769 1624 23802
rect 1582 23760 1638 23769
rect 1582 23695 1638 23704
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1596 21690 1624 23258
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1688 21554 1716 23666
rect 1780 23322 1808 36722
rect 2044 33992 2096 33998
rect 2044 33934 2096 33940
rect 1860 31136 1912 31142
rect 1860 31078 1912 31084
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1768 23180 1820 23186
rect 1768 23122 1820 23128
rect 1780 22098 1808 23122
rect 1768 22092 1820 22098
rect 1768 22034 1820 22040
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1400 21412 1452 21418
rect 1504 21406 1716 21434
rect 1400 21354 1452 21360
rect 1308 20868 1360 20874
rect 1308 20810 1360 20816
rect 1412 18358 1440 21354
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21185 1624 21286
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1492 21072 1544 21078
rect 1492 21014 1544 21020
rect 1400 18352 1452 18358
rect 1400 18294 1452 18300
rect 1398 16552 1454 16561
rect 1398 16487 1454 16496
rect 1412 16114 1440 16487
rect 1504 16182 1532 21014
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1596 20369 1624 20878
rect 1582 20360 1638 20369
rect 1582 20295 1638 20304
rect 1584 19984 1636 19990
rect 1582 19952 1584 19961
rect 1636 19952 1638 19961
rect 1582 19887 1638 19896
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1596 19145 1624 19314
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1584 18624 1636 18630
rect 1582 18592 1584 18601
rect 1636 18592 1638 18601
rect 1582 18527 1638 18536
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17785 1624 18226
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 1582 17368 1638 17377
rect 1582 17303 1584 17312
rect 1636 17303 1638 17312
rect 1584 17274 1636 17280
rect 1688 16574 1716 21406
rect 1780 21146 1808 22034
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1872 21078 1900 31078
rect 1952 27124 2004 27130
rect 1952 27066 2004 27072
rect 1964 25294 1992 27066
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 1964 24206 1992 25230
rect 1952 24200 2004 24206
rect 1952 24142 2004 24148
rect 1964 23186 1992 24142
rect 2056 24018 2084 33934
rect 2148 24970 2176 39374
rect 2596 38956 2648 38962
rect 2596 38898 2648 38904
rect 2412 33516 2464 33522
rect 2412 33458 2464 33464
rect 2228 33312 2280 33318
rect 2228 33254 2280 33260
rect 2240 32842 2268 33254
rect 2228 32836 2280 32842
rect 2228 32778 2280 32784
rect 2424 32570 2452 33458
rect 2412 32564 2464 32570
rect 2412 32506 2464 32512
rect 2412 29164 2464 29170
rect 2412 29106 2464 29112
rect 2228 29096 2280 29102
rect 2228 29038 2280 29044
rect 2240 28098 2268 29038
rect 2320 28484 2372 28490
rect 2320 28426 2372 28432
rect 2332 28218 2360 28426
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 2240 28070 2360 28098
rect 2332 27946 2360 28070
rect 2320 27940 2372 27946
rect 2320 27882 2372 27888
rect 2228 27328 2280 27334
rect 2228 27270 2280 27276
rect 2240 27062 2268 27270
rect 2228 27056 2280 27062
rect 2228 26998 2280 27004
rect 2332 26466 2360 27882
rect 2424 27690 2452 29106
rect 2504 28960 2556 28966
rect 2504 28902 2556 28908
rect 2516 28082 2544 28902
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2424 27662 2544 27690
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 2424 26586 2452 27406
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2332 26450 2452 26466
rect 2332 26444 2464 26450
rect 2332 26438 2412 26444
rect 2412 26386 2464 26392
rect 2148 24942 2360 24970
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 2148 24206 2176 24550
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2056 23990 2176 24018
rect 1952 23180 2004 23186
rect 1952 23122 2004 23128
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1964 21554 1992 22918
rect 2148 22658 2176 23990
rect 2240 23866 2268 24754
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22817 2268 23054
rect 2226 22808 2282 22817
rect 2226 22743 2282 22752
rect 2044 22636 2096 22642
rect 2148 22630 2268 22658
rect 2044 22578 2096 22584
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 1952 21140 2004 21146
rect 1952 21082 2004 21088
rect 1860 21072 1912 21078
rect 1860 21014 1912 21020
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1768 20868 1820 20874
rect 1768 20810 1820 20816
rect 1780 17882 1808 20810
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1872 17134 1900 20878
rect 1964 20466 1992 21082
rect 2056 20890 2084 22578
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 2148 22030 2176 22374
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 2240 21894 2268 22630
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2148 21010 2176 21626
rect 2136 21004 2188 21010
rect 2136 20946 2188 20952
rect 2056 20862 2176 20890
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 2056 19922 2084 20742
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2148 19334 2176 20862
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2240 20534 2268 20742
rect 2228 20528 2280 20534
rect 2228 20470 2280 20476
rect 2226 20360 2282 20369
rect 2226 20295 2282 20304
rect 2056 19306 2176 19334
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 17678 1992 18770
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1964 16658 1992 17614
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1688 16546 1900 16574
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1492 16176 1544 16182
rect 1596 16153 1624 16390
rect 1492 16118 1544 16124
rect 1582 16144 1638 16153
rect 1400 16108 1452 16114
rect 1582 16079 1638 16088
rect 1400 16050 1452 16056
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1400 15360 1452 15366
rect 1596 15337 1624 15438
rect 1400 15302 1452 15308
rect 1582 15328 1638 15337
rect 1412 14482 1440 15302
rect 1582 15263 1638 15272
rect 1582 14920 1638 14929
rect 1582 14855 1584 14864
rect 1636 14855 1638 14864
rect 1584 14826 1636 14832
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13977 1624 14350
rect 1582 13968 1638 13977
rect 1872 13938 1900 16546
rect 1964 16046 1992 16594
rect 2056 16250 2084 19306
rect 2240 18970 2268 20295
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2148 17678 2176 18566
rect 2240 18426 2268 18702
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2332 17202 2360 24942
rect 2424 24614 2452 26386
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 23662 2452 24550
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2424 21690 2452 22578
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2412 20936 2464 20942
rect 2412 20878 2464 20884
rect 2424 20058 2452 20878
rect 2516 20369 2544 27662
rect 2502 20360 2558 20369
rect 2502 20295 2558 20304
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2424 17270 2452 19790
rect 2516 18222 2544 19926
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2412 17264 2464 17270
rect 2412 17206 2464 17212
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2516 17082 2544 18158
rect 2424 17054 2544 17082
rect 2424 16726 2452 17054
rect 2608 16980 2636 38898
rect 2884 38554 2912 41647
rect 3698 41200 3754 42000
rect 11150 41200 11206 42000
rect 18694 41200 18750 42000
rect 26146 41200 26202 42000
rect 33690 41200 33746 42000
rect 41142 41200 41198 42000
rect 48686 41200 48742 42000
rect 56138 41200 56194 42000
rect 3054 40896 3110 40905
rect 3054 40831 3110 40840
rect 3068 39642 3096 40831
rect 3712 39642 3740 41200
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 3056 39636 3108 39642
rect 3056 39578 3108 39584
rect 3700 39636 3752 39642
rect 3700 39578 3752 39584
rect 18708 39506 18736 41200
rect 26160 39658 26188 41200
rect 41156 39930 41184 41200
rect 41156 39902 41460 39930
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 26160 39642 26280 39658
rect 41432 39642 41460 39902
rect 48700 39642 48728 41200
rect 56152 39642 56180 41200
rect 26160 39636 26292 39642
rect 26160 39630 26240 39636
rect 26240 39578 26292 39584
rect 41420 39636 41472 39642
rect 41420 39578 41472 39584
rect 48688 39636 48740 39642
rect 48688 39578 48740 39584
rect 56140 39636 56192 39642
rect 56140 39578 56192 39584
rect 18696 39500 18748 39506
rect 18696 39442 18748 39448
rect 9496 39432 9548 39438
rect 9496 39374 9548 39380
rect 6644 39364 6696 39370
rect 6644 39306 6696 39312
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 2872 38548 2924 38554
rect 2872 38490 2924 38496
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 6656 35894 6684 39306
rect 6656 35866 6776 35894
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 5448 35080 5500 35086
rect 5448 35022 5500 35028
rect 2872 34740 2924 34746
rect 2872 34682 2924 34688
rect 2780 32836 2832 32842
rect 2780 32778 2832 32784
rect 2792 32298 2820 32778
rect 2884 32570 2912 34682
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4988 33380 5040 33386
rect 4988 33322 5040 33328
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4620 33040 4672 33046
rect 4620 32982 4672 32988
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 4632 32502 4660 32982
rect 5000 32978 5028 33322
rect 4988 32972 5040 32978
rect 4988 32914 5040 32920
rect 5080 32972 5132 32978
rect 5080 32914 5132 32920
rect 4804 32768 4856 32774
rect 4804 32710 4856 32716
rect 4896 32768 4948 32774
rect 4896 32710 4948 32716
rect 4620 32496 4672 32502
rect 4620 32438 4672 32444
rect 3332 32428 3384 32434
rect 3332 32370 3384 32376
rect 3148 32360 3200 32366
rect 3148 32302 3200 32308
rect 2780 32292 2832 32298
rect 2780 32234 2832 32240
rect 2792 31278 2820 32234
rect 2964 31952 3016 31958
rect 2964 31894 3016 31900
rect 2872 31680 2924 31686
rect 2872 31622 2924 31628
rect 2884 31414 2912 31622
rect 2872 31408 2924 31414
rect 2872 31350 2924 31356
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2700 29850 2728 30194
rect 2792 30122 2820 31214
rect 2872 31136 2924 31142
rect 2872 31078 2924 31084
rect 2884 30734 2912 31078
rect 2976 30802 3004 31894
rect 3056 31816 3108 31822
rect 3056 31758 3108 31764
rect 3068 30938 3096 31758
rect 3056 30932 3108 30938
rect 3056 30874 3108 30880
rect 3160 30802 3188 32302
rect 2964 30796 3016 30802
rect 2964 30738 3016 30744
rect 3148 30796 3200 30802
rect 3148 30738 3200 30744
rect 2872 30728 2924 30734
rect 2872 30670 2924 30676
rect 2780 30116 2832 30122
rect 2780 30058 2832 30064
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 2792 29322 2820 30058
rect 2872 29504 2924 29510
rect 2872 29446 2924 29452
rect 2700 29294 2820 29322
rect 2884 29306 2912 29446
rect 2872 29300 2924 29306
rect 2700 28558 2728 29294
rect 2872 29242 2924 29248
rect 2780 29164 2832 29170
rect 2780 29106 2832 29112
rect 2688 28552 2740 28558
rect 2688 28494 2740 28500
rect 2700 27962 2728 28494
rect 2792 28422 2820 29106
rect 2780 28416 2832 28422
rect 2780 28358 2832 28364
rect 2700 27934 2820 27962
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2700 26450 2728 27814
rect 2792 27402 2820 27934
rect 3054 27840 3110 27849
rect 3054 27775 3110 27784
rect 3068 27470 3096 27775
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 2780 27396 2832 27402
rect 2780 27338 2832 27344
rect 2792 26994 2820 27338
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 3160 26586 3188 26726
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 2688 26444 2740 26450
rect 2688 26386 2740 26392
rect 2688 24676 2740 24682
rect 2688 24618 2740 24624
rect 2700 23866 2728 24618
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2700 21418 2728 22510
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3252 21690 3280 22170
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 2688 21412 2740 21418
rect 2688 21354 2740 21360
rect 2700 20058 2728 21354
rect 3344 20806 3372 32370
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4632 31414 4660 32438
rect 4712 32428 4764 32434
rect 4712 32370 4764 32376
rect 4724 32026 4752 32370
rect 4712 32020 4764 32026
rect 4712 31962 4764 31968
rect 4816 31822 4844 32710
rect 4908 32570 4936 32710
rect 4896 32564 4948 32570
rect 4896 32506 4948 32512
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 4620 31408 4672 31414
rect 4620 31350 4672 31356
rect 4908 31346 4936 32506
rect 3700 31340 3752 31346
rect 3700 31282 3752 31288
rect 4896 31340 4948 31346
rect 4896 31282 4948 31288
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 3424 25900 3476 25906
rect 3424 25842 3476 25848
rect 3436 24954 3464 25842
rect 3608 25696 3660 25702
rect 3608 25638 3660 25644
rect 3424 24948 3476 24954
rect 3424 24890 3476 24896
rect 3620 24818 3648 25638
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 3344 19854 3372 20538
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18426 2728 19110
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 3528 18290 3556 23666
rect 3712 19514 3740 31282
rect 4804 31136 4856 31142
rect 4804 31078 4856 31084
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4712 30796 4764 30802
rect 4712 30738 4764 30744
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4632 29578 4660 30534
rect 4724 29714 4752 30738
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 4620 29572 4672 29578
rect 4620 29514 4672 29520
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 3792 28416 3844 28422
rect 3792 28358 3844 28364
rect 3804 26314 3832 28358
rect 3884 28076 3936 28082
rect 3884 28018 3936 28024
rect 3896 27334 3924 28018
rect 3976 28008 4028 28014
rect 3976 27950 4028 27956
rect 3988 27674 4016 27950
rect 4068 27872 4120 27878
rect 4068 27814 4120 27820
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 4080 27554 4108 27814
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4080 27526 4200 27554
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 3896 26450 3924 27270
rect 3988 27130 4016 27338
rect 3976 27124 4028 27130
rect 3976 27066 4028 27072
rect 4172 26994 4200 27526
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 3884 26444 3936 26450
rect 3884 26386 3936 26392
rect 3988 26314 4108 26330
rect 3792 26308 3844 26314
rect 3792 26250 3844 26256
rect 3976 26308 4108 26314
rect 4028 26302 4108 26308
rect 3976 26250 4028 26256
rect 3884 25696 3936 25702
rect 3884 25638 3936 25644
rect 3896 25294 3924 25638
rect 4080 25498 4108 26302
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 3884 25288 3936 25294
rect 3884 25230 3936 25236
rect 4080 24954 4108 25434
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 3792 24064 3844 24070
rect 3792 24006 3844 24012
rect 3804 23798 3832 24006
rect 3792 23792 3844 23798
rect 3792 23734 3844 23740
rect 3804 22030 3832 23734
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3896 22778 3924 22918
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3988 22710 4016 22918
rect 4632 22778 4660 22986
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 3976 22704 4028 22710
rect 3976 22646 4028 22652
rect 3988 22098 4016 22646
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3976 22092 4028 22098
rect 4724 22094 4752 29650
rect 4816 22098 4844 31078
rect 5000 30394 5028 31282
rect 5092 30802 5120 32914
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 4988 30388 5040 30394
rect 4988 30330 5040 30336
rect 5000 29646 5028 30330
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 4896 26512 4948 26518
rect 4896 26454 4948 26460
rect 3976 22034 4028 22040
rect 4632 22066 4752 22094
rect 4804 22092 4856 22098
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 20602 4108 21966
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18834 4016 19246
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4172 18426 4200 18634
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2516 16952 2636 16980
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 15638 1992 15982
rect 2148 15706 2176 16526
rect 2516 16454 2544 16952
rect 2700 16810 2728 18022
rect 3252 17542 3280 18226
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 2608 16782 2728 16810
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2240 16182 2268 16390
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1952 15632 2004 15638
rect 1952 15574 2004 15580
rect 1582 13903 1638 13912
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1964 13870 1992 15574
rect 2608 15570 2636 16782
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2700 15570 2728 16662
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1582 13560 1638 13569
rect 1582 13495 1584 13504
rect 1636 13495 1638 13504
rect 1584 13466 1636 13472
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11529 1624 12174
rect 1964 11762 1992 13806
rect 2056 11898 2084 14962
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2240 14006 2268 14758
rect 2332 14618 2360 14962
rect 2700 14618 2728 15506
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2240 11830 2268 12582
rect 2424 12442 2452 12786
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2700 12306 2728 14350
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3068 12753 3096 12786
rect 3054 12744 3110 12753
rect 3054 12679 3110 12688
rect 3160 12434 3188 13874
rect 3068 12406 3188 12434
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1582 11520 1638 11529
rect 1582 11455 1638 11464
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1596 11121 1624 11222
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10305 1624 10610
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1412 9897 1440 9998
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1688 9625 1716 9998
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1964 9518 1992 11698
rect 2608 11558 2636 12038
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 10062 2912 10406
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9722 2912 9862
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2964 9648 3016 9654
rect 2962 9616 2964 9625
rect 3016 9616 3018 9625
rect 2962 9551 3018 9560
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8537 1624 8910
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8634 2084 8774
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1582 8528 1638 8537
rect 2424 8498 2452 9454
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 1582 8463 1638 8472
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 1964 8090 1992 8434
rect 2424 8378 2452 8434
rect 2424 8350 2728 8378
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2700 7970 2728 8350
rect 2792 8129 2820 8910
rect 2778 8120 2834 8129
rect 2778 8055 2834 8064
rect 2700 7942 2820 7970
rect 2976 7954 3004 9046
rect 3068 8974 3096 12406
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 9178 3188 10542
rect 3252 10062 3280 17478
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3436 15502 3464 15846
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 13802 3372 14214
rect 3528 13938 3556 18226
rect 4632 18086 4660 22066
rect 4804 22034 4856 22040
rect 4908 22030 4936 26454
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5276 21010 5304 21830
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 4712 20936 4764 20942
rect 4712 20878 4764 20884
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4080 15706 4108 16458
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 4264 13802 4292 14282
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4356 12782 4384 13126
rect 4632 12918 4660 14486
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4632 12238 4660 12582
rect 4724 12434 4752 20878
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13258 4844 13670
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4724 12406 4936 12434
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11830 4384 12038
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3896 9382 3924 10610
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 1584 7744 1636 7750
rect 1582 7712 1584 7721
rect 1636 7712 1638 7721
rect 1582 7647 1638 7656
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1490 6896 1546 6905
rect 1964 6866 1992 7278
rect 1490 6831 1546 6840
rect 1952 6860 2004 6866
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6497 1440 6734
rect 1398 6488 1454 6497
rect 1398 6423 1454 6432
rect 1504 5710 1532 6831
rect 1952 6802 2004 6808
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6254 1716 6734
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1584 6112 1636 6118
rect 1582 6080 1584 6089
rect 1636 6080 1638 6089
rect 1582 6015 1638 6024
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1412 4282 1440 4558
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4321 1624 4422
rect 1582 4312 1638 4321
rect 1400 4276 1452 4282
rect 1582 4247 1638 4256
rect 1400 4218 1452 4224
rect 204 3392 256 3398
rect 204 3334 256 3340
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 216 800 244 3334
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 676 800 704 2790
rect 1124 2508 1176 2514
rect 1124 2450 1176 2456
rect 1136 800 1164 2450
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1320 649 1348 2382
rect 1412 1873 1440 2926
rect 1398 1864 1454 1873
rect 1398 1799 1454 1808
rect 1688 1714 1716 3334
rect 1964 3058 1992 6802
rect 2516 6746 2544 7346
rect 2608 7002 2636 7346
rect 2792 7342 2820 7942
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 3068 7546 3096 8910
rect 3160 7954 3188 9114
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2516 6730 2636 6746
rect 2516 6724 2648 6730
rect 2516 6718 2596 6724
rect 2596 6666 2648 6672
rect 2608 5930 2636 6666
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 6474 2820 6598
rect 2700 6446 2820 6474
rect 3344 6458 3372 7346
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3332 6452 3384 6458
rect 2700 6322 2728 6446
rect 3332 6394 3384 6400
rect 3528 6322 3556 6666
rect 3620 6322 3648 7890
rect 3804 7750 3832 8230
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 2700 6118 2728 6258
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2608 5902 2728 5930
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2516 4826 2544 5170
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2608 4622 2636 5510
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2136 4208 2188 4214
rect 2136 4150 2188 4156
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1596 1686 1716 1714
rect 1596 800 1624 1686
rect 2148 800 2176 4150
rect 2700 3738 2728 5902
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2884 3534 2912 4014
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2608 800 2636 2926
rect 2792 2281 2820 3334
rect 2870 2680 2926 2689
rect 2870 2615 2872 2624
rect 2924 2615 2926 2624
rect 2872 2586 2924 2592
rect 2778 2272 2834 2281
rect 2778 2207 2834 2216
rect 1306 640 1362 649
rect 1306 575 1362 584
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 2976 241 3004 3878
rect 3068 3602 3096 4422
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 800 3096 2246
rect 3160 1465 3188 4966
rect 3252 4622 3280 5238
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3436 4146 3464 5714
rect 3528 5658 3556 6258
rect 3620 5778 3648 6258
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3528 5630 3740 5658
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3620 5370 3648 5510
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3528 4729 3556 5170
rect 3514 4720 3570 4729
rect 3620 4690 3648 5306
rect 3514 4655 3570 4664
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3528 4214 3556 4558
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3528 3602 3556 4150
rect 3712 4146 3740 5630
rect 3804 5166 3832 7686
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3896 4554 3924 9318
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4540 6798 4568 6870
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4632 4826 4660 6938
rect 4724 6934 4752 7414
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4816 6662 4844 7278
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 4172 4026 4200 4422
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 4080 3998 4200 4026
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3146 1456 3202 1465
rect 3146 1391 3202 1400
rect 3252 1057 3280 3402
rect 3528 3074 3556 3538
rect 3712 3398 3740 3946
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3896 3534 3924 3878
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3620 3194 3648 3334
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3988 3126 4016 3878
rect 4080 3720 4108 3998
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4080 3692 4200 3720
rect 3976 3120 4028 3126
rect 3528 3046 3740 3074
rect 4068 3120 4120 3126
rect 3976 3062 4028 3068
rect 4066 3088 4068 3097
rect 4120 3088 4122 3097
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3238 1048 3294 1057
rect 3238 983 3294 992
rect 3620 800 3648 2858
rect 3712 2378 3740 3046
rect 4172 3058 4200 3692
rect 4066 3023 4122 3032
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3804 2446 3832 2790
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 4632 2122 4660 4082
rect 4724 2650 4752 4558
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 3602 4844 3878
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4908 3194 4936 12406
rect 5092 10146 5120 15846
rect 5184 12434 5212 18022
rect 5368 17252 5396 22170
rect 5460 19310 5488 35022
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5552 22098 5580 23054
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5552 21010 5580 22034
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6564 19378 6592 19790
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5460 18970 5488 19246
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5368 17224 5488 17252
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5368 16250 5396 16458
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5276 13394 5304 15506
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 13938 5396 14214
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5184 12406 5304 12434
rect 5092 10118 5212 10146
rect 5184 10062 5212 10118
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 5166 5212 9998
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5276 4214 5304 12406
rect 5460 10266 5488 17224
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5736 14890 5764 17138
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6656 16114 6684 16526
rect 6748 16114 6776 35866
rect 7564 30320 7616 30326
rect 7564 30262 7616 30268
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7300 20602 7328 20810
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 7484 20466 7512 21490
rect 7576 21078 7604 30262
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7564 21072 7616 21078
rect 7564 21014 7616 21020
rect 7944 20618 7972 25162
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 8036 21690 8064 21898
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 8128 21010 8156 21830
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 7944 20590 8064 20618
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7392 20058 7420 20198
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7300 19514 7328 19722
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7392 19174 7420 19994
rect 7484 19378 7512 20402
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7760 19514 7788 19654
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7484 18834 7512 19314
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7760 18766 7788 19178
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5828 14482 5856 15914
rect 6748 15706 6776 16050
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 7024 15570 7052 15846
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5552 13326 5580 13670
rect 5736 13530 5764 14214
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5644 12442 5672 13466
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5644 11762 5672 12378
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5828 11558 5856 12922
rect 5920 12782 5948 14418
rect 7116 13734 7144 14962
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6288 12832 6316 12922
rect 6288 12804 6500 12832
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6472 12646 6500 12804
rect 6748 12714 6776 12922
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6380 12238 6408 12582
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 10606 5856 11494
rect 6840 11286 6868 13466
rect 7116 12434 7144 13670
rect 7208 12594 7236 17682
rect 7392 17202 7420 17818
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7300 16590 7328 17138
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16794 7420 16934
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7300 16454 7328 16526
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7392 15978 7420 16730
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7484 12730 7512 18634
rect 7576 18290 7604 18702
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7576 17678 7604 18226
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 17338 7696 17478
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7668 15502 7696 16050
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7760 15026 7788 18158
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 16250 7880 16390
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7576 12918 7604 13194
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 7656 12776 7708 12782
rect 7484 12702 7604 12730
rect 7656 12718 7708 12724
rect 7208 12566 7512 12594
rect 7116 12406 7236 12434
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5644 9110 5672 10134
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5828 8566 5856 9998
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9722 6408 9930
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6196 9178 6224 9522
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5920 8498 5948 8774
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5920 7546 5948 8434
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6012 7410 6040 9114
rect 6748 7886 6776 9998
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 6798 5488 7210
rect 6012 7002 6040 7346
rect 6748 7206 6776 7822
rect 6932 7410 6960 8502
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7116 7546 7144 7754
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 5368 4078 5396 6054
rect 5460 5234 5488 6734
rect 6012 6390 6040 6734
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 6748 6322 6776 7142
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 5794 6776 6258
rect 6656 5766 6776 5794
rect 6656 5710 6684 5766
rect 6840 5710 6868 6598
rect 7208 6458 7236 12406
rect 7484 8090 7512 12566
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7576 7478 7604 12702
rect 7668 12102 7696 12718
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7760 11762 7788 14282
rect 7944 12434 7972 20402
rect 8036 19174 8064 20590
rect 8220 20262 8248 21082
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8312 20398 8340 20742
rect 8404 20466 8432 20878
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 19378 8248 20198
rect 8404 19922 8432 20402
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7852 12406 7972 12434
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7852 10146 7880 12406
rect 8036 12186 8064 15438
rect 8220 12434 8248 16050
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8312 15094 8340 15370
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 7944 12158 8064 12186
rect 8128 12406 8248 12434
rect 7944 11098 7972 12158
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11218 8064 12038
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7944 11070 8064 11098
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7944 10266 7972 10610
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7852 10118 7972 10146
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7760 8566 7788 8978
rect 7852 8974 7880 9454
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7760 8090 7788 8502
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7852 7410 7880 8910
rect 7944 7546 7972 10118
rect 8036 8838 8064 11070
rect 8128 8906 8156 12406
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11150 8248 11630
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8220 10674 8248 11086
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8220 8566 8248 9998
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7484 6798 7512 7346
rect 7852 7002 7880 7346
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 8220 6934 8248 8502
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 4690 5488 5170
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5184 3670 5212 4014
rect 5460 3670 5488 4082
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5644 3126 5672 4082
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5736 3058 5764 4966
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3534 6500 3878
rect 6656 3670 6684 5646
rect 7300 5574 7328 6734
rect 8220 6458 8248 6734
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7576 5778 7604 6190
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4826 6776 4966
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6840 4146 6868 5034
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 3126 6316 3334
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4540 2094 4660 2122
rect 4540 800 4568 2094
rect 5092 800 5120 2246
rect 5552 800 5580 2450
rect 6380 2446 6408 2790
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6012 800 6040 2246
rect 6564 1850 6592 3470
rect 6656 3058 6684 3606
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6472 1822 6592 1850
rect 6472 800 6500 1822
rect 7484 800 7512 3470
rect 7852 3466 7880 5510
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 3126 7604 3334
rect 8036 3194 8064 4150
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 8036 2990 8064 3130
rect 8220 3058 8248 4422
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8404 2514 8432 11018
rect 8496 7818 8524 21490
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8588 20806 8616 21422
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 9048 18970 9076 20402
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9232 14414 9260 14758
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8772 12850 8800 14350
rect 9508 13326 9536 39374
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 9692 21554 9720 21966
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10428 21146 10456 21490
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10600 20936 10652 20942
rect 10888 20924 10916 21966
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10980 21078 11008 21286
rect 13096 21146 13124 27406
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 15764 21146 15792 26386
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 10968 21072 11020 21078
rect 10968 21014 11020 21020
rect 10968 20936 11020 20942
rect 10888 20896 10968 20924
rect 10600 20878 10652 20884
rect 10968 20878 11020 20884
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9692 18766 9720 19246
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 16590 9720 18702
rect 9784 18222 9812 19178
rect 10612 18290 10640 20878
rect 10980 18834 11008 20878
rect 11612 20868 11664 20874
rect 12440 20868 12492 20874
rect 11664 20828 11836 20856
rect 11612 20810 11664 20816
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10980 18290 11008 18770
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9784 17202 9812 18158
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 13394 9720 16526
rect 9784 13870 9812 17138
rect 10244 16522 10272 17138
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10244 16114 10272 16458
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10336 15910 10364 16934
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10796 15706 10824 16050
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10888 15502 10916 16390
rect 10980 16046 11008 16526
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15706 11008 15982
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10888 15094 10916 15438
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 10336 14618 10364 14826
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10520 13870 10548 14554
rect 11072 14482 11100 17002
rect 11532 16794 11560 17070
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15502 11192 15846
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11256 14618 11284 14894
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12986 9536 13262
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8772 12442 8800 12786
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 11150 8984 11562
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8864 9450 8892 9862
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8680 8498 8708 8910
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8680 7410 8708 8434
rect 8864 7410 8892 9386
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8864 6866 8892 7346
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 9324 3058 9352 11018
rect 9600 3602 9628 11494
rect 10060 9586 10088 13330
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10152 12442 10180 12786
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10244 9042 10272 13806
rect 10520 13530 10548 13806
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10520 13394 10548 13466
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10520 12238 10548 13126
rect 10796 12850 10824 13670
rect 10888 13326 10916 14350
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10336 11830 10364 12174
rect 10888 11830 10916 12582
rect 11716 12238 11744 13806
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10612 9042 10640 9386
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10244 8498 10272 8978
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 8090 10548 8366
rect 10612 8242 10640 8978
rect 10612 8214 10732 8242
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9784 5234 9812 7278
rect 10520 7206 10548 8026
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7410 10640 7686
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6322 10088 6734
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6458 10456 6666
rect 10520 6662 10548 7142
rect 10612 6662 10640 7346
rect 10704 6798 10732 8214
rect 10796 7886 10824 9454
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7342 10824 7822
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10888 7290 10916 11018
rect 11716 10742 11744 12174
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11716 9450 11744 10678
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9178 11008 9318
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10980 7886 11008 9114
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 8634 11560 8842
rect 11716 8634 11744 9386
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11072 7954 11100 8570
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10888 7262 11008 7290
rect 11256 7274 11284 7958
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9784 4146 9812 4490
rect 9968 4486 9996 5102
rect 10520 5098 10548 6598
rect 10704 6338 10732 6734
rect 10888 6458 10916 7142
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10704 6310 10824 6338
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 5370 10732 6122
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10704 5234 10732 5306
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10796 5166 10824 6310
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9968 4282 9996 4422
rect 10152 4282 10180 4966
rect 10796 4622 10824 5102
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7944 800 7972 2246
rect 8496 800 8524 2790
rect 9048 2446 9076 2858
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 800 8984 2246
rect 9416 800 9444 2382
rect 10336 1850 10364 3470
rect 10428 3194 10456 4082
rect 10888 3738 10916 6258
rect 10980 4010 11008 7262
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11072 6934 11100 7210
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 11716 6390 11744 8434
rect 11808 6458 11836 20828
rect 12440 20810 12492 20816
rect 12452 20602 12480 20810
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12544 20466 12572 20878
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12360 19378 12388 19790
rect 12544 19446 12572 20402
rect 12728 20058 12756 20402
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12544 18766 12572 19382
rect 12820 19174 12848 19926
rect 13096 19854 13124 21082
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14660 20602 14688 20810
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18902 12848 19110
rect 12912 18970 12940 19246
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12820 18290 12848 18838
rect 13188 18766 13216 19110
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12360 16590 12388 16934
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12544 15706 12572 15982
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11900 8090 11928 8434
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11992 8022 12020 15438
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 10266 12112 10610
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12176 9042 12204 14962
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 12360 12442 12388 12650
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12452 12102 12480 15574
rect 12544 13870 12572 15642
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12912 13326 12940 14350
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 12850 12940 13262
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12532 12232 12584 12238
rect 12716 12232 12768 12238
rect 12532 12174 12584 12180
rect 12636 12180 12716 12186
rect 12636 12174 12768 12180
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12268 10062 12296 11562
rect 12544 11286 12572 12174
rect 12636 12158 12756 12174
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12636 11150 12664 12158
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12268 8566 12296 9998
rect 12452 9926 12480 10950
rect 12820 10810 12848 11086
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 13096 9518 13124 13398
rect 13280 12434 13308 18702
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13188 12406 13308 12434
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 4826 11192 5170
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11348 4622 11376 6326
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11348 4078 11376 4558
rect 11532 4554 11560 4966
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10784 3664 10836 3670
rect 10836 3612 10916 3618
rect 10784 3606 10916 3612
rect 10796 3590 10916 3606
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 3194 10824 3334
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10888 3058 10916 3590
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10980 2990 11008 3470
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10336 1822 10456 1850
rect 10428 800 10456 1822
rect 10888 800 10916 2246
rect 11348 800 11376 3470
rect 11624 3194 11652 4558
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 3194 12480 3334
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 11808 2446 11836 2790
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 800 11928 2246
rect 12360 800 12388 2790
rect 12544 2650 12572 8434
rect 13096 7886 13124 9454
rect 13188 8922 13216 12406
rect 13372 12238 13400 12718
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13280 11898 13308 12106
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13360 8968 13412 8974
rect 13188 8894 13308 8922
rect 13360 8910 13412 8916
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8566 13216 8774
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13096 6186 13124 7822
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13280 5370 13308 8894
rect 13372 8090 13400 8910
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 5914 13492 20402
rect 15028 20058 15056 20402
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13544 18692 13596 18698
rect 13544 18634 13596 18640
rect 13556 18222 13584 18634
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13556 16114 13584 18158
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 13682 13676 14282
rect 13740 13870 13768 14350
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13924 13734 13952 14894
rect 13912 13728 13964 13734
rect 13648 13654 13768 13682
rect 13912 13670 13964 13676
rect 13740 13326 13768 13654
rect 13924 13394 13952 13670
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13648 12442 13676 13262
rect 13740 12646 13768 13262
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13636 12436 13688 12442
rect 13556 12396 13636 12424
rect 13556 11354 13584 12396
rect 13636 12378 13688 12384
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11898 13676 12038
rect 13740 11898 13768 12106
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13648 8498 13676 11018
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7546 13860 7686
rect 14016 7546 14044 19450
rect 14660 19378 14688 19790
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14292 18766 14320 19314
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18970 14504 19110
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14476 18358 14504 18702
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 17882 14412 18226
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14660 17678 14688 18566
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14108 13530 14136 13874
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13648 6118 13676 7346
rect 13832 6866 13860 7482
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 14200 4826 14228 17546
rect 14384 16574 14412 17614
rect 14384 16546 14504 16574
rect 14476 16046 14504 16546
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14292 14958 14320 15642
rect 14568 15570 14596 16118
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14618 14320 14894
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14476 14414 14504 15438
rect 14936 14550 14964 15982
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13258 15056 13670
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14568 11830 14596 12922
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7410 14320 7822
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12728 2990 12756 3402
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12728 2446 12756 2926
rect 13004 2446 13032 3334
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13372 800 13400 3470
rect 14384 3194 14412 9998
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 7750 14504 8230
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 7546 14504 7686
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14476 6866 14504 7346
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14476 5710 14504 6258
rect 14568 6254 14596 7346
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14752 6458 14780 6802
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14476 5234 14504 5646
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 13464 2990 13492 3130
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13464 2378 13492 2926
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13832 800 13860 2314
rect 14292 800 14320 2518
rect 14660 1970 14688 6394
rect 14752 5574 14780 6394
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14752 5370 14780 5510
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3058 14780 3470
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14844 2774 14872 7822
rect 15120 5914 15148 20402
rect 15764 19854 15792 21082
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18766 15608 19110
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15212 16998 15240 18362
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15212 8362 15240 16526
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15672 15706 15700 16050
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15304 12238 15332 12786
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12442 15516 12582
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 11762 15332 12174
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15488 11626 15516 12378
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15304 10810 15332 11018
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15580 8634 15608 13262
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15672 10810 15700 11494
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15764 9738 15792 19314
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16868 18970 16896 19178
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17134 16804 17614
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 16658 16436 16934
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15672 9710 15792 9738
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14936 3058 14964 3878
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14844 2746 14964 2774
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 14844 800 14872 2246
rect 14936 2106 14964 2746
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 15028 1902 15056 5646
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15016 1896 15068 1902
rect 15016 1838 15068 1844
rect 15120 1766 15148 5170
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15108 1760 15160 1766
rect 15108 1702 15160 1708
rect 15304 800 15332 3470
rect 15488 2650 15516 7346
rect 15672 5846 15700 9710
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 8634 15792 9522
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15856 5370 15884 16050
rect 16776 14958 16804 17070
rect 17144 16794 17172 17138
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 17144 15502 17172 16458
rect 17236 16250 17264 17546
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17328 15570 17356 21558
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18064 17270 18092 17478
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17420 15706 17448 16662
rect 18064 16658 18092 17206
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17604 16046 17632 16526
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16776 13938 16804 14894
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16868 14074 16896 14350
rect 17144 14346 17172 15438
rect 17420 14634 17448 15642
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17328 14618 17448 14634
rect 17512 14618 17540 14962
rect 17316 14612 17448 14618
rect 17368 14606 17448 14612
rect 17500 14612 17552 14618
rect 17316 14554 17368 14560
rect 17500 14554 17552 14560
rect 17604 14414 17632 15982
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16776 12782 16804 13874
rect 16960 13530 16988 13874
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17236 13326 17264 14214
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17144 12986 17172 13194
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 11354 15976 11630
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 9058 15976 10406
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16040 9178 16068 9522
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15948 9030 16068 9058
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15948 6798 15976 8434
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16040 6610 16068 9030
rect 16132 8974 16160 9318
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15948 6582 16068 6610
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15580 2990 15608 3606
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15856 1698 15884 4558
rect 15948 3058 15976 6582
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 16040 2378 16068 5646
rect 16132 3670 16160 8434
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 15844 1692 15896 1698
rect 15844 1634 15896 1640
rect 16224 800 16252 4082
rect 16316 3126 16344 11766
rect 16776 11150 16804 12718
rect 16960 12442 16988 12786
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17144 12238 17172 12922
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 12238 17356 12582
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16408 5914 16436 6258
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16500 4622 16528 6734
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16500 4078 16528 4558
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16500 3602 16528 4014
rect 16592 3738 16620 10610
rect 16684 8566 16712 11086
rect 17052 9382 17080 11086
rect 17144 10742 17172 12174
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 17052 6186 17080 9318
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7342 17172 7822
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17144 6866 17172 7278
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 16960 5778 16988 6122
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 5234 17080 5510
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17052 4690 17080 5170
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 17052 4486 17080 4626
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17144 4010 17172 5170
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16868 3058 16896 3402
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 3194 16988 3334
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17420 3126 17448 12174
rect 17512 3738 17540 13262
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17604 10810 17632 11018
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17696 8650 17724 16050
rect 17604 8622 17724 8650
rect 17604 5370 17632 8622
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17696 4706 17724 8434
rect 17788 4826 17816 16526
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 16250 18644 16390
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 14414 17908 15302
rect 18616 15162 18644 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 10810 17908 11494
rect 18708 11354 18736 11698
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8294 17908 8910
rect 18064 8838 18092 9318
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8566 18092 8774
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 7954 17908 8230
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17880 5710 17908 6734
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17696 4678 17816 4706
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 16776 800 16804 2450
rect 17328 2446 17356 2858
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17236 800 17264 2246
rect 17696 800 17724 3470
rect 17788 2582 17816 4678
rect 18432 4146 18460 10610
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5642 18920 6054
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18524 4622 18552 5170
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4282 18552 4558
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18708 4146 18736 4422
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18616 3534 18644 4082
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17972 3058 18000 3402
rect 18708 3398 18736 4082
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18064 3126 18092 3334
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 18800 1816 18828 3470
rect 18984 2038 19012 7346
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 19076 2514 19104 5646
rect 19168 3738 19196 8910
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19260 8566 19288 8774
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19260 7818 19288 8502
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19260 7546 19288 7754
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19352 4146 19380 14350
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 19444 8498 19472 8910
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 20364 8634 20392 8842
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 19444 7886 19472 8434
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19444 4486 19472 5238
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19444 4146 19472 4218
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19260 3194 19288 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 18972 2032 19024 2038
rect 18972 1974 19024 1980
rect 18708 1788 18828 1816
rect 18708 800 18736 1788
rect 19168 800 19196 2790
rect 19628 2446 19656 2858
rect 19812 2650 20116 2666
rect 19800 2644 20116 2650
rect 19852 2638 20116 2644
rect 19800 2586 19852 2592
rect 20088 2582 20116 2638
rect 20076 2576 20128 2582
rect 20076 2518 20128 2524
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19720 870 19840 898
rect 19720 800 19748 870
rect 2962 232 3018 241
rect 2962 167 3018 176
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 19812 762 19840 870
rect 19996 762 20024 2246
rect 20180 800 20208 2382
rect 20456 1834 20484 8434
rect 20444 1828 20496 1834
rect 20444 1770 20496 1776
rect 20548 1494 20576 8910
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 1562 20668 7822
rect 20824 1630 20852 8434
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 43812 6452 43864 6458
rect 43812 6394 43864 6400
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 28816 4548 28868 4554
rect 28816 4490 28868 4496
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 21272 3936 21324 3942
rect 21272 3878 21324 3884
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20812 1624 20864 1630
rect 20812 1566 20864 1572
rect 20628 1556 20680 1562
rect 20628 1498 20680 1504
rect 20536 1488 20588 1494
rect 20536 1430 20588 1436
rect 21100 800 21128 3470
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21192 3126 21220 3334
rect 21180 3120 21232 3126
rect 21180 3062 21232 3068
rect 21284 3058 21312 3878
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 22480 2990 22508 3402
rect 23032 3126 23060 4082
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23664 3596 23716 3602
rect 23664 3538 23716 3544
rect 23676 3194 23704 3538
rect 23768 3194 23796 3674
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21652 800 21680 2790
rect 22204 2446 22232 2858
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 22112 800 22140 2246
rect 22572 800 22600 2382
rect 23584 800 23612 2994
rect 24688 2446 24716 4422
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 26068 2650 26096 4014
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 26056 2644 26108 2650
rect 26056 2586 26108 2592
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 24044 800 24072 2382
rect 24964 2310 24992 2586
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 24596 800 24624 2246
rect 25056 800 25084 2382
rect 25976 800 26004 2382
rect 26528 800 26556 2382
rect 27448 800 27476 2994
rect 28828 2650 28856 4490
rect 30300 2650 30328 5170
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 33692 4004 33744 4010
rect 33692 3946 33744 3952
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 27988 2440 28040 2446
rect 27988 2382 28040 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 28000 800 28028 2382
rect 28920 800 28948 2382
rect 29472 800 29500 2382
rect 30392 800 30420 2382
rect 30852 800 30880 2382
rect 31036 1834 31064 2586
rect 31852 2440 31904 2446
rect 31852 2382 31904 2388
rect 31024 1828 31076 1834
rect 31024 1770 31076 1776
rect 31864 800 31892 2382
rect 32324 800 32352 2790
rect 32416 2514 32444 3062
rect 33704 3058 33732 3946
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 33324 2984 33376 2990
rect 33324 2926 33376 2932
rect 32404 2508 32456 2514
rect 32404 2450 32456 2456
rect 32496 2440 32548 2446
rect 32548 2400 32904 2428
rect 32496 2382 32548 2388
rect 32876 2310 32904 2400
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 33336 800 33364 2926
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 39672 2848 39724 2854
rect 39672 2790 39724 2796
rect 42616 2848 42668 2854
rect 42616 2790 42668 2796
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 33796 800 33824 2382
rect 34808 800 34836 2382
rect 35176 1698 35204 2382
rect 35164 1692 35216 1698
rect 35164 1634 35216 1640
rect 35360 1442 35388 2790
rect 36268 2372 36320 2378
rect 36268 2314 36320 2320
rect 35268 1414 35388 1442
rect 35268 800 35296 1414
rect 36280 800 36308 2314
rect 36740 800 36768 2790
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37752 800 37780 2314
rect 38212 800 38240 2382
rect 39212 2372 39264 2378
rect 39212 2314 39264 2320
rect 39224 800 39252 2314
rect 39684 800 39712 2790
rect 41144 2440 41196 2446
rect 41144 2382 41196 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40040 2304 40092 2310
rect 40040 2246 40092 2252
rect 40052 1902 40080 2246
rect 40040 1896 40092 1902
rect 40040 1838 40092 1844
rect 40604 800 40632 2314
rect 40868 2304 40920 2310
rect 40868 2246 40920 2252
rect 40880 1766 40908 2246
rect 40868 1760 40920 1766
rect 40868 1702 40920 1708
rect 41156 800 41184 2382
rect 42064 2372 42116 2378
rect 42064 2314 42116 2320
rect 42076 800 42104 2314
rect 42628 800 42656 2790
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 42984 2304 43036 2310
rect 42984 2246 43036 2252
rect 42996 1970 43024 2246
rect 42984 1964 43036 1970
rect 42984 1906 43036 1912
rect 43548 800 43576 2382
rect 43824 2310 43852 6394
rect 45284 6384 45336 6390
rect 45284 6326 45336 6332
rect 44088 2848 44140 2854
rect 44088 2790 44140 2796
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 44100 800 44128 2790
rect 45008 2440 45060 2446
rect 45008 2382 45060 2388
rect 45020 800 45048 2382
rect 45296 2310 45324 6326
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 59636 3460 59688 3466
rect 59636 3402 59688 3408
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 56692 3052 56744 3058
rect 56692 2994 56744 3000
rect 46940 2848 46992 2854
rect 46940 2790 46992 2796
rect 49884 2848 49936 2854
rect 49884 2790 49936 2796
rect 52828 2848 52880 2854
rect 52828 2790 52880 2796
rect 54300 2848 54352 2854
rect 54300 2790 54352 2796
rect 45468 2440 45520 2446
rect 45468 2382 45520 2388
rect 46480 2440 46532 2446
rect 46480 2382 46532 2388
rect 45284 2304 45336 2310
rect 45284 2246 45336 2252
rect 45480 800 45508 2382
rect 46492 800 46520 2382
rect 46756 2304 46808 2310
rect 46756 2246 46808 2252
rect 46768 2106 46796 2246
rect 46756 2100 46808 2106
rect 46756 2042 46808 2048
rect 46952 800 46980 2790
rect 47952 2440 48004 2446
rect 47952 2382 48004 2388
rect 48412 2440 48464 2446
rect 48412 2382 48464 2388
rect 49424 2440 49476 2446
rect 49424 2382 49476 2388
rect 47964 800 47992 2382
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 48332 2038 48360 2246
rect 48320 2032 48372 2038
rect 48320 1974 48372 1980
rect 48424 800 48452 2382
rect 49436 800 49464 2382
rect 49896 800 49924 2790
rect 50896 2440 50948 2446
rect 50896 2382 50948 2388
rect 51356 2440 51408 2446
rect 51356 2382 51408 2388
rect 52368 2440 52420 2446
rect 52368 2382 52420 2388
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50908 800 50936 2382
rect 51368 800 51396 2382
rect 52380 800 52408 2382
rect 52840 800 52868 2790
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 52920 2304 52972 2310
rect 52920 2246 52972 2252
rect 52932 1562 52960 2246
rect 52920 1556 52972 1562
rect 52920 1498 52972 1504
rect 53852 800 53880 2382
rect 54116 2304 54168 2310
rect 54116 2246 54168 2252
rect 54128 1494 54156 2246
rect 54116 1488 54168 1494
rect 54116 1430 54168 1436
rect 54312 800 54340 2790
rect 55220 2440 55272 2446
rect 55220 2382 55272 2388
rect 55772 2440 55824 2446
rect 55772 2382 55824 2388
rect 55232 800 55260 2382
rect 55496 2304 55548 2310
rect 55496 2246 55548 2252
rect 55508 1630 55536 2246
rect 55496 1624 55548 1630
rect 55496 1566 55548 1572
rect 55784 800 55812 2382
rect 56704 800 56732 2994
rect 58716 2848 58768 2854
rect 58716 2790 58768 2796
rect 57244 2440 57296 2446
rect 57244 2382 57296 2388
rect 57256 800 57284 2382
rect 58164 2372 58216 2378
rect 58164 2314 58216 2320
rect 58176 800 58204 2314
rect 58728 800 58756 2790
rect 59648 800 59676 3402
rect 19812 734 20024 762
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
<< via2 >>
rect 2870 41656 2926 41712
rect 2778 40024 2834 40080
rect 1582 39244 1584 39264
rect 1584 39244 1636 39264
rect 1636 39244 1638 39264
rect 1582 39208 1638 39244
rect 1582 38392 1638 38448
rect 1398 26560 1454 26616
rect 1214 22380 1216 22400
rect 1216 22380 1268 22400
rect 1268 22380 1270 22400
rect 1214 22344 1270 22380
rect 1398 21528 1454 21584
rect 1582 37612 1584 37632
rect 1584 37612 1636 37632
rect 1636 37612 1638 37632
rect 1582 37576 1638 37612
rect 1582 36644 1638 36680
rect 1582 36624 1584 36644
rect 1584 36624 1636 36644
rect 1636 36624 1638 36644
rect 1582 35808 1638 35864
rect 1582 34992 1638 35048
rect 1582 34176 1638 34232
rect 1582 33804 1584 33824
rect 1584 33804 1636 33824
rect 1636 33804 1638 33824
rect 1582 33768 1638 33804
rect 1582 32952 1638 33008
rect 1582 32408 1638 32464
rect 1582 31592 1638 31648
rect 1582 31204 1638 31240
rect 1582 31184 1584 31204
rect 1584 31184 1636 31204
rect 1636 31184 1638 31204
rect 1582 30368 1638 30424
rect 1582 29996 1584 30016
rect 1584 29996 1636 30016
rect 1636 29996 1638 30016
rect 1582 29960 1638 29996
rect 1582 29144 1638 29200
rect 1582 28736 1638 28792
rect 1582 27376 1638 27432
rect 1582 26188 1584 26208
rect 1584 26188 1636 26208
rect 1636 26188 1638 26208
rect 1582 26152 1638 26188
rect 1582 25336 1638 25392
rect 1582 24928 1638 24984
rect 1582 24112 1638 24168
rect 1582 23704 1638 23760
rect 1582 21120 1638 21176
rect 1398 16496 1454 16552
rect 1582 20304 1638 20360
rect 1582 19932 1584 19952
rect 1584 19932 1636 19952
rect 1636 19932 1638 19952
rect 1582 19896 1638 19932
rect 1582 19080 1638 19136
rect 1582 18572 1584 18592
rect 1584 18572 1636 18592
rect 1636 18572 1638 18592
rect 1582 18536 1638 18572
rect 1582 17720 1638 17776
rect 1582 17332 1638 17368
rect 1582 17312 1584 17332
rect 1584 17312 1636 17332
rect 1636 17312 1638 17332
rect 2226 22752 2282 22808
rect 2226 20304 2282 20360
rect 1582 16088 1638 16144
rect 1582 15272 1638 15328
rect 1582 14884 1638 14920
rect 1582 14864 1584 14884
rect 1584 14864 1636 14884
rect 1636 14864 1638 14884
rect 1582 13912 1638 13968
rect 2502 20304 2558 20360
rect 3054 40840 3110 40896
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 3054 27784 3110 27840
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1582 13524 1638 13560
rect 1582 13504 1584 13524
rect 1584 13504 1636 13524
rect 1636 13504 1638 13524
rect 1582 12280 1638 12336
rect 3054 12688 3110 12744
rect 1582 11464 1638 11520
rect 1582 11056 1638 11112
rect 1582 10240 1638 10296
rect 1398 9832 1454 9888
rect 1674 9560 1730 9616
rect 2962 9596 2964 9616
rect 2964 9596 3016 9616
rect 3016 9596 3018 9616
rect 2962 9560 3018 9596
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 1582 8472 1638 8528
rect 2778 8064 2834 8120
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1582 7692 1584 7712
rect 1584 7692 1636 7712
rect 1636 7692 1638 7712
rect 1582 7656 1638 7692
rect 1490 6840 1546 6896
rect 1398 6432 1454 6488
rect 1582 6060 1584 6080
rect 1584 6060 1636 6080
rect 1636 6060 1638 6080
rect 1582 6024 1638 6060
rect 1582 4256 1638 4312
rect 1398 1808 1454 1864
rect 2870 2644 2926 2680
rect 2870 2624 2872 2644
rect 2872 2624 2924 2644
rect 2924 2624 2926 2644
rect 2778 2216 2834 2272
rect 1306 584 1362 640
rect 3514 4664 3570 4720
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3146 1400 3202 1456
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3068 4068 3088
rect 4068 3068 4120 3088
rect 4120 3068 4122 3088
rect 3238 992 3294 1048
rect 4066 3032 4122 3068
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 2962 176 3018 232
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 0 41714 800 41744
rect 2865 41714 2931 41717
rect 0 41712 2931 41714
rect 0 41656 2870 41712
rect 2926 41656 2931 41712
rect 0 41654 2931 41656
rect 0 41624 800 41654
rect 2865 41651 2931 41654
rect 0 41216 800 41336
rect 0 40898 800 40928
rect 3049 40898 3115 40901
rect 0 40896 3115 40898
rect 0 40840 3054 40896
rect 3110 40840 3115 40896
rect 0 40838 3115 40840
rect 0 40808 800 40838
rect 3049 40835 3115 40838
rect 0 40400 800 40520
rect 0 40082 800 40112
rect 2773 40082 2839 40085
rect 0 40080 2839 40082
rect 0 40024 2778 40080
rect 2834 40024 2839 40080
rect 0 40022 2839 40024
rect 0 39992 800 40022
rect 2773 40019 2839 40022
rect 4208 39744 4528 39745
rect 0 39584 800 39704
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39266 800 39296
rect 1577 39266 1643 39269
rect 0 39264 1643 39266
rect 0 39208 1582 39264
rect 1638 39208 1643 39264
rect 0 39206 1643 39208
rect 0 39176 800 39206
rect 1577 39203 1643 39206
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 0 38768 800 38888
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38450 800 38480
rect 1577 38450 1643 38453
rect 0 38448 1643 38450
rect 0 38392 1582 38448
rect 1638 38392 1643 38448
rect 0 38390 1643 38392
rect 0 38360 800 38390
rect 1577 38387 1643 38390
rect 19568 38112 19888 38113
rect 0 37952 800 38072
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 0 37634 800 37664
rect 1577 37634 1643 37637
rect 0 37632 1643 37634
rect 0 37576 1582 37632
rect 1638 37576 1643 37632
rect 0 37574 1643 37576
rect 0 37544 800 37574
rect 1577 37571 1643 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 0 37000 800 37120
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 0 36682 800 36712
rect 1577 36682 1643 36685
rect 0 36680 1643 36682
rect 0 36624 1582 36680
rect 1638 36624 1643 36680
rect 0 36622 1643 36624
rect 0 36592 800 36622
rect 1577 36619 1643 36622
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36184 800 36304
rect 19568 35936 19888 35937
rect 0 35866 800 35896
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 1577 35866 1643 35869
rect 0 35864 1643 35866
rect 0 35808 1582 35864
rect 1638 35808 1643 35864
rect 0 35806 1643 35808
rect 0 35776 800 35806
rect 1577 35803 1643 35806
rect 0 35368 800 35488
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 35050 800 35080
rect 1577 35050 1643 35053
rect 0 35048 1643 35050
rect 0 34992 1582 35048
rect 1638 34992 1643 35048
rect 0 34990 1643 34992
rect 0 34960 800 34990
rect 1577 34987 1643 34990
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 0 34552 800 34672
rect 4208 34304 4528 34305
rect 0 34234 800 34264
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 1577 34234 1643 34237
rect 0 34232 1643 34234
rect 0 34176 1582 34232
rect 1638 34176 1643 34232
rect 0 34174 1643 34176
rect 0 34144 800 34174
rect 1577 34171 1643 34174
rect 0 33826 800 33856
rect 1577 33826 1643 33829
rect 0 33824 1643 33826
rect 0 33768 1582 33824
rect 1638 33768 1643 33824
rect 0 33766 1643 33768
rect 0 33736 800 33766
rect 1577 33763 1643 33766
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 0 33328 800 33448
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 33010 800 33040
rect 1577 33010 1643 33013
rect 0 33008 1643 33010
rect 0 32952 1582 33008
rect 1638 32952 1643 33008
rect 0 32950 1643 32952
rect 0 32920 800 32950
rect 1577 32947 1643 32950
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 0 32466 800 32496
rect 1577 32466 1643 32469
rect 0 32464 1643 32466
rect 0 32408 1582 32464
rect 1638 32408 1643 32464
rect 0 32406 1643 32408
rect 0 32376 800 32406
rect 1577 32403 1643 32406
rect 4208 32128 4528 32129
rect 0 31968 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 0 31650 800 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 800 31590
rect 1577 31587 1643 31590
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31242 800 31272
rect 1577 31242 1643 31245
rect 0 31240 1643 31242
rect 0 31184 1582 31240
rect 1638 31184 1643 31240
rect 0 31182 1643 31184
rect 0 31152 800 31182
rect 1577 31179 1643 31182
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30744 800 30864
rect 19568 30496 19888 30497
rect 0 30426 800 30456
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 1577 30426 1643 30429
rect 0 30424 1643 30426
rect 0 30368 1582 30424
rect 1638 30368 1643 30424
rect 0 30366 1643 30368
rect 0 30336 800 30366
rect 1577 30363 1643 30366
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 0 29520 800 29640
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 0 29202 800 29232
rect 1577 29202 1643 29205
rect 0 29200 1643 29202
rect 0 29144 1582 29200
rect 1638 29144 1643 29200
rect 0 29142 1643 29144
rect 0 29112 800 29142
rect 1577 29139 1643 29142
rect 4208 28864 4528 28865
rect 0 28794 800 28824
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 1577 28794 1643 28797
rect 0 28792 1643 28794
rect 0 28736 1582 28792
rect 1638 28736 1643 28792
rect 0 28734 1643 28736
rect 0 28704 800 28734
rect 1577 28731 1643 28734
rect 0 28296 800 28416
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 0 27842 800 27872
rect 3049 27842 3115 27845
rect 0 27840 3115 27842
rect 0 27784 3054 27840
rect 3110 27784 3115 27840
rect 0 27782 3115 27784
rect 0 27752 800 27782
rect 3049 27779 3115 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27434 800 27464
rect 1577 27434 1643 27437
rect 0 27432 1643 27434
rect 0 27376 1582 27432
rect 1638 27376 1643 27432
rect 0 27374 1643 27376
rect 0 27344 800 27374
rect 1577 27371 1643 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 0 26936 800 27056
rect 4208 26688 4528 26689
rect 0 26618 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 1393 26618 1459 26621
rect 0 26616 1459 26618
rect 0 26560 1398 26616
rect 1454 26560 1459 26616
rect 0 26558 1459 26560
rect 0 26528 800 26558
rect 1393 26555 1459 26558
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 0 25712 800 25832
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25394 800 25424
rect 1577 25394 1643 25397
rect 0 25392 1643 25394
rect 0 25336 1582 25392
rect 1638 25336 1643 25392
rect 0 25334 1643 25336
rect 0 25304 800 25334
rect 1577 25331 1643 25334
rect 19568 25056 19888 25057
rect 0 24986 800 25016
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 800 24926
rect 1577 24923 1643 24926
rect 0 24488 800 24608
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 0 23762 800 23792
rect 1577 23762 1643 23765
rect 0 23760 1643 23762
rect 0 23704 1582 23760
rect 1638 23704 1643 23760
rect 0 23702 1643 23704
rect 0 23672 800 23702
rect 1577 23699 1643 23702
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23128 800 23248
rect 19568 22880 19888 22881
rect 0 22810 800 22840
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 2221 22810 2287 22813
rect 0 22808 2287 22810
rect 0 22752 2226 22808
rect 2282 22752 2287 22808
rect 0 22750 2287 22752
rect 0 22720 800 22750
rect 2221 22747 2287 22750
rect 0 22402 800 22432
rect 1209 22402 1275 22405
rect 0 22400 1275 22402
rect 0 22344 1214 22400
rect 1270 22344 1275 22400
rect 0 22342 1275 22344
rect 0 22312 800 22342
rect 1209 22339 1275 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21904 800 22024
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 0 21586 800 21616
rect 1393 21586 1459 21589
rect 0 21584 1459 21586
rect 0 21528 1398 21584
rect 1454 21528 1459 21584
rect 0 21526 1459 21528
rect 0 21496 800 21526
rect 1393 21523 1459 21526
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 1577 21178 1643 21181
rect 0 21176 1643 21178
rect 0 21120 1582 21176
rect 1638 21120 1643 21176
rect 0 21118 1643 21120
rect 0 21088 800 21118
rect 1577 21115 1643 21118
rect 0 20680 800 20800
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 0 20362 800 20392
rect 1577 20362 1643 20365
rect 0 20360 1643 20362
rect 0 20304 1582 20360
rect 1638 20304 1643 20360
rect 0 20302 1643 20304
rect 0 20272 800 20302
rect 1577 20299 1643 20302
rect 2221 20362 2287 20365
rect 2497 20362 2563 20365
rect 2221 20360 2563 20362
rect 2221 20304 2226 20360
rect 2282 20304 2502 20360
rect 2558 20304 2563 20360
rect 2221 20302 2563 20304
rect 2221 20299 2287 20302
rect 2497 20299 2563 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19954 800 19984
rect 1577 19954 1643 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 800 19894
rect 1577 19891 1643 19894
rect 19568 19616 19888 19617
rect 0 19456 800 19576
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 0 19138 800 19168
rect 1577 19138 1643 19141
rect 0 19136 1643 19138
rect 0 19080 1582 19136
rect 1638 19080 1643 19136
rect 0 19078 1643 19080
rect 0 19048 800 19078
rect 1577 19075 1643 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 0 18594 800 18624
rect 1577 18594 1643 18597
rect 0 18592 1643 18594
rect 0 18536 1582 18592
rect 1638 18536 1643 18592
rect 0 18534 1643 18536
rect 0 18504 800 18534
rect 1577 18531 1643 18534
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 0 18096 800 18216
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 800 17718
rect 1577 17715 1643 17718
rect 19568 17440 19888 17441
rect 0 17370 800 17400
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 0 16872 800 16992
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16554 800 16584
rect 1393 16554 1459 16557
rect 0 16552 1459 16554
rect 0 16496 1398 16552
rect 1454 16496 1459 16552
rect 0 16494 1459 16496
rect 0 16464 800 16494
rect 1393 16491 1459 16494
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 4208 15808 4528 15809
rect 0 15648 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 0 14922 800 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 800 14862
rect 1577 14859 1643 14862
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14424 800 14544
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 4208 13632 4528 13633
rect 0 13562 800 13592
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 1577 13562 1643 13565
rect 0 13560 1643 13562
rect 0 13504 1582 13560
rect 1638 13504 1643 13560
rect 0 13502 1643 13504
rect 0 13472 800 13502
rect 1577 13499 1643 13502
rect 0 13064 800 13184
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 0 12746 800 12776
rect 3049 12746 3115 12749
rect 0 12744 3115 12746
rect 0 12688 3054 12744
rect 3110 12688 3115 12744
rect 0 12686 3115 12688
rect 0 12656 800 12686
rect 3049 12683 3115 12686
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 19568 12000 19888 12001
rect 0 11840 800 11960
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 0 11522 800 11552
rect 1577 11522 1643 11525
rect 0 11520 1643 11522
rect 0 11464 1582 11520
rect 1638 11464 1643 11520
rect 0 11462 1643 11464
rect 0 11432 800 11462
rect 1577 11459 1643 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 11114 800 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 800 11054
rect 1577 11051 1643 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 0 10616 800 10736
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10208 800 10238
rect 1577 10235 1643 10238
rect 0 9890 800 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 800 9830
rect 1393 9827 1459 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 1669 9618 1735 9621
rect 2957 9618 3023 9621
rect 1669 9616 3023 9618
rect 1669 9560 1674 9616
rect 1730 9560 2962 9616
rect 3018 9560 3023 9616
rect 1669 9558 3023 9560
rect 1669 9555 1735 9558
rect 2957 9555 3023 9558
rect 0 9346 800 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 800 9286
rect 1577 9283 1643 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8848 800 8968
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 0 8530 800 8560
rect 1577 8530 1643 8533
rect 0 8528 1643 8530
rect 0 8472 1582 8528
rect 1638 8472 1643 8528
rect 0 8470 1643 8472
rect 0 8440 800 8470
rect 1577 8467 1643 8470
rect 4208 8192 4528 8193
rect 0 8122 800 8152
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 2773 8122 2839 8125
rect 0 8120 2839 8122
rect 0 8064 2778 8120
rect 2834 8064 2839 8120
rect 0 8062 2839 8064
rect 0 8032 800 8062
rect 2773 8059 2839 8062
rect 0 7714 800 7744
rect 1577 7714 1643 7717
rect 0 7712 1643 7714
rect 0 7656 1582 7712
rect 1638 7656 1643 7712
rect 0 7654 1643 7656
rect 0 7624 800 7654
rect 1577 7651 1643 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 0 7216 800 7336
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 19568 6560 19888 6561
rect 0 6490 800 6520
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 1393 6490 1459 6493
rect 0 6488 1459 6490
rect 0 6432 1398 6488
rect 1454 6432 1459 6488
rect 0 6430 1459 6432
rect 0 6400 800 6430
rect 1393 6427 1459 6430
rect 0 6082 800 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 800 6022
rect 1577 6019 1643 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5584 800 5704
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 0 5176 800 5296
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 0 4722 800 4752
rect 3509 4722 3575 4725
rect 0 4720 3575 4722
rect 0 4664 3514 4720
rect 3570 4664 3575 4720
rect 0 4662 3575 4664
rect 0 4632 800 4662
rect 3509 4659 3575 4662
rect 19568 4384 19888 4385
rect 0 4314 800 4344
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 1577 4314 1643 4317
rect 0 4312 1643 4314
rect 0 4256 1582 4312
rect 1638 4256 1643 4312
rect 0 4254 1643 4256
rect 0 4224 800 4254
rect 1577 4251 1643 4254
rect 0 3816 800 3936
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3408 800 3528
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 0 3090 800 3120
rect 4061 3090 4127 3093
rect 0 3088 4127 3090
rect 0 3032 4066 3088
rect 4122 3032 4127 3088
rect 0 3030 4127 3032
rect 0 3000 800 3030
rect 4061 3027 4127 3030
rect 4208 2752 4528 2753
rect 0 2682 800 2712
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 2865 2682 2931 2685
rect 0 2680 2931 2682
rect 0 2624 2870 2680
rect 2926 2624 2931 2680
rect 0 2622 2931 2624
rect 0 2592 800 2622
rect 2865 2619 2931 2622
rect 0 2274 800 2304
rect 2773 2274 2839 2277
rect 0 2272 2839 2274
rect 0 2216 2778 2272
rect 2834 2216 2839 2272
rect 0 2214 2839 2216
rect 0 2184 800 2214
rect 2773 2211 2839 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 0 1866 800 1896
rect 1393 1866 1459 1869
rect 0 1864 1459 1866
rect 0 1808 1398 1864
rect 1454 1808 1459 1864
rect 0 1806 1459 1808
rect 0 1776 800 1806
rect 1393 1803 1459 1806
rect 0 1458 800 1488
rect 3141 1458 3207 1461
rect 0 1456 3207 1458
rect 0 1400 3146 1456
rect 3202 1400 3207 1456
rect 0 1398 3207 1400
rect 0 1368 800 1398
rect 3141 1395 3207 1398
rect 0 1050 800 1080
rect 3233 1050 3299 1053
rect 0 1048 3299 1050
rect 0 992 3238 1048
rect 3294 992 3299 1048
rect 0 990 3299 992
rect 0 960 800 990
rect 3233 987 3299 990
rect 0 642 800 672
rect 1301 642 1367 645
rect 0 640 1367 642
rect 0 584 1306 640
rect 1362 584 1367 640
rect 0 582 1367 584
rect 0 552 800 582
rect 1301 579 1367 582
rect 0 234 800 264
rect 2957 234 3023 237
rect 0 232 3023 234
rect 0 176 2962 232
rect 3018 176 3023 232
rect 0 174 3023 176
rect 0 144 800 174
rect 2957 171 3023 174
<< via3 >>
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 39744 4528 39760
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 39200 19888 39760
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 39744 35248 39760
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 39200 50608 39760
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__decap_8  FILLER_0_19 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1644511149
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47
timestamp 1644511149
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74
timestamp 1644511149
transform 1 0 7912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1644511149
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1644511149
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 1644511149
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_144
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1644511149
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1644511149
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1644511149
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1644511149
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_244
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_260
timestamp 1644511149
transform 1 0 25024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_267
timestamp 1644511149
transform 1 0 25668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_284
timestamp 1644511149
transform 1 0 27232 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_292
timestamp 1644511149
transform 1 0 27968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_296
timestamp 1644511149
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_300
timestamp 1644511149
transform 1 0 28704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_312
timestamp 1644511149
transform 1 0 29808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_316
timestamp 1644511149
transform 1 0 30176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1644511149
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1644511149
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_347
timestamp 1644511149
transform 1 0 33028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_355
timestamp 1644511149
transform 1 0 33764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1644511149
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1644511149
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1644511149
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1644511149
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_425
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_434
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_441
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1644511149
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1644511149
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1644511149
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1644511149
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_493
timestamp 1644511149
transform 1 0 46460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1644511149
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_509
timestamp 1644511149
transform 1 0 47932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_514
timestamp 1644511149
transform 1 0 48392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_521
timestamp 1644511149
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_537
timestamp 1644511149
transform 1 0 50508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_541
timestamp 1644511149
transform 1 0 50876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_546
timestamp 1644511149
transform 1 0 51336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_553
timestamp 1644511149
transform 1 0 51980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1644511149
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_565
timestamp 1644511149
transform 1 0 53084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1644511149
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1644511149
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_593
timestamp 1644511149
transform 1 0 55660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_600
timestamp 1644511149
transform 1 0 56304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1644511149
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1644511149
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1644511149
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1644511149
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1644511149
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1644511149
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1644511149
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1644511149
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_130
timestamp 1644511149
transform 1 0 13064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1644511149
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_151
timestamp 1644511149
transform 1 0 14996 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_176
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_186
timestamp 1644511149
transform 1 0 18216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1644511149
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_203 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19780 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_215
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_228
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_244
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_248
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_260
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1644511149
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_290
timestamp 1644511149
transform 1 0 27784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_302
timestamp 1644511149
transform 1 0 28888 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_314
timestamp 1644511149
transform 1 0 29992 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1644511149
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1644511149
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_343
timestamp 1644511149
transform 1 0 32660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_369
timestamp 1644511149
transform 1 0 35052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_375
timestamp 1644511149
transform 1 0 35604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1644511149
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_396
timestamp 1644511149
transform 1 0 37536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_408
timestamp 1644511149
transform 1 0 38640 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_423
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_435
timestamp 1644511149
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_455
timestamp 1644511149
transform 1 0 42964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_467
timestamp 1644511149
transform 1 0 44068 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_471
timestamp 1644511149
transform 1 0 44436 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_483
timestamp 1644511149
transform 1 0 45540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1644511149
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_508
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_520
timestamp 1644511149
transform 1 0 48944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_528
timestamp 1644511149
transform 1 0 49680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_534
timestamp 1644511149
transform 1 0 50232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_546
timestamp 1644511149
transform 1 0 51336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1644511149
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_566
timestamp 1644511149
transform 1 0 53176 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_578
timestamp 1644511149
transform 1 0 54280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_582
timestamp 1644511149
transform 1 0 54648 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_594
timestamp 1644511149
transform 1 0 55752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_602
timestamp 1644511149
transform 1 0 56488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1644511149
transform 1 0 58236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1644511149
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1644511149
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_100
timestamp 1644511149
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1644511149
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1644511149
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_178
timestamp 1644511149
transform 1 0 17480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_212
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1644511149
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1644511149
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_66
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_78
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_100
timestamp 1644511149
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_194
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_204
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_13
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1644511149
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_60
timestamp 1644511149
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_72
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_101
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_115
timestamp 1644511149
transform 1 0 11684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1644511149
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1644511149
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_207
timestamp 1644511149
transform 1 0 20148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_219
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_231
timestamp 1644511149
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1644511149
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_256
timestamp 1644511149
transform 1 0 24656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_268
timestamp 1644511149
transform 1 0 25760 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1644511149
transform 1 0 26864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_292
timestamp 1644511149
transform 1 0 27968 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1644511149
transform 1 0 6808 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1644511149
transform 1 0 7912 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_86
timestamp 1644511149
transform 1 0 9016 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1644511149
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1644511149
transform 1 0 12972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1644511149
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1644511149
transform 1 0 14996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1644511149
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_175
timestamp 1644511149
transform 1 0 17204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1644511149
transform 1 0 19136 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_6
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1644511149
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1644511149
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_159
timestamp 1644511149
transform 1 0 15732 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_185
timestamp 1644511149
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1644511149
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_30
timestamp 1644511149
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_42
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1644511149
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_63
timestamp 1644511149
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1644511149
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1644511149
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_92
timestamp 1644511149
transform 1 0 9568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_100
timestamp 1644511149
transform 1 0 10304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1644511149
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_143
timestamp 1644511149
transform 1 0 14260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1644511149
transform 1 0 14996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1644511149
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1644511149
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_194
timestamp 1644511149
transform 1 0 18952 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_206
timestamp 1644511149
transform 1 0 20056 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1644511149
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1644511149
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1644511149
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_47
timestamp 1644511149
transform 1 0 5428 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_56
timestamp 1644511149
transform 1 0 6256 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_71
timestamp 1644511149
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp 1644511149
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_96
timestamp 1644511149
transform 1 0 9936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_113
timestamp 1644511149
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_125
timestamp 1644511149
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1644511149
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_159
timestamp 1644511149
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1644511149
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1644511149
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_19
timestamp 1644511149
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 1644511149
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1644511149
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_66
timestamp 1644511149
transform 1 0 7176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1644511149
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_89
timestamp 1644511149
transform 1 0 9292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1644511149
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1644511149
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_147
timestamp 1644511149
transform 1 0 14628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp 1644511149
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1644511149
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp 1644511149
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1644511149
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_194
timestamp 1644511149
transform 1 0 18952 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_206
timestamp 1644511149
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1644511149
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1644511149
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1644511149
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_126
timestamp 1644511149
transform 1 0 12696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_147
timestamp 1644511149
transform 1 0 14628 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_159
timestamp 1644511149
transform 1 0 15732 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_171
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_203
timestamp 1644511149
transform 1 0 19780 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1644511149
transform 1 0 20884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1644511149
transform 1 0 21988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1644511149
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1644511149
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_60
timestamp 1644511149
transform 1 0 6624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_77
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_89
timestamp 1644511149
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1644511149
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_119
timestamp 1644511149
transform 1 0 12052 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_127
timestamp 1644511149
transform 1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_146
timestamp 1644511149
transform 1 0 14536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1644511149
transform 1 0 17204 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_183
timestamp 1644511149
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_195
timestamp 1644511149
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1644511149
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1644511149
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1644511149
transform 1 0 2852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1644511149
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1644511149
transform 1 0 7360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1644511149
transform 1 0 10120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1644511149
transform 1 0 10488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_119
timestamp 1644511149
transform 1 0 12052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1644511149
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_164
timestamp 1644511149
transform 1 0 16192 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_176
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1644511149
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_203
timestamp 1644511149
transform 1 0 19780 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1644511149
transform 1 0 20884 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1644511149
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1644511149
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_31
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1644511149
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_60
timestamp 1644511149
transform 1 0 6624 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_72
timestamp 1644511149
transform 1 0 7728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1644511149
transform 1 0 9016 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_94
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1644511149
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_185
timestamp 1644511149
transform 1 0 18124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_197
timestamp 1644511149
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_209
timestamp 1644511149
transform 1 0 20332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1644511149
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1644511149
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_48
timestamp 1644511149
transform 1 0 5520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1644511149
transform 1 0 11868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_125
timestamp 1644511149
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1644511149
transform 1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_25
timestamp 1644511149
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1644511149
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1644511149
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_77
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_85
timestamp 1644511149
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_97
timestamp 1644511149
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1644511149
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_141
timestamp 1644511149
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_153
timestamp 1644511149
transform 1 0 15180 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1644511149
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1644511149
transform 1 0 18032 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1644511149
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1644511149
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1644511149
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1644511149
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1644511149
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_123
timestamp 1644511149
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1644511149
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_162
timestamp 1644511149
transform 1 0 16008 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1644511149
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_24
timestamp 1644511149
transform 1 0 3312 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_77
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_85
timestamp 1644511149
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_97
timestamp 1644511149
transform 1 0 10028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1644511149
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_121
timestamp 1644511149
transform 1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_129
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_138
timestamp 1644511149
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1644511149
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1644511149
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_177
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_201
timestamp 1644511149
transform 1 0 19596 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1644511149
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1644511149
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_6
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1644511149
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_38
timestamp 1644511149
transform 1 0 4600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_50
timestamp 1644511149
transform 1 0 5704 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_72
timestamp 1644511149
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_104
timestamp 1644511149
transform 1 0 10672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_112
timestamp 1644511149
transform 1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1644511149
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_146
timestamp 1644511149
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_158
timestamp 1644511149
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1644511149
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1644511149
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1644511149
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1644511149
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_22
timestamp 1644511149
transform 1 0 3128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_30
timestamp 1644511149
transform 1 0 3864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_42
timestamp 1644511149
transform 1 0 4968 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_48
timestamp 1644511149
transform 1 0 5520 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1644511149
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1644511149
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1644511149
transform 1 0 8280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_82
timestamp 1644511149
transform 1 0 8648 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1644511149
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1644511149
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_148
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_156
timestamp 1644511149
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_189
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_201
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_213
timestamp 1644511149
transform 1 0 20700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1644511149
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 1644511149
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_37
timestamp 1644511149
transform 1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1644511149
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_63
timestamp 1644511149
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1644511149
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1644511149
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_108
timestamp 1644511149
transform 1 0 11040 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_120
timestamp 1644511149
transform 1 0 12144 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_147
timestamp 1644511149
transform 1 0 14628 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_159
timestamp 1644511149
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1644511149
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_33
timestamp 1644511149
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_45
timestamp 1644511149
transform 1 0 5244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_152
timestamp 1644511149
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_185
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_197
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_209
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_6
timestamp 1644511149
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_12
timestamp 1644511149
transform 1 0 2208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1644511149
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_37
timestamp 1644511149
transform 1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_45
timestamp 1644511149
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_55
timestamp 1644511149
transform 1 0 6164 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_67
timestamp 1644511149
transform 1 0 7268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1644511149
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1644511149
transform 1 0 10488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1644511149
transform 1 0 11316 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 1644511149
transform 1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 1644511149
transform 1 0 13156 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_151
timestamp 1644511149
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_163
timestamp 1644511149
transform 1 0 16100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1644511149
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_11
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_79
timestamp 1644511149
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1644511149
transform 1 0 9476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1644511149
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1644511149
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_191
timestamp 1644511149
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_203
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1644511149
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_10
timestamp 1644511149
transform 1 0 2024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1644511149
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_62
timestamp 1644511149
transform 1 0 6808 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1644511149
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1644511149
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1644511149
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_150
timestamp 1644511149
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_162
timestamp 1644511149
transform 1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1644511149
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_26
timestamp 1644511149
transform 1 0 3496 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_38
timestamp 1644511149
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1644511149
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_65
timestamp 1644511149
transform 1 0 7084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_75
timestamp 1644511149
transform 1 0 8004 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1644511149
transform 1 0 9108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_99
timestamp 1644511149
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1644511149
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_150
timestamp 1644511149
transform 1 0 14904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_49
timestamp 1644511149
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_61
timestamp 1644511149
transform 1 0 6716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_72
timestamp 1644511149
transform 1 0 7728 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1644511149
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_115
timestamp 1644511149
transform 1 0 11684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1644511149
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_182
timestamp 1644511149
transform 1 0 17848 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1644511149
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_19
timestamp 1644511149
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_31
timestamp 1644511149
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_43
timestamp 1644511149
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1644511149
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_72
timestamp 1644511149
transform 1 0 7728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_84
timestamp 1644511149
transform 1 0 8832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1644511149
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_104
timestamp 1644511149
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_187
timestamp 1644511149
transform 1 0 18308 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_211
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_49
timestamp 1644511149
transform 1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1644511149
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1644511149
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_150
timestamp 1644511149
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_162
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_168
timestamp 1644511149
transform 1 0 16560 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_185
timestamp 1644511149
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1644511149
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_6
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1644511149
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1644511149
transform 1 0 8648 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1644511149
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1644511149
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1644511149
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_7
timestamp 1644511149
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_48
timestamp 1644511149
transform 1 0 5520 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_60
timestamp 1644511149
transform 1 0 6624 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 1644511149
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1644511149
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_89
timestamp 1644511149
transform 1 0 9292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_101
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1644511149
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_148
timestamp 1644511149
transform 1 0 14720 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_172
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_184
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_6
timestamp 1644511149
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_18
timestamp 1644511149
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_30
timestamp 1644511149
transform 1 0 3864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1644511149
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_64
timestamp 1644511149
transform 1 0 6992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1644511149
transform 1 0 7912 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_86
timestamp 1644511149
transform 1 0 9016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_97
timestamp 1644511149
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1644511149
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1644511149
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_132
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_144
timestamp 1644511149
transform 1 0 14352 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1644511149
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1644511149
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_73
timestamp 1644511149
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1644511149
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_152
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_164
timestamp 1644511149
transform 1 0 16192 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_176
timestamp 1644511149
transform 1 0 17296 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1644511149
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_25
timestamp 1644511149
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_37
timestamp 1644511149
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1644511149
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp 1644511149
transform 1 0 7084 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_73
timestamp 1644511149
transform 1 0 7820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1644511149
transform 1 0 8648 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1644511149
transform 1 0 9752 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1644511149
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_121
timestamp 1644511149
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_141
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_153
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1644511149
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_6
timestamp 1644511149
transform 1 0 1656 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_33
timestamp 1644511149
transform 1 0 4140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_44
timestamp 1644511149
transform 1 0 5152 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_52
timestamp 1644511149
transform 1 0 5888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_71
timestamp 1644511149
transform 1 0 7636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_95
timestamp 1644511149
transform 1 0 9844 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_107
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1644511149
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_160
timestamp 1644511149
transform 1 0 15824 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_184
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_11
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_21
timestamp 1644511149
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_33
timestamp 1644511149
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1644511149
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1644511149
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_89
timestamp 1644511149
transform 1 0 9292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_35
timestamp 1644511149
transform 1 0 4324 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_45
timestamp 1644511149
transform 1 0 5244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_57
timestamp 1644511149
transform 1 0 6348 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_63
timestamp 1644511149
transform 1 0 6900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_23
timestamp 1644511149
transform 1 0 3220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1644511149
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_41
timestamp 1644511149
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1644511149
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1644511149
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_13
timestamp 1644511149
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1644511149
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_21
timestamp 1644511149
transform 1 0 3036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_29
timestamp 1644511149
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1644511149
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1644511149
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_6
timestamp 1644511149
transform 1 0 1656 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_34
timestamp 1644511149
transform 1 0 4232 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_46
timestamp 1644511149
transform 1 0 5336 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1644511149
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1644511149
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_45
timestamp 1644511149
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_57
timestamp 1644511149
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_69
timestamp 1644511149
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1644511149
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_6
timestamp 1644511149
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_18
timestamp 1644511149
transform 1 0 2760 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_26
timestamp 1644511149
transform 1 0 3496 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_31
timestamp 1644511149
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_43
timestamp 1644511149
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1644511149
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_35
timestamp 1644511149
transform 1 0 4324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_47
timestamp 1644511149
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_59
timestamp 1644511149
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_71
timestamp 1644511149
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_23
timestamp 1644511149
transform 1 0 3220 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_34
timestamp 1644511149
transform 1 0 4232 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_46
timestamp 1644511149
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1644511149
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_11
timestamp 1644511149
transform 1 0 2116 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1644511149
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_49
timestamp 1644511149
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_73
timestamp 1644511149
transform 1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1644511149
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_6
timestamp 1644511149
transform 1 0 1656 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_12
timestamp 1644511149
transform 1 0 2208 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_16
timestamp 1644511149
transform 1 0 2576 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_24
timestamp 1644511149
transform 1 0 3312 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_35
timestamp 1644511149
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1644511149
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_7
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_13
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_23
timestamp 1644511149
transform 1 0 3220 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_6
timestamp 1644511149
transform 1 0 1656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_18
timestamp 1644511149
transform 1 0 2760 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1644511149
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_38
timestamp 1644511149
transform 1 0 4600 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_50
timestamp 1644511149
transform 1 0 5704 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_62
timestamp 1644511149
transform 1 0 6808 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_74
timestamp 1644511149
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1644511149
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_7
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_18
timestamp 1644511149
transform 1 0 2760 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_38
timestamp 1644511149
transform 1 0 4600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1644511149
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_6
timestamp 1644511149
transform 1 0 1656 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_14
timestamp 1644511149
transform 1 0 2392 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_7
timestamp 1644511149
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_35
timestamp 1644511149
transform 1 0 4324 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1644511149
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1644511149
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_18
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1644511149
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_37
timestamp 1644511149
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_43
timestamp 1644511149
transform 1 0 5060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_55
timestamp 1644511149
transform 1 0 6164 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_67
timestamp 1644511149
transform 1 0 7268 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1644511149
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_13
timestamp 1644511149
transform 1 0 2300 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_23
timestamp 1644511149
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_35
timestamp 1644511149
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_46
timestamp 1644511149
transform 1 0 5336 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_58
timestamp 1644511149
transform 1 0 6440 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_70
timestamp 1644511149
transform 1 0 7544 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1644511149
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_6
timestamp 1644511149
transform 1 0 1656 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1644511149
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_6
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_18
timestamp 1644511149
transform 1 0 2760 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1644511149
transform 1 0 3864 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_42
timestamp 1644511149
transform 1 0 4968 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1644511149
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1644511149
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_31
timestamp 1644511149
transform 1 0 3956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_43
timestamp 1644511149
transform 1 0 5060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_7
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_19
timestamp 1644511149
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_31
timestamp 1644511149
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_43
timestamp 1644511149
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_517
timestamp 1644511149
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_529
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_541
timestamp 1644511149
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1644511149
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_7
timestamp 1644511149
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1644511149
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_513
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_545
timestamp 1644511149
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_557
timestamp 1644511149
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_569
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1644511149
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1644511149
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_7
timestamp 1644511149
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_19
timestamp 1644511149
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_529
timestamp 1644511149
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_541
timestamp 1644511149
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1644511149
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_23
timestamp 1644511149
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1644511149
transform 1 0 4048 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1644511149
transform 1 0 5152 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_57
timestamp 1644511149
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_69
timestamp 1644511149
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1644511149
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_113
timestamp 1644511149
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_125
timestamp 1644511149
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 1644511149
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_169
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_181
timestamp 1644511149
transform 1 0 17756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1644511149
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_200
timestamp 1644511149
transform 1 0 19504 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_212
timestamp 1644511149
transform 1 0 20608 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_225
timestamp 1644511149
transform 1 0 21804 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_237
timestamp 1644511149
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1644511149
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_276
timestamp 1644511149
transform 1 0 26496 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_281
timestamp 1644511149
transform 1 0 26956 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_293
timestamp 1644511149
transform 1 0 28060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1644511149
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1644511149
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_349
timestamp 1644511149
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1644511149
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_393
timestamp 1644511149
transform 1 0 37260 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_405
timestamp 1644511149
transform 1 0 38364 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_417
timestamp 1644511149
transform 1 0 39468 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_439
timestamp 1644511149
transform 1 0 41492 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_447
timestamp 1644511149
transform 1 0 42228 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_449
timestamp 1644511149
transform 1 0 42412 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_461
timestamp 1644511149
transform 1 0 43516 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1644511149
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_505
timestamp 1644511149
transform 1 0 47564 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_517
timestamp 1644511149
transform 1 0 48668 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_521
timestamp 1644511149
transform 1 0 49036 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_529
timestamp 1644511149
transform 1 0 49772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_561
timestamp 1644511149
transform 1 0 52716 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_573
timestamp 1644511149
transform 1 0 53820 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_585
timestamp 1644511149
transform 1 0 54924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_597
timestamp 1644511149
transform 1 0 56028 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_602
timestamp 1644511149
transform 1 0 56488 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_614
timestamp 1644511149
transform 1 0 57592 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_617
timestamp 1644511149
transform 1 0 57868 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1644511149
transform 1 0 16836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 42320 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 47472 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 52624 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 57776 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _220_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _221_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _222_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _223_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _224_
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _225_
timestamp 1644511149
transform 1 0 14628 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _226_
timestamp 1644511149
transform 1 0 12328 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1644511149
transform 1 0 14260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _228_
timestamp 1644511149
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _229_
timestamp 1644511149
transform 1 0 12788 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _230_
timestamp 1644511149
transform 1 0 14444 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _231_
timestamp 1644511149
transform 1 0 12788 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _232_
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _233_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9016 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _234_
timestamp 1644511149
transform 1 0 9384 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _235_
timestamp 1644511149
transform 1 0 14444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _236_
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1644511149
transform 1 0 7360 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _238_
timestamp 1644511149
transform 1 0 17112 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _239_
timestamp 1644511149
transform 1 0 14076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _240_
timestamp 1644511149
transform 1 0 7728 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _241_
timestamp 1644511149
transform 1 0 7360 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _242_
timestamp 1644511149
transform 1 0 8188 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _243_
timestamp 1644511149
transform 1 0 13156 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _244_
timestamp 1644511149
transform 1 0 7268 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _245_
timestamp 1644511149
transform 1 0 8004 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _246_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _247_
timestamp 1644511149
transform 1 0 8004 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _248_
timestamp 1644511149
transform 1 0 6532 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _249_
timestamp 1644511149
transform 1 0 14996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _250_
timestamp 1644511149
transform 1 0 7360 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1644511149
transform 1 0 9568 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1644511149
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _253_
timestamp 1644511149
transform 1 0 7268 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _254_
timestamp 1644511149
transform 1 0 18124 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _255_
timestamp 1644511149
transform 1 0 18400 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _256_
timestamp 1644511149
transform 1 0 7728 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _257_
timestamp 1644511149
transform 1 0 10212 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _258_
timestamp 1644511149
transform 1 0 17572 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _259_
timestamp 1644511149
transform 1 0 19412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _260_
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _261_
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _262_
timestamp 1644511149
transform 1 0 10304 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _263_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1644511149
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _265_
timestamp 1644511149
transform 1 0 7268 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _266_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _267_
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _268_
timestamp 1644511149
transform 1 0 6624 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _269_
timestamp 1644511149
transform 1 0 20332 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1644511149
transform 1 0 7452 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _271_
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _272_
timestamp 1644511149
transform 1 0 17664 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _273_
timestamp 1644511149
transform 1 0 9844 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _274_
timestamp 1644511149
transform 1 0 9292 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _275_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _276_
timestamp 1644511149
transform 1 0 10120 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _277_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _278_
timestamp 1644511149
transform 1 0 15640 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _279_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _280_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _281_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6808 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _282_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1932 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _283_
timestamp 1644511149
transform 1 0 2944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _284_
timestamp 1644511149
transform 1 0 3220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _285_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp 1644511149
transform 1 0 2576 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _291_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _292_
timestamp 1644511149
transform 1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1644511149
transform 1 0 2208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1644511149
transform 1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1644511149
transform 1 0 4324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1644511149
transform 1 0 2300 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _301_
timestamp 1644511149
transform 1 0 5336 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1644511149
transform 1 0 5520 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _303_
timestamp 1644511149
transform 1 0 4140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _304_
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1644511149
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1644511149
transform 1 0 2208 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1644511149
transform 1 0 2208 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1644511149
transform 1 0 2208 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _310_
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1644511149
transform 1 0 2208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _312_
timestamp 1644511149
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1644511149
transform 1 0 4600 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1644511149
transform 1 0 3404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1644511149
transform 1 0 2208 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1644511149
transform 1 0 2208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _317_
timestamp 1644511149
transform 1 0 3404 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 3680 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1644511149
transform 1 0 2208 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1644511149
transform 1 0 2208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1644511149
transform 1 0 3496 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1644511149
transform 1 0 3956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _323_
timestamp 1644511149
transform 1 0 2392 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1644511149
transform 1 0 2300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _325_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _328_
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1644511149
transform 1 0 4508 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1644511149
transform 1 0 4784 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1644511149
transform 1 0 2392 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1644511149
transform 1 0 2208 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _335_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5612 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _337_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _338_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _340_
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1644511149
transform 1 0 16376 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1644511149
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1644511149
transform 1 0 12788 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1644511149
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1644511149
transform 1 0 15364 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1644511149
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _349_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _350_
timestamp 1644511149
transform 1 0 4508 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _351_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _353_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _355_
timestamp 1644511149
transform 1 0 7544 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _356_
timestamp 1644511149
transform 1 0 4968 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _357_
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _358_
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _359_
timestamp 1644511149
transform 1 0 4692 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _360_
timestamp 1644511149
transform 1 0 4232 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _361_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _363_
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _365_
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1644511149
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1644511149
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _368_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _369_
timestamp 1644511149
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _370_
timestamp 1644511149
transform 1 0 8004 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _371_
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _372_
timestamp 1644511149
transform 1 0 8464 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _374_
timestamp 1644511149
transform 1 0 8464 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _376_
timestamp 1644511149
transform 1 0 9752 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _378_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _379_
timestamp 1644511149
transform 1 0 10120 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _380_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _381_
timestamp 1644511149
transform 1 0 10028 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _382_
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _383_
timestamp 1644511149
transform 1 0 13156 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_2  _384_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _385_
timestamp 1644511149
transform 1 0 15824 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _386_
timestamp 1644511149
transform 1 0 14628 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _387_
timestamp 1644511149
transform 1 0 10396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _388_
timestamp 1644511149
transform 1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _389_
timestamp 1644511149
transform 1 0 10672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _390_
timestamp 1644511149
transform 1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _391_
timestamp 1644511149
transform 1 0 9752 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _392_
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _393_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _394_
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _395_
timestamp 1644511149
transform 1 0 10488 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _396_
timestamp 1644511149
transform 1 0 10672 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _397_
timestamp 1644511149
transform 1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _398_
timestamp 1644511149
transform 1 0 10764 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _399_
timestamp 1644511149
transform 1 0 12512 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _400_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _401_
timestamp 1644511149
transform 1 0 10120 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _402_
timestamp 1644511149
transform 1 0 12696 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _403_
timestamp 1644511149
transform 1 0 10120 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _404_
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _405_
timestamp 1644511149
transform 1 0 12604 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _406_
timestamp 1644511149
transform 1 0 14444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _407_
timestamp 1644511149
transform 1 0 12052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _408_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _409_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _410_
timestamp 1644511149
transform 1 0 16744 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _411_
timestamp 1644511149
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _412_
timestamp 1644511149
transform 1 0 13248 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _413_
timestamp 1644511149
transform 1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _414_
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _415_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _416_
timestamp 1644511149
transform 1 0 15272 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _417_
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _418_
timestamp 1644511149
transform 1 0 15272 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _419_
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _420_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _421_
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _422_
timestamp 1644511149
transform 1 0 17480 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _423_
timestamp 1644511149
transform 1 0 13892 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _424_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _425_
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _426_
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _427_
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _428_
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _429_
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _430_
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _431_
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _432_
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _433_
timestamp 1644511149
transform 1 0 18216 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _434_
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _435_
timestamp 1644511149
transform 1 0 17204 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _436_
timestamp 1644511149
transform 1 0 17204 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _437_
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _438_
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _439_
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _440_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _441_
timestamp 1644511149
transform 1 0 15272 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _442_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _443_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _444_
timestamp 1644511149
transform 1 0 14260 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _445_
timestamp 1644511149
transform 1 0 15364 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _446_
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _447_
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _448_
timestamp 1644511149
transform 1 0 17112 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _449_
timestamp 1644511149
transform 1 0 17572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _450_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1644511149
transform 1 0 11684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp 1644511149
transform 1 0 17020 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1644511149
transform 1 0 14536 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1644511149
transform 1 0 16836 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1644511149
transform 1 0 16652 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1644511149
transform 1 0 17204 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1644511149
transform 1 0 13432 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1644511149
transform 1 0 13524 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _465_
timestamp 1644511149
transform 1 0 15456 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _466_
timestamp 1644511149
transform 1 0 14352 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _467_
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _468_
timestamp 1644511149
transform 1 0 10948 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _469_
timestamp 1644511149
transform 1 0 9568 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _470_
timestamp 1644511149
transform 1 0 3956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _471_
timestamp 1644511149
transform 1 0 6164 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _472_
timestamp 1644511149
transform 1 0 6992 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _473_
timestamp 1644511149
transform 1 0 4048 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1644511149
transform 1 0 5888 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _475_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _476_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _477_
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _478_
timestamp 1644511149
transform 1 0 5244 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _479_
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _480_
timestamp 1644511149
transform 1 0 8740 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _481_
timestamp 1644511149
transform 1 0 12696 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1644511149
transform 1 0 6532 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1644511149
transform 1 0 2208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1644511149
transform 1 0 2392 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1644511149
transform 1 0 1840 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1644511149
transform 1 0 6256 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1644511149
transform 1 0 4416 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1644511149
transform 1 0 5428 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1644511149
transform 1 0 1840 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1644511149
transform 1 0 1932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1644511149
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1644511149
transform 1 0 4508 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1644511149
transform 1 0 1840 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1644511149
transform 1 0 4140 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1644511149
transform 1 0 1840 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1644511149
transform 1 0 3128 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1644511149
transform 1 0 2852 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1644511149
transform 1 0 4416 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1644511149
transform 1 0 1840 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1644511149
transform 1 0 6072 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1644511149
transform 1 0 6716 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _508_
timestamp 1644511149
transform 1 0 3772 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1644511149
transform 1 0 6532 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1644511149
transform 1 0 17480 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1644511149
transform 1 0 13064 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _513__157 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514__158
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _515__159
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _516__160
timestamp 1644511149
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _517__161
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _518__162
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _519__163
timestamp 1644511149
transform 1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _520__110
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _521__111
timestamp 1644511149
transform 1 0 26220 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _522__112
timestamp 1644511149
transform 1 0 41216 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _523__113
timestamp 1644511149
transform 1 0 48760 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _524__114
timestamp 1644511149
transform 1 0 56212 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _525__115
timestamp 1644511149
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _526__116
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _527__117
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _528__118
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _529__119
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _530__120
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _531__121
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _532__122
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _533__123
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _534__124
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _535__125
timestamp 1644511149
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _536__126
timestamp 1644511149
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _537__127
timestamp 1644511149
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _538__128
timestamp 1644511149
transform 1 0 15916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539__129
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _540__130
timestamp 1644511149
transform 1 0 20516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _541__131
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _542__132
timestamp 1644511149
transform 1 0 25392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _543__133
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _544__134
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _545__135
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _546__136
timestamp 1644511149
transform 1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _547__137
timestamp 1644511149
transform 1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _548__138
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _549__139
timestamp 1644511149
transform 1 0 35328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _550__140
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _551__141
timestamp 1644511149
transform 1 0 38548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _552__142
timestamp 1644511149
transform 1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _553__143
timestamp 1644511149
transform 1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _554__144
timestamp 1644511149
transform 1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _555__145
timestamp 1644511149
transform 1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _556__146
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _557__147
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _558__148
timestamp 1644511149
transform 1 0 48760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _559__149
timestamp 1644511149
transform 1 0 49956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _560__150
timestamp 1644511149
transform 1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _561__151
timestamp 1644511149
transform 1 0 52900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _562__152
timestamp 1644511149
transform 1 0 54372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _563__153
timestamp 1644511149
transform 1 0 56028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _564__154
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _565__155
timestamp 1644511149
transform 1 0 57960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _566__156
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1644511149
transform 1 0 33396 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform 1 0 34868 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform 1 0 36340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1644511149
transform 1 0 40664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1644511149
transform 1 0 45080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1644511149
transform 1 0 48024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1644511149
transform 1 0 50968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1644511149
transform 1 0 53912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1644511149
transform 1 0 56764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1644511149
transform 1 0 56856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1644511149
transform 1 0 57684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 26036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 2852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input55 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 11776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 2116 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 2852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 2852 0 1 3264
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3698 41200 3754 42000 6 flash_csb
port 0 nsew signal tristate
rlabel metal2 s 11150 41200 11206 42000 6 flash_io0_read
port 1 nsew signal input
rlabel metal2 s 18694 41200 18750 42000 6 flash_io0_we
port 2 nsew signal tristate
rlabel metal2 s 26146 41200 26202 42000 6 flash_io0_write
port 3 nsew signal tristate
rlabel metal2 s 33690 41200 33746 42000 6 flash_io1_read
port 4 nsew signal input
rlabel metal2 s 41142 41200 41198 42000 6 flash_io1_we
port 5 nsew signal tristate
rlabel metal2 s 48686 41200 48742 42000 6 flash_io1_write
port 6 nsew signal tristate
rlabel metal2 s 56138 41200 56194 42000 6 flash_sck
port 7 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 sram_addr0[0]
port 8 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 sram_addr0[1]
port 9 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 sram_addr0[2]
port 10 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 sram_addr0[3]
port 11 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 sram_addr0[4]
port 12 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 sram_addr0[5]
port 13 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 sram_addr0[6]
port 14 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 sram_addr0[7]
port 15 nsew signal tristate
rlabel metal2 s 24030 0 24086 800 6 sram_addr0[8]
port 16 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 sram_addr1[0]
port 17 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 sram_addr1[1]
port 18 nsew signal tristate
rlabel metal2 s 8942 0 8998 800 6 sram_addr1[2]
port 19 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 sram_addr1[3]
port 20 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 sram_addr1[4]
port 21 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 sram_addr1[5]
port 22 nsew signal tristate
rlabel metal2 s 19706 0 19762 800 6 sram_addr1[6]
port 23 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 sram_addr1[7]
port 24 nsew signal tristate
rlabel metal2 s 24582 0 24638 800 6 sram_addr1[8]
port 25 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 sram_clk0
port 26 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 sram_clk1
port 27 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 sram_csb0
port 28 nsew signal tristate
rlabel metal2 s 1582 0 1638 800 6 sram_csb1
port 29 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 sram_din0[0]
port 30 nsew signal tristate
rlabel metal2 s 27986 0 28042 800 6 sram_din0[10]
port 31 nsew signal tristate
rlabel metal2 s 29458 0 29514 800 6 sram_din0[11]
port 32 nsew signal tristate
rlabel metal2 s 30838 0 30894 800 6 sram_din0[12]
port 33 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 sram_din0[13]
port 34 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 sram_din0[14]
port 35 nsew signal tristate
rlabel metal2 s 35254 0 35310 800 6 sram_din0[15]
port 36 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 sram_din0[16]
port 37 nsew signal tristate
rlabel metal2 s 38198 0 38254 800 6 sram_din0[17]
port 38 nsew signal tristate
rlabel metal2 s 39670 0 39726 800 6 sram_din0[18]
port 39 nsew signal tristate
rlabel metal2 s 41142 0 41198 800 6 sram_din0[19]
port 40 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 sram_din0[1]
port 41 nsew signal tristate
rlabel metal2 s 42614 0 42670 800 6 sram_din0[20]
port 42 nsew signal tristate
rlabel metal2 s 44086 0 44142 800 6 sram_din0[21]
port 43 nsew signal tristate
rlabel metal2 s 45466 0 45522 800 6 sram_din0[22]
port 44 nsew signal tristate
rlabel metal2 s 46938 0 46994 800 6 sram_din0[23]
port 45 nsew signal tristate
rlabel metal2 s 48410 0 48466 800 6 sram_din0[24]
port 46 nsew signal tristate
rlabel metal2 s 49882 0 49938 800 6 sram_din0[25]
port 47 nsew signal tristate
rlabel metal2 s 51354 0 51410 800 6 sram_din0[26]
port 48 nsew signal tristate
rlabel metal2 s 52826 0 52882 800 6 sram_din0[27]
port 49 nsew signal tristate
rlabel metal2 s 54298 0 54354 800 6 sram_din0[28]
port 50 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 sram_din0[29]
port 51 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 sram_din0[2]
port 52 nsew signal tristate
rlabel metal2 s 57242 0 57298 800 6 sram_din0[30]
port 53 nsew signal tristate
rlabel metal2 s 58714 0 58770 800 6 sram_din0[31]
port 54 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 sram_din0[3]
port 55 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 sram_din0[4]
port 56 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 sram_din0[5]
port 57 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 sram_din0[6]
port 58 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 sram_din0[7]
port 59 nsew signal tristate
rlabel metal2 s 25042 0 25098 800 6 sram_din0[8]
port 60 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 sram_din0[9]
port 61 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 sram_dout0[0]
port 62 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 sram_dout0[10]
port 63 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[11]
port 64 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 sram_dout0[12]
port 65 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 sram_dout0[13]
port 66 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 sram_dout0[14]
port 67 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 sram_dout0[15]
port 68 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 sram_dout0[16]
port 69 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 sram_dout0[17]
port 70 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 sram_dout0[18]
port 71 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 sram_dout0[19]
port 72 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 sram_dout0[1]
port 73 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 sram_dout0[20]
port 74 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 sram_dout0[21]
port 75 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 sram_dout0[22]
port 76 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout0[23]
port 77 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 sram_dout0[24]
port 78 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 sram_dout0[25]
port 79 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 sram_dout0[26]
port 80 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 sram_dout0[27]
port 81 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout0[28]
port 82 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 sram_dout0[29]
port 83 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 sram_dout0[2]
port 84 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 sram_dout0[30]
port 85 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 sram_dout0[31]
port 86 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 sram_dout0[3]
port 87 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 sram_dout0[4]
port 88 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 sram_dout0[5]
port 89 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 sram_dout0[6]
port 90 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 sram_dout0[7]
port 91 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 sram_dout0[8]
port 92 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 sram_dout0[9]
port 93 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 sram_dout1[0]
port 94 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 sram_dout1[10]
port 95 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 sram_dout1[11]
port 96 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 sram_dout1[12]
port 97 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 sram_dout1[13]
port 98 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 sram_dout1[14]
port 99 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 sram_dout1[15]
port 100 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 sram_dout1[16]
port 101 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 sram_dout1[17]
port 102 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 sram_dout1[18]
port 103 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 sram_dout1[19]
port 104 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 sram_dout1[1]
port 105 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 sram_dout1[20]
port 106 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 sram_dout1[21]
port 107 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 sram_dout1[22]
port 108 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 sram_dout1[23]
port 109 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 sram_dout1[24]
port 110 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 sram_dout1[25]
port 111 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[26]
port 112 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 sram_dout1[27]
port 113 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 sram_dout1[28]
port 114 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 sram_dout1[29]
port 115 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 sram_dout1[2]
port 116 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 sram_dout1[30]
port 117 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 sram_dout1[31]
port 118 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 sram_dout1[3]
port 119 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 sram_dout1[4]
port 120 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 sram_dout1[5]
port 121 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 sram_dout1[6]
port 122 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 sram_dout1[7]
port 123 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout1[8]
port 124 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 sram_dout1[9]
port 125 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 sram_web0
port 126 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 sram_wmask0[0]
port 127 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 sram_wmask0[1]
port 128 nsew signal tristate
rlabel metal2 s 10874 0 10930 800 6 sram_wmask0[2]
port 129 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 sram_wmask0[3]
port 130 nsew signal tristate
rlabel metal4 s 4208 2128 4528 39760 6 vccd1
port 131 nsew power input
rlabel metal4 s 34928 2128 35248 39760 6 vccd1
port 131 nsew power input
rlabel metal4 s 19568 2128 19888 39760 6 vssd1
port 132 nsew ground input
rlabel metal4 s 50288 2128 50608 39760 6 vssd1
port 132 nsew ground input
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 133 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 wb_adr_i[0]
port 134 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wb_adr_i[10]
port 135 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[11]
port 136 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[12]
port 137 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[13]
port 138 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[14]
port 139 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wb_adr_i[15]
port 140 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 wb_adr_i[16]
port 141 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wb_adr_i[17]
port 142 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wb_adr_i[18]
port 143 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wb_adr_i[19]
port 144 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wb_adr_i[1]
port 145 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_adr_i[20]
port 146 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wb_adr_i[21]
port 147 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_adr_i[22]
port 148 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[23]
port 149 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wb_adr_i[2]
port 150 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 wb_adr_i[3]
port 151 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wb_adr_i[4]
port 152 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 wb_adr_i[5]
port 153 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 wb_adr_i[6]
port 154 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 wb_adr_i[7]
port 155 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 wb_adr_i[8]
port 156 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wb_adr_i[9]
port 157 nsew signal input
rlabel metal3 s 0 552 800 672 6 wb_clk_i
port 158 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wb_cyc_i
port 159 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 wb_data_i[0]
port 160 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wb_data_i[10]
port 161 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[11]
port 162 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[12]
port 163 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[13]
port 164 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[14]
port 165 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wb_data_i[15]
port 166 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_data_i[16]
port 167 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wb_data_i[17]
port 168 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wb_data_i[18]
port 169 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wb_data_i[19]
port 170 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wb_data_i[1]
port 171 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wb_data_i[20]
port 172 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wb_data_i[21]
port 173 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 wb_data_i[22]
port 174 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_data_i[23]
port 175 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wb_data_i[24]
port 176 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 wb_data_i[25]
port 177 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 wb_data_i[26]
port 178 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 wb_data_i[27]
port 179 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 wb_data_i[28]
port 180 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 wb_data_i[29]
port 181 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 wb_data_i[2]
port 182 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 wb_data_i[30]
port 183 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 wb_data_i[31]
port 184 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 wb_data_i[3]
port 185 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wb_data_i[4]
port 186 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_data_i[5]
port 187 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wb_data_i[6]
port 188 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wb_data_i[7]
port 189 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wb_data_i[8]
port 190 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wb_data_i[9]
port 191 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 wb_data_o[0]
port 192 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 wb_data_o[10]
port 193 nsew signal tristate
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[11]
port 194 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[12]
port 195 nsew signal tristate
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[13]
port 196 nsew signal tristate
rlabel metal3 s 0 23672 800 23792 6 wb_data_o[14]
port 197 nsew signal tristate
rlabel metal3 s 0 24896 800 25016 6 wb_data_o[15]
port 198 nsew signal tristate
rlabel metal3 s 0 26120 800 26240 6 wb_data_o[16]
port 199 nsew signal tristate
rlabel metal3 s 0 27344 800 27464 6 wb_data_o[17]
port 200 nsew signal tristate
rlabel metal3 s 0 28704 800 28824 6 wb_data_o[18]
port 201 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 wb_data_o[19]
port 202 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 wb_data_o[1]
port 203 nsew signal tristate
rlabel metal3 s 0 31152 800 31272 6 wb_data_o[20]
port 204 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[21]
port 205 nsew signal tristate
rlabel metal3 s 0 33736 800 33856 6 wb_data_o[22]
port 206 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wb_data_o[23]
port 207 nsew signal tristate
rlabel metal3 s 0 35776 800 35896 6 wb_data_o[24]
port 208 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 wb_data_o[25]
port 209 nsew signal tristate
rlabel metal3 s 0 37544 800 37664 6 wb_data_o[26]
port 210 nsew signal tristate
rlabel metal3 s 0 38360 800 38480 6 wb_data_o[27]
port 211 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wb_data_o[28]
port 212 nsew signal tristate
rlabel metal3 s 0 39992 800 40112 6 wb_data_o[29]
port 213 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 wb_data_o[2]
port 214 nsew signal tristate
rlabel metal3 s 0 40808 800 40928 6 wb_data_o[30]
port 215 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 wb_data_o[31]
port 216 nsew signal tristate
rlabel metal3 s 0 9256 800 9376 6 wb_data_o[3]
port 217 nsew signal tristate
rlabel metal3 s 0 11024 800 11144 6 wb_data_o[4]
port 218 nsew signal tristate
rlabel metal3 s 0 12248 800 12368 6 wb_data_o[5]
port 219 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 wb_data_o[6]
port 220 nsew signal tristate
rlabel metal3 s 0 14832 800 14952 6 wb_data_o[7]
port 221 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 wb_data_o[8]
port 222 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 wb_data_o[9]
port 223 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wb_error_o
port 224 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 wb_rst_i
port 225 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wb_sel_i[0]
port 226 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wb_sel_i[1]
port 227 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 wb_sel_i[2]
port 228 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wb_sel_i[3]
port 229 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wb_stall_o
port 230 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 wb_stb_i
port 231 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 wb_we_i
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 42000
<< end >>
