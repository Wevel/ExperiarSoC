* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

.subckt CaravelHost caravel_irq[0] caravel_irq[1] caravel_irq[2] caravel_irq[3] caravel_uart_rx
+ caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0] caravel_wb_adr_o[10] caravel_wb_adr_o[11]
+ caravel_wb_adr_o[12] caravel_wb_adr_o[13] caravel_wb_adr_o[14] caravel_wb_adr_o[15]
+ caravel_wb_adr_o[16] caravel_wb_adr_o[17] caravel_wb_adr_o[18] caravel_wb_adr_o[19]
+ caravel_wb_adr_o[1] caravel_wb_adr_o[20] caravel_wb_adr_o[21] caravel_wb_adr_o[22]
+ caravel_wb_adr_o[23] caravel_wb_adr_o[24] caravel_wb_adr_o[25] caravel_wb_adr_o[26]
+ caravel_wb_adr_o[27] caravel_wb_adr_o[2] caravel_wb_adr_o[3] caravel_wb_adr_o[4]
+ caravel_wb_adr_o[5] caravel_wb_adr_o[6] caravel_wb_adr_o[7] caravel_wb_adr_o[8]
+ caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0] caravel_wb_data_i[10]
+ caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13] caravel_wb_data_i[14]
+ caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17] caravel_wb_data_i[18]
+ caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20] caravel_wb_data_i[21]
+ caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24] caravel_wb_data_i[25]
+ caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28] caravel_wb_data_i[29]
+ caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31] caravel_wb_data_i[3]
+ caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6] caravel_wb_data_i[7]
+ caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0] caravel_wb_data_o[10]
+ caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13] caravel_wb_data_o[14]
+ caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17] caravel_wb_data_o[18]
+ caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20] caravel_wb_data_o[21]
+ caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24] caravel_wb_data_o[25]
+ caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28] caravel_wb_data_o[29]
+ caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31] caravel_wb_data_o[3]
+ caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6] caravel_wb_data_o[7]
+ caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i caravel_wb_sel_o[0]
+ caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3] caravel_wb_stall_i caravel_wb_stb_o
+ caravel_wb_we_o core0Index[0] core0Index[1] core0Index[2] core0Index[3] core0Index[4]
+ core0Index[5] core0Index[6] core0Index[7] core1Index[0] core1Index[1] core1Index[2]
+ core1Index[3] core1Index[4] core1Index[5] core1Index[6] core1Index[7] manufacturerID[0]
+ manufacturerID[10] manufacturerID[1] manufacturerID[2] manufacturerID[3] manufacturerID[4]
+ manufacturerID[5] manufacturerID[6] manufacturerID[7] manufacturerID[8] manufacturerID[9]
+ partID[0] partID[10] partID[11] partID[12] partID[13] partID[14] partID[15] partID[1]
+ partID[2] partID[3] partID[4] partID[5] partID[6] partID[7] partID[8] partID[9]
+ vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12]
+ wbs_data_i[13] wbs_data_i[14] wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18]
+ wbs_data_i[19] wbs_data_i[1] wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23]
+ wbs_data_i[24] wbs_data_i[25] wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29]
+ wbs_data_i[2] wbs_data_i[30] wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5]
+ wbs_data_i[6] wbs_data_i[7] wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10]
+ wbs_data_o[11] wbs_data_o[12] wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16]
+ wbs_data_o[17] wbs_data_o[18] wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21]
+ wbs_data_o[22] wbs_data_o[23] wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27]
+ wbs_data_o[28] wbs_data_o[29] wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3]
+ wbs_data_o[4] wbs_data_o[5] wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7963_ _8570_/CLK _7963_/D vssd1 vssd1 vccd1 vccd1 _7963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7894_ _8436_/CLK _7894_/D vssd1 vssd1 vccd1 vccd1 _7894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6845_ _7808_/A _7548_/B vssd1 vssd1 vccd1 vccd1 _7586_/A sky130_fd_sc_hd__xor2_1
X_3988_ _3959_/X _8584_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__mux2_1
X_5727_ _5727_/A vssd1 vssd1 vccd1 vccd1 _8020_/D sky130_fd_sc_hd__clkbuf_1
X_8515_ _8515_/CLK _8515_/D vssd1 vssd1 vccd1 vccd1 _8515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7481__151 _7483__153/A vssd1 vssd1 vccd1 vccd1 _8490_/CLK sky130_fd_sc_hd__inv_2
X_8446_ _8604_/CLK _8446_/D vssd1 vssd1 vccd1 vccd1 _8446_/Q sky130_fd_sc_hd__dfxtp_1
X_5658_ _5658_/A vssd1 vssd1 vccd1 vccd1 _8058_/D sky130_fd_sc_hd__clkbuf_1
X_8377_ _8377_/CLK _8377_/D vssd1 vssd1 vccd1 vccd1 _8377_/Q sky130_fd_sc_hd__dfxtp_1
X_5589_ _5424_/X _8105_/Q _5591_/S vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3456_ _7104_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3456_/X sky130_fd_sc_hd__clkbuf_16
X_4609_ _5826_/A _4646_/A vssd1 vssd1 vccd1 vccd1 _4625_/S sky130_fd_sc_hd__nor2_2
XFILLER_117_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7328_ _7588_/A _7394_/A _7394_/B vssd1 vssd1 vccd1 vccd1 _7328_/X sky130_fd_sc_hd__and3_1
XFILLER_117_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7259_ _8429_/Q vssd1 vssd1 vccd1 vccd1 _7282_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7178__60 _7178__60/A vssd1 vssd1 vccd1 vccd1 _8369_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6928__380 _6928__380/A vssd1 vssd1 vccd1 vccd1 _8176_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4960_ _4990_/B _4939_/X _4946_/X _4959_/X vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__a31o_1
X_4891_ _8281_/Q _4812_/X _4665_/X _8243_/Q vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__a22o_1
X_3911_ _7961_/Q _7962_/Q _6499_/A _6376_/B vssd1 vssd1 vccd1 vccd1 _7790_/B sky130_fd_sc_hd__or4_2
XFILLER_20_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6561_ _6561_/A vssd1 vssd1 vccd1 vccd1 _7981_/D sky130_fd_sc_hd__clkbuf_1
X_5512_ _5512_/A vssd1 vssd1 vccd1 vccd1 _8140_/D sky130_fd_sc_hd__clkbuf_1
X_8300_ _8300_/CLK _8300_/D vssd1 vssd1 vccd1 vccd1 _8300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6760_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6492_ _8614_/Q _6494_/B _6492_/C vssd1 vssd1 vccd1 vccd1 _6492_/X sky130_fd_sc_hd__and3_1
X_8231_ _8231_/CLK _8231_/D vssd1 vssd1 vccd1 vccd1 _8231_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3310_ _6767_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3310_/X sky130_fd_sc_hd__clkbuf_16
X_5443_ _5420_/X _8174_/Q _5447_/S vssd1 vssd1 vccd1 vccd1 _5444_/A sky130_fd_sc_hd__mux2_1
X_8162_ _8162_/CLK _8162_/D vssd1 vssd1 vccd1 vccd1 _8162_/Q sky130_fd_sc_hd__dfxtp_1
X_5374_ _5377_/A vssd1 vssd1 vccd1 vccd1 _5374_/X sky130_fd_sc_hd__clkbuf_2
X_4325_ _4325_/A vssd1 vssd1 vccd1 vccd1 _8404_/D sky130_fd_sc_hd__clkbuf_1
X_8680__245 vssd1 vssd1 vccd1 vccd1 _8680__245/HI partID[13] sky130_fd_sc_hd__conb_1
XFILLER_99_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8093_ _8617_/CLK _8093_/D vssd1 vssd1 vccd1 vccd1 _8093_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4256_ _4256_/A vssd1 vssd1 vccd1 vccd1 _8462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7120__514 _7121__515/A vssd1 vssd1 vccd1 vccd1 _8323_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4187_ _4981_/A _4965_/A vssd1 vssd1 vccd1 vccd1 _4970_/C sky130_fd_sc_hd__nand2_1
X_7077__479 _7078__480/A vssd1 vssd1 vccd1 vccd1 _8288_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7946_ _8633_/CLK _7946_/D vssd1 vssd1 vccd1 vccd1 _7946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7877_ _8622_/CLK _7877_/D vssd1 vssd1 vccd1 vccd1 _7877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6828_ _8554_/Q _8553_/Q _8552_/Q _8551_/Q vssd1 vssd1 vccd1 vccd1 _6843_/A sky130_fd_sc_hd__and4_1
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8429_ _8440_/CLK _8429_/D vssd1 vssd1 vccd1 vccd1 _8429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3439_ _7020_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3439_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6327__200 _6327__200/A vssd1 vssd1 vccd1 vccd1 _7912_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7488__157 _7488__157/A vssd1 vssd1 vccd1 vccd1 _8496_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8664__229 vssd1 vssd1 vccd1 vccd1 _8664__229/HI manufacturerID[1] sky130_fd_sc_hd__conb_1
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4110_ _8576_/Q vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5090_ _5221_/A _5222_/B _8198_/Q vssd1 vssd1 vccd1 vccd1 _5103_/B sky130_fd_sc_hd__a21oi_2
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4041_ _4041_/A vssd1 vssd1 vccd1 vccd1 _8527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5992_ _5992_/A vssd1 vssd1 vccd1 vccd1 _5992_/X sky130_fd_sc_hd__clkbuf_1
X_7800_ _7806_/A vssd1 vssd1 vccd1 vccd1 _7800_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7539__24 _7540__25/A vssd1 vssd1 vccd1 vccd1 _8538_/CLK sky130_fd_sc_hd__inv_2
X_4943_ _4849_/A _8112_/Q _8064_/Q _4847_/A vssd1 vssd1 vccd1 vccd1 _4943_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7662_ _7661_/X _7662_/B vssd1 vssd1 vccd1 vccd1 _7663_/A sky130_fd_sc_hd__and2b_1
X_6613_ _6619_/A vssd1 vssd1 vccd1 vccd1 _6613_/X sky130_fd_sc_hd__buf_1
X_4874_ _4874_/A vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__buf_2
X_7593_ _7593_/A _7593_/B _7593_/C _7593_/D vssd1 vssd1 vccd1 vccd1 _7688_/B sky130_fd_sc_hd__and4_2
X_6544_ _8091_/Q _7976_/Q _6548_/S vssd1 vssd1 vccd1 vccd1 _6545_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7172__55 _7172__55/A vssd1 vssd1 vccd1 vccd1 _8364_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3256_ clkbuf_0__3256_/X vssd1 vssd1 vccd1 vccd1 _6626__271/A sky130_fd_sc_hd__clkbuf_4
X_6475_ _8619_/Q vssd1 vssd1 vccd1 vccd1 _7588_/A sky130_fd_sc_hd__clkbuf_4
X_5426_ _5426_/A vssd1 vssd1 vccd1 vccd1 _8181_/D sky130_fd_sc_hd__clkbuf_1
X_8214_ _8214_/CLK _8214_/D vssd1 vssd1 vccd1 vccd1 _8214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5357_ _5305_/A _5355_/X _5356_/X _5189_/A vssd1 vssd1 vccd1 vccd1 _5357_/X sky130_fd_sc_hd__o211a_1
X_8145_ _8633_/CLK _8145_/D vssd1 vssd1 vccd1 vccd1 _8145_/Q sky130_fd_sc_hd__dfxtp_1
X_8076_ _8076_/CLK _8076_/D vssd1 vssd1 vccd1 vccd1 _8076_/Q sky130_fd_sc_hd__dfxtp_1
X_4308_ _8411_/Q _4226_/X _4310_/S vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_4 _4197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5288_ _8527_/Q _5276_/X _5230_/B _8519_/Q vssd1 vssd1 vccd1 vccd1 _5288_/X sky130_fd_sc_hd__o22a_1
X_4239_ _8469_/Q _4238_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3472_ clkbuf_0__3472_/X vssd1 vssd1 vccd1 vccd1 _7188__68/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7929_ _7929_/CLK _7929_/D vssd1 vssd1 vccd1 vccd1 _7929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _4590_/A vssd1 vssd1 vccd1 vccd1 _8303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _6257_/X _8090_/Q _6253_/X _6255_/X _7879_/Q vssd1 vssd1 vccd1 vccd1 _7879_/D
+ sky130_fd_sc_hd__o32a_1
X_5211_ _5135_/X _5210_/X _5171_/X vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__a21o_1
X_6191_ _7958_/Q _6195_/C _6072_/A vssd1 vssd1 vccd1 vccd1 _6191_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5142_ _5139_/X _5141_/X _5142_/S vssd1 vssd1 vccd1 vccd1 _5142_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5073_ _5073_/A vssd1 vssd1 vccd1 vccd1 _8217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4024_ _4024_/A vssd1 vssd1 vccd1 vccd1 _8533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5975_ _5975_/A vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4926_ _4849_/A _8165_/Q _7993_/Q _4852_/A vssd1 vssd1 vccd1 vccd1 _4926_/X sky130_fd_sc_hd__a22o_1
X_7714_ _7714_/A _7716_/B _7714_/C vssd1 vssd1 vccd1 vccd1 _7715_/A sky130_fd_sc_hd__and3_1
XFILLER_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4857_ _4855_/X _8035_/Q _7848_/Q _4856_/X _4834_/X vssd1 vssd1 vccd1 vccd1 _4857_/X
+ sky130_fd_sc_hd__o221a_1
X_7645_ _7645_/A vssd1 vssd1 vccd1 vccd1 _8552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7576_ _7581_/A _7579_/A vssd1 vssd1 vccd1 vccd1 _7642_/A sky130_fd_sc_hd__nand2_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7050__460 _7050__460/A vssd1 vssd1 vccd1 vccd1 _8267_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3308_ clkbuf_0__3308_/X vssd1 vssd1 vccd1 vccd1 _6765__325/A sky130_fd_sc_hd__clkbuf_4
X_4788_ _8299_/Q _8283_/Q _8245_/Q _8315_/Q _4700_/X _4714_/X vssd1 vssd1 vccd1 vccd1
+ _4788_/X sky130_fd_sc_hd__mux4_1
X_6527_ _6527_/A vssd1 vssd1 vccd1 vccd1 _7968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6458_ _6501_/A _6396_/A _6436_/Y _6647_/A vssd1 vssd1 vccd1 vccd1 _6472_/A sky130_fd_sc_hd__a31o_2
X_5409_ _5408_/X _8185_/Q _5417_/S vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6389_ _6416_/A _6389_/B _6389_/C vssd1 vssd1 vccd1 vccd1 _6389_/Y sky130_fd_sc_hd__nor3_2
X_6764__324 _6765__325/A vssd1 vssd1 vccd1 vccd1 _8116_/CLK sky130_fd_sc_hd__inv_2
X_7439__118 _7441__120/A vssd1 vssd1 vccd1 vccd1 _8457_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8128_ _8128_/CLK _8128_/D vssd1 vssd1 vccd1 vccd1 _8128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8059_ _8059_/CLK _8059_/D vssd1 vssd1 vccd1 vccd1 _8059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3455_ clkbuf_0__3455_/X vssd1 vssd1 vccd1 vccd1 _7122_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7533__19 _7534__20/A vssd1 vssd1 vccd1 vccd1 _8533_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7342__109 _7342__109/A vssd1 vssd1 vccd1 vccd1 _8420_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6665__288 _6667__290/A vssd1 vssd1 vccd1 vccd1 _8056_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _8005_/Q _5627_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5761_/A sky130_fd_sc_hd__mux2_1
X_5691_ _5691_/A vssd1 vssd1 vccd1 vccd1 _8036_/D sky130_fd_sc_hd__clkbuf_1
X_4711_ _8302_/Q _8286_/Q _8248_/Q _8318_/Q _4710_/X _4702_/X vssd1 vssd1 vccd1 vccd1
+ _4711_/X sky130_fd_sc_hd__mux4_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4642_ _4475_/X _8280_/Q _4644_/S vssd1 vssd1 vccd1 vccd1 _4643_/A sky130_fd_sc_hd__mux2_1
X_7430_ _8451_/Q _7430_/B vssd1 vssd1 vccd1 vccd1 _7430_/X sky130_fd_sc_hd__or2_1
XFILLER_30_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _4573_/A _4646_/A vssd1 vssd1 vccd1 vccd1 _4589_/S sky130_fd_sc_hd__or2_2
X_7361_ _7361_/A _7361_/B vssd1 vssd1 vccd1 vccd1 _7361_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7292_ _8632_/Q _7292_/B vssd1 vssd1 vccd1 vccd1 _7292_/Y sky130_fd_sc_hd__xnor2_1
X_6312_ _8443_/Q _6312_/B vssd1 vssd1 vccd1 vccd1 _6312_/X sky130_fd_sc_hd__and2b_1
XFILLER_116_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6243_ _6240_/X _8080_/Q _6236_/X _6238_/X _7869_/Q vssd1 vssd1 vccd1 vccd1 _7869_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174_ _7886_/Q _6159_/X _6163_/X _6172_/X _6173_/X vssd1 vssd1 vccd1 vccd1 _6174_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5125_ _5144_/B _5125_/B vssd1 vssd1 vccd1 vccd1 _5204_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _5898_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5072_/S sky130_fd_sc_hd__or2_2
XFILLER_84_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4007_ _4646_/A _5539_/B vssd1 vssd1 vccd1 vccd1 _4023_/S sky130_fd_sc_hd__nor2_2
XFILLER_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _7818_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__or2_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7205__81 _7209__85/A vssd1 vssd1 vccd1 vccd1 _8390_/CLK sky130_fd_sc_hd__inv_2
X_4909_ _8017_/Q _4821_/X _4908_/X _4861_/X vssd1 vssd1 vccd1 vccd1 _4909_/X sky130_fd_sc_hd__o22a_1
X_5889_ _5889_/A vssd1 vssd1 vccd1 vccd1 _7857_/D sky130_fd_sc_hd__clkbuf_1
X_7628_ _7627_/X _7628_/B vssd1 vssd1 vccd1 vccd1 _7629_/A sky130_fd_sc_hd__and2b_1
XFILLER_119_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7559_ _7611_/A _7611_/B _8630_/Q vssd1 vssd1 vccd1 vccd1 _7562_/B sky130_fd_sc_hd__a21boi_1
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3438_ clkbuf_0__3438_/X vssd1 vssd1 vccd1 vccd1 _7019__435/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8561_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7001__421 _7002__422/A vssd1 vssd1 vccd1 vccd1 _8227_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6861_ _6861_/A _6891_/C _6852_/B vssd1 vssd1 vccd1 vccd1 _7566_/B sky130_fd_sc_hd__or3b_1
XFILLER_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5812_ _5598_/X _7934_/Q _5818_/S vssd1 vssd1 vccd1 vccd1 _5813_/A sky130_fd_sc_hd__mux2_1
X_8600_ _8600_/CLK _8600_/D vssd1 vssd1 vccd1 vccd1 _8600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5743_ _5743_/A vssd1 vssd1 vccd1 vccd1 _8013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8531_ _8531_/CLK _8531_/D vssd1 vssd1 vccd1 vccd1 _8531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8462_ _8462_/CLK _8462_/D vssd1 vssd1 vccd1 vccd1 _8462_/Q sky130_fd_sc_hd__dfxtp_1
X_5674_ _5607_/X _8043_/Q _5674_/S vssd1 vssd1 vccd1 vccd1 _5675_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3472_ _7185_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3472_/X sky130_fd_sc_hd__clkbuf_16
X_8393_ _8393_/CLK _8393_/D vssd1 vssd1 vccd1 vccd1 _8393_/Q sky130_fd_sc_hd__dfxtp_1
X_4625_ _8287_/Q _4504_/X _4625_/S vssd1 vssd1 vccd1 vccd1 _4626_/A sky130_fd_sc_hd__mux2_1
X_7413_ _7413_/A vssd1 vssd1 vccd1 vccd1 _7413_/X sky130_fd_sc_hd__clkbuf_2
X_7344_ _7436_/A vssd1 vssd1 vccd1 vccd1 _7344_/X sky130_fd_sc_hd__buf_1
X_4556_ _4571_/S vssd1 vssd1 vccd1 vccd1 _4565_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4487_ _8341_/Q _4486_/X _4496_/S vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__mux2_1
X_7275_ _8429_/Q _7266_/A _7274_/A vssd1 vssd1 vccd1 vccd1 _7369_/B sky130_fd_sc_hd__a21o_1
X_6226_ _7902_/Q _7901_/Q vssd1 vssd1 vccd1 vccd1 _6306_/B sky130_fd_sc_hd__or2b_4
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6173_/A vssd1 vssd1 vccd1 vccd1 _6157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5108_ _5358_/S vssd1 vssd1 vccd1 vccd1 _5345_/S sky130_fd_sc_hd__buf_4
XFILLER_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _7863_/Q _6088_/B vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__or2_1
X_5039_ _8232_/Q _4507_/X _5047_/S vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6215__188 _6216__189/A vssd1 vssd1 vccd1 vccd1 _7857_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6777__334 _6778__335/A vssd1 vssd1 vccd1 vccd1 _8126_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7070__474 _7071__475/A vssd1 vssd1 vccd1 vccd1 _8283_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ _4425_/S vssd1 vssd1 vccd1 vccd1 _4419_/S sky130_fd_sc_hd__clkbuf_2
X_5390_ _5112_/A _5385_/X _5389_/Y _5374_/X vssd1 vssd1 vccd1 vccd1 _8199_/D sky130_fd_sc_hd__o211a_1
X_4341_ _4111_/X _8397_/Q _4347_/S vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7060_ _7066_/A vssd1 vssd1 vccd1 vccd1 _7060_/X sky130_fd_sc_hd__buf_1
X_4272_ _8456_/Q _4203_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4273_/A sky130_fd_sc_hd__mux2_1
X_6011_ _6011_/A vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7962_ _8570_/CLK _7962_/D vssd1 vssd1 vccd1 vccd1 _7962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7893_ _8436_/CLK _7893_/D vssd1 vssd1 vccd1 vccd1 _7893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6844_ _6838_/Y _7555_/B _6900_/B vssd1 vssd1 vccd1 vccd1 _7548_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3987_ _3987_/A vssd1 vssd1 vccd1 vccd1 _8585_/D sky130_fd_sc_hd__clkbuf_1
X_5726_ _8020_/Q _5630_/X _5728_/S vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__mux2_1
X_8514_ _8514_/CLK _8514_/D vssd1 vssd1 vccd1 vccd1 _8514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8445_ _8604_/CLK _8445_/D vssd1 vssd1 vccd1 vccd1 _8445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5657_ _5610_/X _8058_/Q _5661_/S vssd1 vssd1 vccd1 vccd1 _5658_/A sky130_fd_sc_hd__mux2_1
X_8376_ _8376_/CLK _8376_/D vssd1 vssd1 vccd1 vccd1 _8376_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3455_ _7103_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3455_/X sky130_fd_sc_hd__clkbuf_16
X_5588_ _5588_/A vssd1 vssd1 vccd1 vccd1 _8106_/D sky130_fd_sc_hd__clkbuf_1
X_4608_ _4608_/A vssd1 vssd1 vccd1 vccd1 _8295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4539_ _4539_/A vssd1 vssd1 vccd1 vccd1 _8325_/D sky130_fd_sc_hd__clkbuf_1
X_7327_ _7327_/A _7327_/B _7327_/C _7327_/D vssd1 vssd1 vccd1 vccd1 _7334_/C sky130_fd_sc_hd__and4_1
X_7258_ _8430_/Q vssd1 vssd1 vccd1 vccd1 _7274_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7732__33 _7732__33/A vssd1 vssd1 vccd1 vccd1 _8584_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3410_ clkbuf_0__3410_/X vssd1 vssd1 vccd1 vccd1 _6920__374/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4890_ _4827_/X _4888_/X _4889_/X vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__o21a_1
X_3910_ _7963_/Q _7964_/Q _7965_/Q _7966_/Q vssd1 vssd1 vccd1 vccd1 _6376_/B sky130_fd_sc_hd__or4_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6560_ _7836_/A _6560_/B _6563_/C vssd1 vssd1 vccd1 vccd1 _6561_/A sky130_fd_sc_hd__and3_1
X_5511_ _8140_/Q _4492_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5512_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6797_/A sky130_fd_sc_hd__clkbuf_4
X_6491_ _7954_/Q _6483_/X _6474_/X _6490_/X _6472_/A vssd1 vssd1 vccd1 vccd1 _7954_/D
+ sky130_fd_sc_hd__a221o_1
X_8230_ _8230_/CLK _8230_/D vssd1 vssd1 vccd1 vccd1 _8230_/Q sky130_fd_sc_hd__dfxtp_1
X_5442_ _5442_/A vssd1 vssd1 vccd1 vccd1 _8175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8161_ _8161_/CLK _8161_/D vssd1 vssd1 vccd1 vccd1 _8161_/Q sky130_fd_sc_hd__dfxtp_1
X_5373_ _5373_/A _5377_/B vssd1 vssd1 vccd1 vccd1 _5373_/Y sky130_fd_sc_hd__nand2_1
X_4324_ _8404_/Q _4223_/X _4328_/S vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8092_ _8617_/CLK _8092_/D vssd1 vssd1 vccd1 vccd1 _8092_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _8462_/Q _4235_/X _4257_/S vssd1 vssd1 vccd1 vccd1 _4256_/A sky130_fd_sc_hd__mux2_1
X_4186_ _8269_/Q _7753_/B vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__and2_1
XFILLER_103_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6645__286 _6646__287/A vssd1 vssd1 vccd1 vccd1 _8046_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7945_ _8623_/CLK _7945_/D vssd1 vssd1 vccd1 vccd1 _7945_/Q sky130_fd_sc_hd__dfxtp_1
X_7876_ _8630_/CLK _7876_/D vssd1 vssd1 vccd1 vccd1 _7876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6827_ _7683_/A vssd1 vssd1 vccd1 vccd1 _7662_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5709_ _5709_/A vssd1 vssd1 vccd1 vccd1 _8028_/D sky130_fd_sc_hd__clkbuf_1
X_8428_ _8441_/CLK _8428_/D vssd1 vssd1 vccd1 vccd1 _8428_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3438_ _7014_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3438_/X sky130_fd_sc_hd__clkbuf_16
X_8359_ _8359_/CLK _8359_/D vssd1 vssd1 vccd1 vccd1 _8359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6334__205 _6334__205/A vssd1 vssd1 vccd1 vccd1 _7917_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _3971_/X _8527_/Q _4044_/S vssd1 vssd1 vccd1 vccd1 _4041_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5991_ _5991_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5992_/A sky130_fd_sc_hd__or2_4
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942_ _4861_/X _4940_/X _4941_/X vssd1 vssd1 vccd1 vccd1 _4946_/B sky130_fd_sc_hd__o21a_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7661_ _6835_/A _7642_/A _7647_/X _6846_/B vssd1 vssd1 vccd1 vccd1 _7661_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4873_ _4469_/X _4669_/X _4872_/X _4744_/X vssd1 vssd1 vccd1 vccd1 _8264_/D sky130_fd_sc_hd__o211a_1
X_7592_ _7587_/Y _7588_/X _7589_/Y _7590_/X _7591_/X vssd1 vssd1 vccd1 vccd1 _7593_/D
+ sky130_fd_sc_hd__o2111a_1
X_6543_ _6543_/A vssd1 vssd1 vccd1 vccd1 _7975_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3255_ clkbuf_0__3255_/X vssd1 vssd1 vccd1 vccd1 _6624__270/A sky130_fd_sc_hd__clkbuf_4
X_6474_ _6474_/A vssd1 vssd1 vccd1 vccd1 _6474_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5425_ _5424_/X _8181_/Q _5429_/S vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__mux2_1
X_8213_ _8213_/CLK _8213_/D vssd1 vssd1 vccd1 vccd1 _8213_/Q sky130_fd_sc_hd__dfxtp_1
X_7083__484 _7083__484/A vssd1 vssd1 vccd1 vccd1 _8293_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5356_ _8578_/Q _5220_/X _5238_/X _8594_/Q vssd1 vssd1 vccd1 vccd1 _5356_/X sky130_fd_sc_hd__o22a_1
X_8144_ _8610_/CLK _8144_/D vssd1 vssd1 vccd1 vccd1 _8144_/Q sky130_fd_sc_hd__dfxtp_1
X_4307_ _4307_/A vssd1 vssd1 vccd1 vccd1 _8412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8075_ _8075_/CLK _8075_/D vssd1 vssd1 vccd1 vccd1 _8075_/Q sky130_fd_sc_hd__dfxtp_1
X_5287_ _7914_/Q _8511_/Q _5345_/S vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_5 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3471_ clkbuf_0__3471_/X vssd1 vssd1 vccd1 vccd1 _7184__65/A sky130_fd_sc_hd__clkbuf_4
X_4238_ _8570_/Q vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__clkbuf_4
X_7026_ _7032_/A vssd1 vssd1 vccd1 vccd1 _7026_/X sky130_fd_sc_hd__buf_1
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _4259_/A _4852_/A _4172_/A vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__or3_1
XFILLER_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7928_ _7928_/CLK _7928_/D vssd1 vssd1 vccd1 vccd1 _7928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7859_ _7859_/CLK _7859_/D vssd1 vssd1 vccd1 vccd1 _7859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6587__240 _6587__240/A vssd1 vssd1 vccd1 vccd1 _8000_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494__162 _7496__164/A vssd1 vssd1 vccd1 vccd1 _8501_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5210_ _8291_/Q _8275_/Q _8537_/Q _8307_/Q _5341_/S _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5210_/X sky130_fd_sc_hd__mux4_2
X_6190_ input35/X input2/X _6172_/B vssd1 vssd1 vccd1 vccd1 _6190_/X sky130_fd_sc_hd__o21a_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5141_ _8508_/Q _8406_/Q _8143_/Q _8358_/Q _5123_/A _5140_/X vssd1 vssd1 vccd1 vccd1
+ _5141_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5072_ _4478_/X _8217_/Q _5072_/S vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4023_ _8533_/Q _3949_/X _4023_/S vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5974_ _7796_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__or2_1
XFILLER_80_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7713_ _7713_/A vssd1 vssd1 vccd1 vccd1 _8572_/D sky130_fd_sc_hd__clkbuf_1
X_4925_ _4831_/X _7985_/Q _4833_/X _8218_/Q _4758_/A vssd1 vssd1 vccd1 vccd1 _4925_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4856_ _4856_/A vssd1 vssd1 vccd1 vccd1 _4856_/X sky130_fd_sc_hd__clkbuf_2
X_7644_ _7643_/X _7649_/B vssd1 vssd1 vccd1 vccd1 _7645_/A sky130_fd_sc_hd__and2b_1
X_7575_ _7575_/A input1/X vssd1 vssd1 vccd1 vccd1 _7575_/X sky130_fd_sc_hd__or2_1
XFILLER_119_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4787_ _8457_/Q _8347_/Q _8060_/Q _8481_/Q _4710_/X _4694_/X vssd1 vssd1 vccd1 vccd1
+ _4787_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1_0__3307_ clkbuf_0__3307_/X vssd1 vssd1 vccd1 vccd1 _6758__319/A sky130_fd_sc_hd__clkbuf_4
X_6526_ _6034_/A _7968_/Q _6526_/S vssd1 vssd1 vccd1 vccd1 _6527_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6457_ _7814_/A _6471_/B _6469_/C vssd1 vssd1 vccd1 vccd1 _6457_/X sky130_fd_sc_hd__and3_1
X_5408_ _5601_/A vssd1 vssd1 vccd1 vccd1 _5408_/X sky130_fd_sc_hd__buf_2
X_6388_ _6436_/B _6383_/Y _6385_/X _6386_/Y _6387_/X vssd1 vssd1 vccd1 vccd1 _6389_/C
+ sky130_fd_sc_hd__o221a_1
X_8127_ _8127_/CLK _8127_/D vssd1 vssd1 vccd1 vccd1 _8127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5339_ _8303_/Q _5271_/X _5257_/X _8287_/Q _5135_/A vssd1 vssd1 vccd1 vccd1 _5339_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8058_ _8058_/CLK _8058_/D vssd1 vssd1 vccd1 vccd1 _8058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3454_ clkbuf_0__3454_/X vssd1 vssd1 vccd1 vccd1 _7099__497/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7133__525 _7133__525/A vssd1 vssd1 vccd1 vccd1 _8334_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6771__329 _6772__330/A vssd1 vssd1 vccd1 vccd1 _8121_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7027__441 _7028__442/A vssd1 vssd1 vccd1 vccd1 _8247_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6602__251 _6603__252/A vssd1 vssd1 vccd1 vccd1 _8011_/CLK sky130_fd_sc_hd__inv_2
X_4710_ _4710_/A vssd1 vssd1 vccd1 vccd1 _4710_/X sky130_fd_sc_hd__clkbuf_4
X_5690_ _8036_/Q _5630_/X _5692_/S vssd1 vssd1 vccd1 vccd1 _5691_/A sky130_fd_sc_hd__mux2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641_ _4641_/A vssd1 vssd1 vccd1 vccd1 _8281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4572_ _4572_/A vssd1 vssd1 vccd1 vccd1 _8311_/D sky130_fd_sc_hd__clkbuf_1
X_7360_ _7360_/A vssd1 vssd1 vccd1 vccd1 _7360_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7291_ _8426_/Q _7294_/B vssd1 vssd1 vccd1 vccd1 _7292_/B sky130_fd_sc_hd__xor2_1
X_6311_ _8444_/Q _8445_/Q _8446_/Q _8447_/Q _8441_/Q _8442_/Q vssd1 vssd1 vccd1 vccd1
+ _6312_/B sky130_fd_sc_hd__mux4_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6242_ _6240_/X _7900_/Q _6236_/X _6238_/X _7868_/Q vssd1 vssd1 vccd1 vccd1 _7868_/D
+ sky130_fd_sc_hd__o32a_1
X_6683__301 _6685__303/A vssd1 vssd1 vccd1 vccd1 _8069_/CLK sky130_fd_sc_hd__inv_2
X_6173_ _6173_/A vssd1 vssd1 vccd1 vccd1 _6173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _8524_/Q _8516_/Q _7919_/Q _8532_/Q _5122_/X _5123_/X vssd1 vssd1 vccd1 vccd1
+ _5124_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5055_ _5055_/A _5055_/B _5055_/C vssd1 vssd1 vccd1 vccd1 _5790_/B sky130_fd_sc_hd__nand3_4
X_4006_ _5844_/A vssd1 vssd1 vccd1 vccd1 _5539_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _5957_/A vssd1 vssd1 vccd1 vccd1 _5957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4908_ _4812_/A _8113_/Q _8065_/Q _4853_/A vssd1 vssd1 vccd1 vccd1 _4908_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5888_ _4200_/X _7857_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__mux2_1
X_7445__123 _7447__125/A vssd1 vssd1 vccd1 vccd1 _8462_/CLK sky130_fd_sc_hd__inv_2
X_7627_ _7624_/Y _7620_/X _7625_/X _7626_/Y vssd1 vssd1 vccd1 vccd1 _7627_/X sky130_fd_sc_hd__o22a_1
X_4839_ _8480_/Q _4680_/A _4838_/X _8456_/Q _4713_/A vssd1 vssd1 vccd1 vccd1 _4839_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7558_ _8632_/Q _7603_/A vssd1 vssd1 vccd1 vccd1 _7562_/A sky130_fd_sc_hd__xnor2_1
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6509_ _6017_/A _7790_/A _6515_/S vssd1 vssd1 vccd1 vccd1 _6510_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3437_ clkbuf_0__3437_/X vssd1 vssd1 vccd1 vccd1 _7013__430/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7739__39 _7740__40/A vssd1 vssd1 vccd1 vccd1 _8590_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6671__293 _6673__295/A vssd1 vssd1 vccd1 vccd1 _8061_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ _8546_/Q _7610_/A _7607_/A _6876_/A vssd1 vssd1 vccd1 vccd1 _6891_/C sky130_fd_sc_hd__nand4_2
XFILLER_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6791_ _6791_/A vssd1 vssd1 vccd1 vccd1 _6791_/X sky130_fd_sc_hd__buf_1
X_5811_ _5811_/A vssd1 vssd1 vccd1 vccd1 _7935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5742_ _8013_/Q _5627_/X _5746_/S vssd1 vssd1 vccd1 vccd1 _5743_/A sky130_fd_sc_hd__mux2_1
X_8530_ _8530_/CLK _8530_/D vssd1 vssd1 vccd1 vccd1 _8530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ _5673_/A vssd1 vssd1 vccd1 vccd1 _8044_/D sky130_fd_sc_hd__clkbuf_1
X_8461_ _8461_/CLK _8461_/D vssd1 vssd1 vccd1 vccd1 _8461_/Q sky130_fd_sc_hd__dfxtp_1
X_7509__175 _7509__175/A vssd1 vssd1 vccd1 vccd1 _8514_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3471_ _7179_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3471_/X sky130_fd_sc_hd__clkbuf_16
X_8392_ _8392_/CLK _8392_/D vssd1 vssd1 vccd1 vccd1 _8392_/Q sky130_fd_sc_hd__dfxtp_1
X_4624_ _4624_/A vssd1 vssd1 vccd1 vccd1 _8288_/D sky130_fd_sc_hd__clkbuf_1
X_7412_ _7412_/A vssd1 vssd1 vccd1 vccd1 _7413_/A sky130_fd_sc_hd__clkbuf_2
X_4555_ _5682_/A _5000_/A vssd1 vssd1 vccd1 vccd1 _4571_/S sky130_fd_sc_hd__nor2_2
XFILLER_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4486_ _8576_/Q vssd1 vssd1 vccd1 vccd1 _4486_/X sky130_fd_sc_hd__clkbuf_4
X_7274_ _7274_/A _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _7369_/A sky130_fd_sc_hd__nand3_1
X_6225_ _6236_/A vssd1 vssd1 vccd1 vccd1 _6225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _7881_/Q _6175_/A vssd1 vssd1 vccd1 vccd1 _6156_/X sky130_fd_sc_hd__or2_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5107_ _5258_/S vssd1 vssd1 vccd1 vccd1 _5358_/S sky130_fd_sc_hd__buf_2
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6609__257 _6611__259/A vssd1 vssd1 vccd1 vccd1 _8017_/CLK sky130_fd_sc_hd__inv_2
X_6087_ _7938_/Q input25/X _6188_/B vssd1 vssd1 vccd1 vccd1 _6087_/X sky130_fd_sc_hd__mux2_1
X_5038_ _5053_/S vssd1 vssd1 vccd1 vccd1 _5047_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_53_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7146__535 _7146__535/A vssd1 vssd1 vccd1 vccd1 _8344_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4340_ _4340_/A vssd1 vssd1 vccd1 vccd1 _8398_/D sky130_fd_sc_hd__clkbuf_1
X_4271_ _4271_/A vssd1 vssd1 vccd1 vccd1 _8457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _6010_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__and2_1
XFILLER_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7961_ _8570_/CLK _7961_/D vssd1 vssd1 vccd1 vccd1 _7961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6912_ _6912_/A vssd1 vssd1 vccd1 vccd1 _8163_/D sky130_fd_sc_hd__clkbuf_1
X_7892_ _8561_/CLK _7892_/D vssd1 vssd1 vccd1 vccd1 _7892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6843_ _6843_/A _6850_/A _6843_/C vssd1 vssd1 vccd1 vccd1 _6900_/B sky130_fd_sc_hd__and3_2
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6678__299 _6678__299/A vssd1 vssd1 vccd1 vccd1 _8067_/CLK sky130_fd_sc_hd__inv_2
X_3986_ _3952_/X _8585_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3987_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5725_ _5725_/A vssd1 vssd1 vccd1 vccd1 _8021_/D sky130_fd_sc_hd__clkbuf_1
X_8513_ _8513_/CLK _8513_/D vssd1 vssd1 vccd1 vccd1 _8513_/Q sky130_fd_sc_hd__dfxtp_1
X_5656_ _5656_/A vssd1 vssd1 vccd1 vccd1 _8059_/D sky130_fd_sc_hd__clkbuf_1
X_8444_ _8604_/CLK _8444_/D vssd1 vssd1 vccd1 vccd1 _8444_/Q sky130_fd_sc_hd__dfxtp_1
X_4607_ _4478_/X _8295_/Q _4607_/S vssd1 vssd1 vccd1 vccd1 _4608_/A sky130_fd_sc_hd__mux2_1
X_8375_ _8375_/CLK _8375_/D vssd1 vssd1 vccd1 vccd1 _8375_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3454_ _7097_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3454_/X sky130_fd_sc_hd__clkbuf_16
X_5587_ _5420_/X _8106_/Q _5591_/S vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4538_ _4432_/X _8325_/Q _4544_/S vssd1 vssd1 vccd1 vccd1 _4539_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7326_ _7811_/A _7268_/B _7323_/Y _7324_/X _7325_/Y vssd1 vssd1 vccd1 vccd1 _7327_/D
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7257_ _7308_/A _7308_/B vssd1 vssd1 vccd1 vccd1 _7324_/B sky130_fd_sc_hd__nand2_1
X_4469_ _8191_/Q vssd1 vssd1 vccd1 vccd1 _4469_/X sky130_fd_sc_hd__buf_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6139_ _6173_/A vssd1 vssd1 vccd1 vccd1 _6139_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6581__235 _6581__235/A vssd1 vssd1 vccd1 vccd1 _7995_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7458__133 _7458__133/A vssd1 vssd1 vccd1 vccd1 _8472_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _5510_/A vssd1 vssd1 vccd1 vccd1 _8141_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3271_ clkbuf_0__3271_/X vssd1 vssd1 vccd1 vccd1 _6679__300/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7184__65 _7184__65/A vssd1 vssd1 vccd1 vccd1 _8374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6490_ _8615_/Q _6490_/B _6492_/C vssd1 vssd1 vccd1 vccd1 _6490_/X sky130_fd_sc_hd__and3_1
X_5441_ _5416_/X _8175_/Q _5441_/S vssd1 vssd1 vccd1 vccd1 _5442_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8160_ _8160_/CLK _8160_/D vssd1 vssd1 vccd1 vccd1 _8160_/Q sky130_fd_sc_hd__dfxtp_1
X_5372_ _3877_/B _5377_/B _5371_/X _5303_/X vssd1 vssd1 vccd1 vccd1 _8205_/D sky130_fd_sc_hd__o211a_1
X_4323_ _4323_/A vssd1 vssd1 vccd1 vccd1 _8405_/D sky130_fd_sc_hd__clkbuf_1
X_8091_ _8091_/CLK _8091_/D vssd1 vssd1 vccd1 vccd1 _8091_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4254_ _4254_/A vssd1 vssd1 vccd1 vccd1 _8463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4185_ _4169_/X _4173_/X _4180_/Y _4184_/Y vssd1 vssd1 vccd1 vccd1 _7753_/B sky130_fd_sc_hd__a211o_2
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7944_ _8633_/CLK _7944_/D vssd1 vssd1 vccd1 vccd1 _7944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ _8622_/CLK _7875_/D vssd1 vssd1 vccd1 vccd1 _7875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6826_ _7600_/A vssd1 vssd1 vccd1 vccd1 _7683_/A sky130_fd_sc_hd__buf_2
XFILLER_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5708_ _5604_/X _8028_/Q _5710_/S vssd1 vssd1 vccd1 vccd1 _5709_/A sky130_fd_sc_hd__mux2_1
X_3969_ _3968_/X _8589_/Q _3969_/S vssd1 vssd1 vccd1 vccd1 _3970_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6688_ _6694_/A vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3469_ clkbuf_0__3469_/X vssd1 vssd1 vccd1 vccd1 _7172__55/A sky130_fd_sc_hd__clkbuf_4
X_8427_ _8441_/CLK _8427_/D vssd1 vssd1 vccd1 vccd1 _8427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5639_ _8189_/Q vssd1 vssd1 vccd1 vccd1 _5639_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8358_ _8358_/CLK _8358_/D vssd1 vssd1 vccd1 vccd1 _8358_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3437_ _7008_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3437_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_88_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7309_ _8435_/Q _7308_/A _7308_/B _7266_/C _8436_/Q vssd1 vssd1 vccd1 vccd1 _7310_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8289_ _8289_/CLK _8289_/D vssd1 vssd1 vccd1 vccd1 _8289_/Q sky130_fd_sc_hd__dfxtp_1
X_7021__436 _7023__438/A vssd1 vssd1 vccd1 vccd1 _8242_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _5990_/A vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4941_ _8417_/Q _4855_/A _8225_/Q _4865_/A _4724_/A vssd1 vssd1 vccd1 vccd1 _4941_/X
+ sky130_fd_sc_hd__o221a_1
X_7660_ _7660_/A vssd1 vssd1 vccd1 vccd1 _8556_/D sky130_fd_sc_hd__clkbuf_1
X_4872_ _4872_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4872_/X sky130_fd_sc_hd__or2_1
X_7591_ _6893_/Y _6894_/X _6881_/X vssd1 vssd1 vccd1 vccd1 _7591_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6542_ _8090_/Q _7975_/Q _6548_/S vssd1 vssd1 vccd1 vccd1 _6543_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_9_wb_clk_i _6197_/A vssd1 vssd1 vccd1 vccd1 _8052_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1_0__3254_ clkbuf_0__3254_/X vssd1 vssd1 vccd1 vccd1 _6616__263/A sky130_fd_sc_hd__clkbuf_4
X_6473_ _7949_/Q _6464_/X _6452_/X _6471_/X _6472_/X vssd1 vssd1 vccd1 vccd1 _7949_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5424_ _5613_/A vssd1 vssd1 vccd1 vccd1 _5424_/X sky130_fd_sc_hd__clkbuf_2
Xoutput200 _6187_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__buf_2
X_8212_ _8212_/CLK _8212_/D vssd1 vssd1 vccd1 vccd1 _8212_/Q sky130_fd_sc_hd__dfxtp_1
X_8143_ _8143_/CLK _8143_/D vssd1 vssd1 vccd1 vccd1 _8143_/Q sky130_fd_sc_hd__dfxtp_1
X_5355_ _8120_/Q _8147_/Q _5355_/S vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__mux2_1
X_4306_ _8412_/Q _4223_/X _4310_/S vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__mux2_1
X_8074_ _8074_/CLK _8074_/D vssd1 vssd1 vccd1 vccd1 _8074_/Q sky130_fd_sc_hd__dfxtp_1
X_5286_ _5351_/A _5286_/B _5286_/C vssd1 vssd1 vccd1 vccd1 _5286_/X sky130_fd_sc_hd__or3_1
XFILLER_59_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_6 _4209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4237_ _4237_/A vssd1 vssd1 vccd1 vccd1 _8470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3470_ clkbuf_0__3470_/X vssd1 vssd1 vccd1 vccd1 _7177__59/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4168_ _8256_/Q _8251_/Q vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__xor2_1
XFILLER_82_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4099_ _8502_/Q _3946_/X _4101_/S vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7927_ _7927_/CLK _7927_/D vssd1 vssd1 vccd1 vccd1 _7927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7858_ _7858_/CLK _7858_/D vssd1 vssd1 vccd1 vccd1 _7858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7789_ _8145_/Q vssd1 vssd1 vccd1 vccd1 _7791_/A sky130_fd_sc_hd__clkinv_2
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6999__420 _6999__420/A vssd1 vssd1 vccd1 vccd1 _8226_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6340__210 _6340__210/A vssd1 vssd1 vccd1 vccd1 _7922_/CLK sky130_fd_sc_hd__inv_2
X_8670__235 vssd1 vssd1 vccd1 vccd1 _8670__235/HI manufacturerID[7] sky130_fd_sc_hd__conb_1
XFILLER_42_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5140_ _5358_/S vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__buf_2
X_5071_ _5071_/A vssd1 vssd1 vccd1 vccd1 _8218_/D sky130_fd_sc_hd__clkbuf_1
X_4022_ _4022_/A vssd1 vssd1 vccd1 vccd1 _8534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5973_ _5995_/A vssd1 vssd1 vccd1 vccd1 _5982_/B sky130_fd_sc_hd__clkbuf_1
X_7217__91 _7219__93/A vssd1 vssd1 vccd1 vccd1 _8400_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924_ _4874_/X _8105_/Q _8001_/Q _4847_/X _4809_/A vssd1 vssd1 vccd1 vccd1 _4924_/X
+ sky130_fd_sc_hd__a221o_1
X_7712_ _7838_/A _7716_/B _7714_/C vssd1 vssd1 vccd1 vccd1 _7713_/A sky130_fd_sc_hd__and3_1
XFILLER_100_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4855_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4855_/X sky130_fd_sc_hd__clkbuf_2
X_7643_ _7641_/Y _7642_/X _7625_/X _7590_/B vssd1 vssd1 vccd1 vccd1 _7643_/X sky130_fd_sc_hd__o22a_1
X_7574_ _8541_/Q _8542_/Q vssd1 vssd1 vccd1 vccd1 _7681_/A sky130_fd_sc_hd__or2b_2
X_4786_ _4463_/X _4669_/X _4785_/X _4744_/X vssd1 vssd1 vccd1 vccd1 _8266_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6525_ _6525_/A vssd1 vssd1 vccd1 vccd1 _7967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6456_ _8145_/Q vssd1 vssd1 vccd1 vccd1 _6469_/C sky130_fd_sc_hd__clkbuf_1
X_5407_ _8193_/Q vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6387_ _6387_/A vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8126_ _8126_/CLK _8126_/D vssd1 vssd1 vccd1 vccd1 _8126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5338_ _8533_/Q _8271_/Q _5345_/S vssd1 vssd1 vccd1 vccd1 _5338_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8057_ _8057_/CLK _8057_/D vssd1 vssd1 vccd1 vccd1 _8057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7008_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7008_/X sky130_fd_sc_hd__buf_1
X_5269_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__buf_2
XFILLER_68_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3453_ clkbuf_0__3453_/X vssd1 vssd1 vccd1 vccd1 _7096__495/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8654__219 vssd1 vssd1 vccd1 vccd1 _8654__219/HI core0Index[6] sky130_fd_sc_hd__conb_1
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4472_/X _8281_/Q _4644_/S vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__mux2_1
X_4571_ _8311_/Q _4531_/X _4571_/S vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__mux2_1
X_6310_ _8448_/Q _8449_/Q _8450_/Q _8451_/Q _8441_/Q _8442_/Q vssd1 vssd1 vccd1 vccd1
+ _6310_/X sky130_fd_sc_hd__mux4_1
X_7290_ _8425_/Q vssd1 vssd1 vccd1 vccd1 _7294_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6241_ _6240_/X _7899_/Q _6236_/X _6238_/X _7867_/Q vssd1 vssd1 vccd1 vccd1 _7867_/D
+ sky130_fd_sc_hd__o32a_1
X_6172_ _6172_/A _6172_/B vssd1 vssd1 vccd1 vccd1 _6172_/X sky130_fd_sc_hd__and2_4
X_5123_ _5123_/A vssd1 vssd1 vccd1 vccd1 _5123_/X sky130_fd_sc_hd__buf_2
XFILLER_97_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5054_ _5054_/A vssd1 vssd1 vccd1 vccd1 _8225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4005_ _5150_/A _5376_/B vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__nand2_4
XFILLER_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5956_ _7723_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__or2_1
XFILLER_111_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5887_ _5887_/A vssd1 vssd1 vccd1 vccd1 _7858_/D sky130_fd_sc_hd__clkbuf_1
X_4907_ _4845_/X _4905_/X _4906_/X vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__o21a_1
X_4838_ _4865_/A vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__clkbuf_4
X_7626_ _7626_/A _7626_/B vssd1 vssd1 vccd1 vccd1 _7626_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4769_ _8300_/Q _8284_/Q _8246_/Q _8316_/Q _4700_/X _4714_/X vssd1 vssd1 vccd1 vccd1
+ _4769_/X sky130_fd_sc_hd__mux4_1
X_7557_ _7552_/X _7553_/Y _7554_/Y _7555_/Y _7556_/X vssd1 vssd1 vccd1 vccd1 _7557_/X
+ sky130_fd_sc_hd__o2111a_1
X_6508_ _6508_/A vssd1 vssd1 vccd1 vccd1 _7959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6439_ _6501_/A _6437_/X _6438_/X vssd1 vssd1 vccd1 vccd1 _7942_/D sky130_fd_sc_hd__a21o_1
X_8109_ _8109_/CLK _8109_/D vssd1 vssd1 vccd1 vccd1 _8109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6961__393 _6963__395/A vssd1 vssd1 vccd1 vccd1 _8197_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7452__128 _7453__129/A vssd1 vssd1 vccd1 vccd1 _8467_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3436_ clkbuf_0__3436_/X vssd1 vssd1 vccd1 vccd1 _7032_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7096__495 _7096__495/A vssd1 vssd1 vccd1 vccd1 _8304_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7211__86 _7214__89/A vssd1 vssd1 vccd1 vccd1 _8395_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7516__5 _7516__5/A vssd1 vssd1 vccd1 vccd1 _8519_/CLK sky130_fd_sc_hd__inv_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8610_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8676__241 vssd1 vssd1 vccd1 vccd1 _8676__241/HI partID[5] sky130_fd_sc_hd__conb_1
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5810_ _5593_/X _7935_/Q _5818_/S vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ _5741_/A vssd1 vssd1 vccd1 vccd1 _8014_/D sky130_fd_sc_hd__clkbuf_1
X_8460_ _8460_/CLK _8460_/D vssd1 vssd1 vccd1 vccd1 _8460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5672_ _5604_/X _8044_/Q _5674_/S vssd1 vssd1 vccd1 vccd1 _5673_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7411_ _7411_/A vssd1 vssd1 vccd1 vccd1 _7756_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__3470_ _7173_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3470_/X sky130_fd_sc_hd__clkbuf_16
X_8391_ _8391_/CLK _8391_/D vssd1 vssd1 vccd1 vccd1 _8391_/Q sky130_fd_sc_hd__dfxtp_1
X_4623_ _8288_/Q _4501_/X _4625_/S vssd1 vssd1 vccd1 vccd1 _4624_/A sky130_fd_sc_hd__mux2_1
X_4554_ _4508_/B _5055_/C _5055_/A vssd1 vssd1 vccd1 vccd1 _5000_/A sky130_fd_sc_hd__nand3b_4
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7273_ _7373_/A _7373_/B _7569_/A vssd1 vssd1 vccd1 vccd1 _7331_/A sky130_fd_sc_hd__a21o_1
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4485_ _4485_/A vssd1 vssd1 vccd1 vccd1 _8342_/D sky130_fd_sc_hd__clkbuf_1
X_6224_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__buf_4
XFILLER_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7956_/Q input15/X _6177_/A vssd1 vssd1 vccd1 vccd1 _6155_/X sky130_fd_sc_hd__mux2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5222_/B vssd1 vssd1 vccd1 vccd1 _5258_/S sky130_fd_sc_hd__clkbuf_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6073_/X _6084_/X _6085_/X _6082_/X vssd1 vssd1 vccd1 vccd1 _6086_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5862_/A _5594_/A vssd1 vssd1 vccd1 vccd1 _5053_/S sky130_fd_sc_hd__nor2_2
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6988_ _7000_/A vssd1 vssd1 vccd1 vccd1 _6988_/X sky130_fd_sc_hd__buf_1
X_5939_ _6008_/B vssd1 vssd1 vccd1 vccd1 _5949_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7744__43 _7746__45/A vssd1 vssd1 vccd1 vccd1 _8594_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8589_ _8589_/CLK _8589_/D vssd1 vssd1 vccd1 vccd1 _8589_/Q sky130_fd_sc_hd__dfxtp_1
X_7609_ _7607_/X _7608_/X _7601_/X vssd1 vssd1 vccd1 vccd1 _8544_/D sky130_fd_sc_hd__o21a_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput100 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _7818_/A sky130_fd_sc_hd__buf_4
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6968__399 _6968__399/A vssd1 vssd1 vccd1 vccd1 _8203_/CLK sky130_fd_sc_hd__inv_2
X_4270_ _8457_/Q _4200_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7960_ _8570_/CLK _7960_/D vssd1 vssd1 vccd1 vccd1 _7960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6911_ _7662_/B _6911_/B _7681_/B vssd1 vssd1 vccd1 vccd1 _6912_/A sky130_fd_sc_hd__and3_1
X_7891_ _8561_/CLK _7891_/D vssd1 vssd1 vccd1 vccd1 _7891_/Q sky130_fd_sc_hd__dfxtp_1
X_6842_ _8553_/Q _6886_/A _6842_/C _6886_/C vssd1 vssd1 vccd1 vccd1 _7555_/B sky130_fd_sc_hd__nand4_4
XFILLER_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6773_ _6785_/A vssd1 vssd1 vccd1 vccd1 _6773_/X sky130_fd_sc_hd__buf_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _4000_/S vssd1 vssd1 vccd1 vccd1 _3994_/S sky130_fd_sc_hd__clkbuf_2
X_5724_ _8021_/Q _5627_/X _5728_/S vssd1 vssd1 vccd1 vccd1 _5725_/A sky130_fd_sc_hd__mux2_1
X_8512_ _8512_/CLK _8512_/D vssd1 vssd1 vccd1 vccd1 _8512_/Q sky130_fd_sc_hd__dfxtp_1
X_5655_ _5607_/X _8059_/Q _5655_/S vssd1 vssd1 vccd1 vccd1 _5656_/A sky130_fd_sc_hd__mux2_1
X_8443_ _8452_/CLK _8443_/D vssd1 vssd1 vccd1 vccd1 _8443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8374_ _8374_/CLK _8374_/D vssd1 vssd1 vccd1 vccd1 _8374_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3453_ _7091_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3453_/X sky130_fd_sc_hd__clkbuf_16
X_4606_ _4606_/A vssd1 vssd1 vccd1 vccd1 _8296_/D sky130_fd_sc_hd__clkbuf_1
X_6615__262 _6616__263/A vssd1 vssd1 vccd1 vccd1 _8022_/CLK sky130_fd_sc_hd__inv_2
X_5586_ _5586_/A vssd1 vssd1 vccd1 vccd1 _8107_/D sky130_fd_sc_hd__clkbuf_1
X_7325_ _7324_/B _7324_/C _7324_/A vssd1 vssd1 vccd1 vccd1 _7325_/Y sky130_fd_sc_hd__a21oi_1
X_4537_ _4537_/A vssd1 vssd1 vccd1 vccd1 _8326_/D sky130_fd_sc_hd__clkbuf_1
X_4468_ _4468_/A vssd1 vssd1 vccd1 vccd1 _8347_/D sky130_fd_sc_hd__clkbuf_1
X_6318__192 _6321__195/A vssd1 vssd1 vccd1 vccd1 _7904_/CLK sky130_fd_sc_hd__inv_2
X_7256_ _7280_/C vssd1 vssd1 vccd1 vccd1 _7308_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4399_ _4119_/X _8371_/Q _4401_/S vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__mux2_1
X_6138_ _7876_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6138_/X sky130_fd_sc_hd__or2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6069_ _8099_/Q _6069_/B vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__and2_2
XFILLER_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6993__415 _6993__415/A vssd1 vssd1 vccd1 vccd1 _8221_/CLK sky130_fd_sc_hd__inv_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7152__540 _7152__540/A vssd1 vssd1 vccd1 vccd1 _8349_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7169__52 _7169__52/A vssd1 vssd1 vccd1 vccd1 _8361_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3270_ clkbuf_0__3270_/X vssd1 vssd1 vccd1 vccd1 _6673__295/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _5440_/A vssd1 vssd1 vccd1 vccd1 _8176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5371_ _4336_/B _5370_/A _5382_/B _4299_/A vssd1 vssd1 vccd1 vccd1 _5371_/X sky130_fd_sc_hd__a31o_1
X_4322_ _8405_/Q _4220_/X _4328_/S vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__mux2_1
X_7110_ _7122_/A vssd1 vssd1 vccd1 vccd1 _7110_/X sky130_fd_sc_hd__buf_1
X_8090_ _8091_/CLK _8090_/D vssd1 vssd1 vccd1 vccd1 _8090_/Q sky130_fd_sc_hd__dfxtp_4
X_4253_ _8463_/Q _4232_/X _4257_/S vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4184_ _4666_/D _4183_/X _4969_/B vssd1 vssd1 vccd1 vccd1 _4184_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7943_ _8610_/CLK _7943_/D vssd1 vssd1 vccd1 vccd1 _7943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7874_ _8623_/CLK _7874_/D vssd1 vssd1 vccd1 vccd1 _7874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6825_ _7842_/A _4164_/X _6280_/A vssd1 vssd1 vccd1 vccd1 _7600_/A sky130_fd_sc_hd__a21oi_4
XFILLER_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3968_ _8573_/Q vssd1 vssd1 vccd1 vccd1 _3968_/X sky130_fd_sc_hd__buf_2
X_5707_ _5707_/A vssd1 vssd1 vccd1 vccd1 _8029_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3468_ clkbuf_0__3468_/X vssd1 vssd1 vccd1 vccd1 _7191_/A sky130_fd_sc_hd__clkbuf_4
X_3899_ _3899_/A _3899_/B _3899_/C _3899_/D vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__or4_1
X_5638_ _5638_/A vssd1 vssd1 vccd1 vccd1 _8066_/D sky130_fd_sc_hd__clkbuf_1
X_8426_ _8441_/CLK _8426_/D vssd1 vssd1 vccd1 vccd1 _8426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8357_ _8357_/CLK _8357_/D vssd1 vssd1 vccd1 vccd1 _8357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5569_ _5420_/X _8114_/Q _5573_/S vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3436_ _7007_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3436_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7308_ _7308_/A _7308_/B _7308_/C vssd1 vssd1 vccd1 vccd1 _7310_/A sky130_fd_sc_hd__nand3_1
XFILLER_78_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8288_ _8288_/CLK _8288_/D vssd1 vssd1 vccd1 vccd1 _8288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7239_ _8428_/Q _8427_/Q _8426_/Q _8425_/Q vssd1 vssd1 vccd1 vccd1 _7260_/A sky130_fd_sc_hd__and4_1
X_6808__354 _6809__355/A vssd1 vssd1 vccd1 vccd1 _8149_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _4812_/A _8180_/Q _8072_/Q _4822_/A vssd1 vssd1 vccd1 vccd1 _4940_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4871_ _4672_/A _8264_/Q _4859_/X _4870_/X _4741_/A vssd1 vssd1 vccd1 vccd1 _4872_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7590_ _7590_/A _7590_/B vssd1 vssd1 vccd1 vccd1 _7590_/X sky130_fd_sc_hd__xor2_1
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6541_ _6541_/A vssd1 vssd1 vccd1 vccd1 _7974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3253_ clkbuf_0__3253_/X vssd1 vssd1 vccd1 vccd1 _6612__260/A sky130_fd_sc_hd__clkbuf_4
X_6472_ _6472_/A vssd1 vssd1 vccd1 vccd1 _6472_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput201 _6189_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__buf_2
X_8211_ _8211_/CLK _8211_/D vssd1 vssd1 vccd1 vccd1 _8211_/Q sky130_fd_sc_hd__dfxtp_1
X_5423_ _8189_/Q vssd1 vssd1 vccd1 vccd1 _5613_/A sky130_fd_sc_hd__clkbuf_2
X_8142_ _8142_/CLK _8142_/D vssd1 vssd1 vccd1 vccd1 _8142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5354_ _5305_/A _5352_/X _5353_/X vssd1 vssd1 vccd1 vccd1 _5354_/X sky130_fd_sc_hd__o21a_1
X_4305_ _4305_/A vssd1 vssd1 vccd1 vccd1 _8413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8073_ _8073_/CLK _8073_/D vssd1 vssd1 vccd1 vccd1 _8073_/Q sky130_fd_sc_hd__dfxtp_1
X_5285_ _8503_/Q _5238_/X _5142_/S _5284_/X vssd1 vssd1 vccd1 vccd1 _5286_/C sky130_fd_sc_hd__o211a_1
XFILLER_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_7 _4209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _8470_/Q _4235_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4237_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4167_ _4171_/B vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__buf_2
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4098_ _4098_/A vssd1 vssd1 vccd1 vccd1 _8503_/D sky130_fd_sc_hd__clkbuf_1
X_7926_ _7926_/CLK _7926_/D vssd1 vssd1 vccd1 vccd1 _7926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7857_ _7857_/CLK _7857_/D vssd1 vssd1 vccd1 vccd1 _7857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7788_ _8617_/Q _7777_/X _7787_/X _7763_/A vssd1 vssd1 vccd1 vccd1 _8617_/D sky130_fd_sc_hd__o211a_1
X_6739_ _6739_/A vssd1 vssd1 vccd1 vccd1 _8098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8409_ _8409_/CLK _8409_/D vssd1 vssd1 vccd1 vccd1 _8409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5070_ _4475_/X _8218_/Q _5072_/S vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4021_ _8534_/Q _3946_/X _4023_/S vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5972_ _5972_/A vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6796__350 _6796__350/A vssd1 vssd1 vccd1 vccd1 _8142_/CLK sky130_fd_sc_hd__inv_2
X_4923_ _4827_/X _4921_/X _4922_/X vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7711_ _7711_/A vssd1 vssd1 vccd1 vccd1 _8571_/D sky130_fd_sc_hd__clkbuf_1
X_4854_ _4853_/X _7931_/Q _7856_/Q _4829_/X vssd1 vssd1 vccd1 vccd1 _4854_/X sky130_fd_sc_hd__a22o_1
X_7642_ _7642_/A vssd1 vssd1 vccd1 vccd1 _7642_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7573_ _7573_/A _7573_/B _7573_/C _7573_/D vssd1 vssd1 vccd1 vccd1 _7573_/X sky130_fd_sc_hd__and4_1
X_4785_ _4671_/X _8266_/Q _4988_/A _4784_/X _4741_/X vssd1 vssd1 vccd1 vccd1 _4785_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6524_ _6032_/A _7967_/Q _6526_/S vssd1 vssd1 vccd1 vccd1 _6525_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6455_ _6494_/B vssd1 vssd1 vccd1 vccd1 _6471_/B sky130_fd_sc_hd__clkbuf_1
X_5406_ _5406_/A vssd1 vssd1 vccd1 vccd1 _8186_/D sky130_fd_sc_hd__clkbuf_1
X_6386_ _8607_/Q vssd1 vssd1 vccd1 vccd1 _6386_/Y sky130_fd_sc_hd__inv_2
X_8125_ _8125_/CLK _8125_/D vssd1 vssd1 vccd1 vccd1 _8125_/Q sky130_fd_sc_hd__dfxtp_1
X_5337_ _3974_/X _5078_/A _5336_/X _5303_/X vssd1 vssd1 vccd1 vccd1 _8208_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8056_ _8056_/CLK _8056_/D vssd1 vssd1 vccd1 vccd1 _8056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5268_ _3968_/X _5078_/X _5267_/X _5152_/X vssd1 vssd1 vccd1 vccd1 _8210_/D sky130_fd_sc_hd__o211a_1
X_4219_ _4219_/A vssd1 vssd1 vccd1 vccd1 _8476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7007_ _7072_/A vssd1 vssd1 vccd1 vccd1 _7007_/X sky130_fd_sc_hd__buf_1
X_5199_ _5095_/X _5196_/X _5198_/X vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0_0__3452_ clkbuf_0__3452_/X vssd1 vssd1 vccd1 vccd1 _7089__489/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7909_ _7909_/CLK _7909_/D vssd1 vssd1 vccd1 vccd1 _7909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6973__402 _6975__404/A vssd1 vssd1 vccd1 vccd1 _8206_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7034__447 _7034__447/A vssd1 vssd1 vccd1 vccd1 _8254_/CLK sky130_fd_sc_hd__inv_2
X_4570_ _4570_/A vssd1 vssd1 vccd1 vccd1 _8312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6240_ _6423_/A vssd1 vssd1 vccd1 vccd1 _6240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6171_ _7885_/Q _6159_/X _6163_/X _6170_/X _6157_/X vssd1 vssd1 vccd1 vccd1 _6171_/X
+ sky130_fd_sc_hd__o221a_1
X_5122_ _5283_/S vssd1 vssd1 vccd1 vccd1 _5122_/X sky130_fd_sc_hd__buf_2
XFILLER_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5053_ _8225_/Q _4531_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4004_ _4004_/A _5382_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5376_/B sky130_fd_sc_hd__and3_1
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5955_ _5955_/A vssd1 vssd1 vccd1 vccd1 _5955_/X sky130_fd_sc_hd__clkbuf_1
X_5886_ _4197_/X _7858_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__mux2_1
X_4906_ _8418_/Q _4855_/X _8226_/Q _4856_/X _4834_/X vssd1 vssd1 vccd1 vccd1 _4906_/X
+ sky130_fd_sc_hd__o221a_1
X_6690__307 _6690__307/A vssd1 vssd1 vccd1 vccd1 _8075_/CLK sky130_fd_sc_hd__inv_2
X_4837_ _8346_/Q _4812_/X _4665_/X _8059_/Q vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__a22o_1
X_7625_ _7647_/A vssd1 vssd1 vccd1 vccd1 _7625_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4768_ _8458_/Q _8348_/Q _8061_/Q _8482_/Q _4691_/X _4694_/X vssd1 vssd1 vccd1 vccd1
+ _4768_/X sky130_fd_sc_hd__mux4_1
X_7556_ _7554_/B _7554_/C _7589_/A vssd1 vssd1 vccd1 vccd1 _7556_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4699_ _4801_/S vssd1 vssd1 vccd1 vccd1 _4699_/X sky130_fd_sc_hd__buf_2
X_6507_ _6014_/A _7959_/Q _6515_/S vssd1 vssd1 vccd1 vccd1 _6508_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6438_ _7942_/Q _6430_/A _6265_/X vssd1 vssd1 vccd1 vccd1 _6438_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8108_ _8108_/CLK _8108_/D vssd1 vssd1 vccd1 vccd1 _8108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6369_ _7959_/Q _7967_/Q _7968_/Q vssd1 vssd1 vccd1 vccd1 _7790_/D sky130_fd_sc_hd__or3_1
XFILLER_76_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8039_ _8039_/CLK _8039_/D vssd1 vssd1 vccd1 vccd1 _8039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3435_ clkbuf_0__3435_/X vssd1 vssd1 vccd1 vccd1 _7072_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7040__451 _7041__452/A vssd1 vssd1 vccd1 vccd1 _8258_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5740_ _8014_/Q _5624_/X _5746_/S vssd1 vssd1 vccd1 vccd1 _5741_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5671_/A vssd1 vssd1 vccd1 vccd1 _8045_/D sky130_fd_sc_hd__clkbuf_1
X_7410_ _7410_/A vssd1 vssd1 vccd1 vccd1 _7411_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8390_ _8390_/CLK _8390_/D vssd1 vssd1 vccd1 vccd1 _8390_/Q sky130_fd_sc_hd__dfxtp_1
X_4622_ _4622_/A vssd1 vssd1 vccd1 vccd1 _8289_/D sky130_fd_sc_hd__clkbuf_1
X_4553_ _5663_/A vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__clkbuf_4
X_4484_ _8342_/Q _4481_/X _4496_/S vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7272_ _7569_/A _7373_/A _7373_/B vssd1 vssd1 vccd1 vccd1 _7330_/A sky130_fd_sc_hd__nand3_1
X_6223_ _7901_/Q _7902_/Q vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__or2b_1
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6136_/X _6152_/X _6153_/X _6139_/X vssd1 vssd1 vccd1 vccd1 _6154_/X sky130_fd_sc_hd__o211a_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5391_/B sky130_fd_sc_hd__buf_2
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _7862_/Q _6088_/B vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__or2_1
XFILLER_111_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5036_ _5036_/A vssd1 vssd1 vccd1 vccd1 _8233_/D sky130_fd_sc_hd__clkbuf_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6987_ _6987_/A vssd1 vssd1 vccd1 vccd1 _8216_/D sky130_fd_sc_hd__clkbuf_1
X_5938_ _5995_/A vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0_0__3082_ clkbuf_0__3082_/X vssd1 vssd1 vccd1 vccd1 _6568__225/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5869_ _5869_/A vssd1 vssd1 vccd1 vccd1 _7909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7608_ _7604_/X _7608_/B vssd1 vssd1 vccd1 vccd1 _7608_/X sky130_fd_sc_hd__and2b_1
X_8588_ _8588_/CLK _8588_/D vssd1 vssd1 vccd1 vccd1 _8588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput101 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _7815_/A sky130_fd_sc_hd__buf_4
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7196__75 _7196__75/A vssd1 vssd1 vccd1 vccd1 _8384_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6910_ _8561_/Q _8560_/Q _8559_/Q vssd1 vssd1 vccd1 vccd1 _7681_/B sky130_fd_sc_hd__and3_2
X_7890_ _8561_/CLK _7890_/D vssd1 vssd1 vccd1 vccd1 _7890_/Q sky130_fd_sc_hd__dfxtp_1
X_6841_ _6843_/C vssd1 vssd1 vccd1 vccd1 _6886_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8511_ _8511_/CLK _8511_/D vssd1 vssd1 vccd1 vccd1 _8511_/Q sky130_fd_sc_hd__dfxtp_1
X_3984_ _5539_/A _5467_/A vssd1 vssd1 vccd1 vccd1 _4000_/S sky130_fd_sc_hd__or2_2
X_5723_ _5723_/A vssd1 vssd1 vccd1 vccd1 _8022_/D sky130_fd_sc_hd__clkbuf_1
X_5654_ _5654_/A vssd1 vssd1 vccd1 vccd1 _8060_/D sky130_fd_sc_hd__clkbuf_1
X_8442_ _8452_/CLK _8442_/D vssd1 vssd1 vccd1 vccd1 _8442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8373_ _8373_/CLK _8373_/D vssd1 vssd1 vccd1 vccd1 _8373_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3452_ _7085_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3452_/X sky130_fd_sc_hd__clkbuf_16
X_4605_ _4475_/X _8296_/Q _4607_/S vssd1 vssd1 vccd1 vccd1 _4606_/A sky130_fd_sc_hd__mux2_1
X_5585_ _5416_/X _8107_/Q _5585_/S vssd1 vssd1 vccd1 vccd1 _5586_/A sky130_fd_sc_hd__mux2_1
X_7324_ _7324_/A _7324_/B _7324_/C vssd1 vssd1 vccd1 vccd1 _7324_/X sky130_fd_sc_hd__and3_1
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4536_ _4427_/X _8326_/Q _4544_/S vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__mux2_1
X_7047__457 _7049__459/A vssd1 vssd1 vccd1 vccd1 _8264_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4467_ _4466_/X _8347_/Q _4470_/S vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__mux2_1
X_7255_ _7266_/A vssd1 vssd1 vccd1 vccd1 _7308_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4398_ _4398_/A vssd1 vssd1 vccd1 vccd1 _8372_/D sky130_fd_sc_hd__clkbuf_1
X_6206_ _6212_/A vssd1 vssd1 vccd1 vccd1 _6206_/X sky130_fd_sc_hd__buf_1
X_6137_ _7951_/Q input9/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6137_/X sky130_fd_sc_hd__mux2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6068_/A vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5019_ _5682_/A _5772_/B vssd1 vssd1 vccd1 vccd1 _5035_/S sky130_fd_sc_hd__nor2_2
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7465__139 _7466__140/A vssd1 vssd1 vccd1 vccd1 _8478_/CLK sky130_fd_sc_hd__inv_2
X_6790__345 _6790__345/A vssd1 vssd1 vccd1 vccd1 _8137_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5370_ _5370_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5377_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4321_ _4321_/A vssd1 vssd1 vccd1 vccd1 _8406_/D sky130_fd_sc_hd__clkbuf_1
X_4252_ _4252_/A vssd1 vssd1 vccd1 vccd1 _8464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _4454_/A _4259_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4183_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7942_ _8610_/CLK _7942_/D vssd1 vssd1 vccd1 vccd1 _7942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7873_ _8623_/CLK _7873_/D vssd1 vssd1 vccd1 vccd1 _7873_/Q sky130_fd_sc_hd__dfxtp_1
X_3967_ _3967_/A vssd1 vssd1 vccd1 vccd1 _8590_/D sky130_fd_sc_hd__clkbuf_1
X_5706_ _5601_/X _8029_/Q _5710_/S vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3467_ clkbuf_0__3467_/X vssd1 vssd1 vccd1 vccd1 _7448_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8425_ _8440_/CLK _8425_/D vssd1 vssd1 vccd1 vccd1 _8425_/Q sky130_fd_sc_hd__dfxtp_1
X_3898_ _8202_/Q _3983_/B _5074_/A _3897_/Y vssd1 vssd1 vccd1 vccd1 _3899_/D sky130_fd_sc_hd__a31o_1
X_7227__100 _7226__99/A vssd1 vssd1 vccd1 vccd1 _8409_/CLK sky130_fd_sc_hd__inv_2
X_5637_ _8066_/Q _5636_/X _5643_/S vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__mux2_1
X_7129__521 _7133__525/A vssd1 vssd1 vccd1 vccd1 _8330_/CLK sky130_fd_sc_hd__inv_2
X_8356_ _8356_/CLK _8356_/D vssd1 vssd1 vccd1 vccd1 _8356_/Q sky130_fd_sc_hd__dfxtp_1
X_5568_ _5568_/A vssd1 vssd1 vccd1 vccd1 _8115_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3435_ _7006_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3435_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4519_ _8192_/Q vssd1 vssd1 vccd1 vccd1 _4519_/X sky130_fd_sc_hd__buf_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8287_ _8287_/CLK _8287_/D vssd1 vssd1 vccd1 vccd1 _8287_/Q sky130_fd_sc_hd__dfxtp_1
X_7307_ _7590_/A _7281_/X _7306_/X vssd1 vssd1 vccd1 vccd1 _7307_/Y sky130_fd_sc_hd__a21boi_1
X_5499_ _8148_/Q _4501_/X _5501_/S vssd1 vssd1 vccd1 vccd1 _5500_/A sky130_fd_sc_hd__mux2_1
X_7238_ _8443_/Q _8416_/Q _7407_/C vssd1 vssd1 vccd1 vccd1 _7399_/B sky130_fd_sc_hd__and3_1
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4870_ _4737_/X _4864_/X _4868_/X _4869_/X _4673_/A vssd1 vssd1 vccd1 vccd1 _4870_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3321_ clkbuf_0__3321_/X vssd1 vssd1 vccd1 vccd1 _6821__365/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6540_ _8089_/Q _7974_/Q _6548_/S vssd1 vssd1 vccd1 vccd1 _6541_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3252_ clkbuf_0__3252_/X vssd1 vssd1 vccd1 vccd1 _6606__255/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6471_ _8620_/Q _6471_/B _6481_/C vssd1 vssd1 vccd1 vccd1 _6471_/X sky130_fd_sc_hd__and3_1
X_5422_ _5422_/A vssd1 vssd1 vccd1 vccd1 _8182_/D sky130_fd_sc_hd__clkbuf_1
X_8210_ _8210_/CLK _8210_/D vssd1 vssd1 vccd1 vccd1 _8210_/Q sky130_fd_sc_hd__dfxtp_1
X_8141_ _8141_/CLK _8141_/D vssd1 vssd1 vccd1 vccd1 _8141_/Q sky130_fd_sc_hd__dfxtp_1
X_5353_ _5254_/X _8155_/Q _7920_/Q _5249_/A _5135_/A vssd1 vssd1 vccd1 vccd1 _5353_/X
+ sky130_fd_sc_hd__o221a_1
Xoutput202 _6094_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__buf_2
X_4304_ _8413_/Q _4220_/X _4310_/S vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8072_ _8072_/CLK _8072_/D vssd1 vssd1 vccd1 vccd1 _8072_/Q sky130_fd_sc_hd__dfxtp_1
X_5284_ _8353_/Q _5103_/B _5283_/X _5274_/A vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__o22a_1
X_4235_ _8571_/Q vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__buf_2
Xclkbuf_0__3082_ _6353_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3082_/X sky130_fd_sc_hd__clkbuf_16
XINSDIODE2_8 _4212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4166_ _8250_/Q vssd1 vssd1 vccd1 vccd1 _4171_/B sky130_fd_sc_hd__inv_2
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4097_ _8503_/Q _3943_/X _4101_/S vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__mux2_1
X_7925_ _7925_/CLK _7925_/D vssd1 vssd1 vccd1 vccd1 _7925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7856_ _7856_/CLK _7856_/D vssd1 vssd1 vccd1 vccd1 _7856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6918__372 _6920__374/A vssd1 vssd1 vccd1 vccd1 _8168_/CLK sky130_fd_sc_hd__inv_2
X_7787_ _5976_/A _7778_/X _7776_/A vssd1 vssd1 vccd1 vccd1 _7787_/X sky130_fd_sc_hd__a21bo_1
X_4999_ _4691_/X _4988_/X _4998_/Y vssd1 vssd1 vccd1 vccd1 _8250_/D sky130_fd_sc_hd__a21oi_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6738_ _8098_/Q _5998_/A _6742_/S vssd1 vssd1 vccd1 vccd1 _6739_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8408_ _8408_/CLK _8408_/D vssd1 vssd1 vccd1 vccd1 _8408_/Q sky130_fd_sc_hd__dfxtp_1
X_8339_ _8339_/CLK _8339_/D vssd1 vssd1 vccd1 vccd1 _8339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6628__273 _6630__275/A vssd1 vssd1 vccd1 vccd1 _8033_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7884_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _4020_/A vssd1 vssd1 vccd1 vccd1 _8535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5971_ _7799_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5972_/A sky130_fd_sc_hd__or2_1
XFILLER_65_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4922_ _8312_/Q _4815_/X _4838_/X _8296_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4922_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7710_ _7840_/A _7716_/B _7714_/C vssd1 vssd1 vccd1 vccd1 _7711_/A sky130_fd_sc_hd__and3_1
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7641_ _8552_/Q vssd1 vssd1 vccd1 vccd1 _7641_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4853_ _4853_/A vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__buf_2
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4784_ _4683_/X _4771_/X _4775_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__a31o_2
X_7572_ _7814_/A _7551_/Y _7557_/X _7565_/Y _7571_/X vssd1 vssd1 vccd1 vccd1 _7573_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_119_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6523_ _6523_/A vssd1 vssd1 vccd1 vccd1 _7966_/D sky130_fd_sc_hd__clkbuf_1
X_6454_ _6454_/A vssd1 vssd1 vccd1 vccd1 _6494_/B sky130_fd_sc_hd__clkbuf_2
X_5405_ _5404_/X _8186_/Q _5417_/S vssd1 vssd1 vccd1 vccd1 _5406_/A sky130_fd_sc_hd__mux2_1
X_6385_ _6385_/A vssd1 vssd1 vccd1 vccd1 _6385_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8124_ _8124_/CLK _8124_/D vssd1 vssd1 vccd1 vccd1 _8124_/Q sky130_fd_sc_hd__dfxtp_1
X_5336_ _8208_/Q _5081_/A _5386_/A _5335_/Y _5148_/A vssd1 vssd1 vccd1 vccd1 _5336_/X
+ sky130_fd_sc_hd__a221o_1
X_8055_ _8608_/CLK _8055_/D vssd1 vssd1 vccd1 vccd1 _8055_/Q sky130_fd_sc_hd__dfxtp_1
X_5267_ _8210_/Q _5080_/X _5386_/A _5266_/X _5148_/X vssd1 vssd1 vccd1 vccd1 _5267_/X
+ sky130_fd_sc_hd__a221o_1
X_4218_ _8476_/Q _4215_/X _4230_/S vssd1 vssd1 vccd1 vccd1 _4219_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3451_ clkbuf_0__3451_/X vssd1 vssd1 vccd1 vccd1 _7084__485/A sky130_fd_sc_hd__clkbuf_4
X_7006_ _7541_/A vssd1 vssd1 vccd1 vccd1 _7006_/X sky130_fd_sc_hd__buf_1
X_5198_ _5121_/X _5197_/X _5333_/A vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4149_ _4149_/A vssd1 vssd1 vccd1 vccd1 _8488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7908_ _7908_/CLK _7908_/D vssd1 vssd1 vccd1 vccd1 _7908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7223__96 _7224__97/A vssd1 vssd1 vccd1 vccd1 _8405_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7839_ _6872_/A _7826_/X _7838_/X _6423_/X vssd1 vssd1 vccd1 vccd1 _8631_/D sky130_fd_sc_hd__a211o_1
XFILLER_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3649_ clkbuf_0__3649_/X vssd1 vssd1 vccd1 vccd1 _7471__144/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3020_ clkbuf_0__3020_/X vssd1 vssd1 vccd1 vccd1 _6219__191/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6170_ _6170_/A _6172_/B vssd1 vssd1 vccd1 vccd1 _6170_/X sky130_fd_sc_hd__and2_4
XFILLER_115_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _5142_/S vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _5052_/A vssd1 vssd1 vccd1 vccd1 _8226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4003_ _4299_/A _5373_/A _4027_/B vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__or3b_4
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5954_ _7828_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__or2_1
XFILLER_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6577__231 _6578__232/A vssd1 vssd1 vccd1 vccd1 _7991_/CLK sky130_fd_sc_hd__inv_2
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _7859_/D sky130_fd_sc_hd__clkbuf_1
X_4905_ _4874_/X _8181_/Q _8073_/Q _4853_/X vssd1 vssd1 vccd1 vccd1 _4905_/X sky130_fd_sc_hd__a22o_1
X_4836_ _4827_/X _4830_/X _4835_/X vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__o21a_1
X_7624_ _8548_/Q vssd1 vssd1 vccd1 vccd1 _7624_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7555_ _8622_/Q _7555_/B _7555_/C vssd1 vssd1 vccd1 vccd1 _7555_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6506_ _6550_/A vssd1 vssd1 vccd1 vccd1 _6515_/S sky130_fd_sc_hd__clkbuf_2
X_4767_ _4460_/X _4669_/X _4766_/X _4744_/X vssd1 vssd1 vccd1 vccd1 _8267_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7486_ _7504_/A vssd1 vssd1 vccd1 vccd1 _7486_/X sky130_fd_sc_hd__buf_1
X_4698_ _4724_/A vssd1 vssd1 vccd1 vccd1 _4801_/S sky130_fd_sc_hd__buf_4
X_6437_ _8627_/Q _6363_/X _6452_/A _6435_/X _6436_/Y vssd1 vssd1 vccd1 vccd1 _6437_/X
+ sky130_fd_sc_hd__a32o_1
X_6368_ _6368_/A _6454_/A vssd1 vssd1 vccd1 vccd1 _6501_/B sky130_fd_sc_hd__or2b_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8107_ _8107_/CLK _8107_/D vssd1 vssd1 vccd1 vccd1 _8107_/Q sky130_fd_sc_hd__dfxtp_1
X_5319_ _5389_/B _5315_/Y _5318_/Y _5087_/A vssd1 vssd1 vccd1 vccd1 _5319_/X sky130_fd_sc_hd__a31o_1
X_8660__225 vssd1 vssd1 vccd1 vccd1 _8660__225/HI core1Index[5] sky130_fd_sc_hd__conb_1
XFILLER_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6299_ _6072_/A _6505_/A _6080_/A _7901_/Q vssd1 vssd1 vccd1 vccd1 _6299_/X sky130_fd_sc_hd__a31o_1
X_8038_ _8038_/CLK _8038_/D vssd1 vssd1 vccd1 vccd1 _8038_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3434_ clkbuf_0__3434_/X vssd1 vssd1 vccd1 vccd1 _7002__422/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5670_ _5601_/X _8045_/Q _5674_/S vssd1 vssd1 vccd1 vccd1 _5671_/A sky130_fd_sc_hd__mux2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4621_ _8289_/Q _4498_/X _4625_/S vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__mux2_1
X_4552_ _5663_/B vssd1 vssd1 vccd1 vccd1 _5055_/C sky130_fd_sc_hd__clkbuf_4
X_4483_ _4505_/S vssd1 vssd1 vccd1 vccd1 _4496_/S sky130_fd_sc_hd__buf_2
X_7271_ _8430_/Q _8429_/Q _7266_/A _8431_/Q vssd1 vssd1 vccd1 vccd1 _7373_/B sky130_fd_sc_hd__a31o_1
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8644__209 vssd1 vssd1 vccd1 vccd1 _8644__209/HI caravel_irq[0] sky130_fd_sc_hd__conb_1
X_6222_ _6390_/A vssd1 vssd1 vccd1 vccd1 _6222_/X sky130_fd_sc_hd__buf_4
X_7123__516 _7124__517/A vssd1 vssd1 vccd1 vccd1 _8325_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _7880_/Q _6175_/A vssd1 vssd1 vccd1 vccd1 _6153_/X sky130_fd_sc_hd__or2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5120_/A vssd1 vssd1 vccd1 vccd1 _5165_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _7937_/Q input14/X _6188_/B vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__mux2_1
X_5035_ _8233_/Q _4531_/X _5035_/S vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__mux2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6986_ _8452_/Q _6986_/B _6986_/C _7053_/A vssd1 vssd1 vccd1 vccd1 _6987_/A sky130_fd_sc_hd__and4b_1
X_5937_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3081_ clkbuf_0__3081_/X vssd1 vssd1 vccd1 vccd1 _6351__219/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _7909_/Q _5601_/A _5872_/S vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__mux2_1
X_7607_ _7607_/A _7664_/B _7664_/C vssd1 vssd1 vccd1 vccd1 _7607_/X sky130_fd_sc_hd__and3_1
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5799_ _5799_/A vssd1 vssd1 vccd1 vccd1 _7988_/D sky130_fd_sc_hd__clkbuf_1
X_4819_ _4996_/B _4813_/X _4818_/X vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__o21a_1
X_8587_ _8587_/CLK _8587_/D vssd1 vssd1 vccd1 vccd1 _8587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _6281_/A sky130_fd_sc_hd__buf_6
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7750__48 _7752__50/A vssd1 vssd1 vccd1 vccd1 _8599_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6840_ _6850_/A vssd1 vssd1 vccd1 vccd1 _6842_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_23_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5722_ _8022_/Q _5624_/X _5728_/S vssd1 vssd1 vccd1 vccd1 _5723_/A sky130_fd_sc_hd__mux2_1
X_8510_ _8510_/CLK _8510_/D vssd1 vssd1 vccd1 vccd1 _8510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3983_ _4004_/A _3983_/B _4064_/B _5150_/A vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__or4b_4
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5653_ _5604_/X _8060_/Q _5655_/S vssd1 vssd1 vccd1 vccd1 _5654_/A sky130_fd_sc_hd__mux2_1
X_8441_ _8441_/CLK _8441_/D vssd1 vssd1 vccd1 vccd1 _8441_/Q sky130_fd_sc_hd__dfxtp_1
X_8372_ _8372_/CLK _8372_/D vssd1 vssd1 vccd1 vccd1 _8372_/Q sky130_fd_sc_hd__dfxtp_1
X_5584_ _5584_/A vssd1 vssd1 vccd1 vccd1 _8108_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3451_ _7079_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3451_/X sky130_fd_sc_hd__clkbuf_16
X_4604_ _4604_/A vssd1 vssd1 vccd1 vccd1 _8297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4535_ _4550_/S vssd1 vssd1 vccd1 vccd1 _4544_/S sky130_fd_sc_hd__buf_2
X_7323_ _7303_/A _7303_/B _6901_/A vssd1 vssd1 vccd1 vccd1 _7323_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7254_ _7260_/A vssd1 vssd1 vccd1 vccd1 _7266_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4466_ _8192_/Q vssd1 vssd1 vccd1 vccd1 _4466_/X sky130_fd_sc_hd__clkbuf_4
X_4397_ _4115_/X _8372_/Q _4401_/S vssd1 vssd1 vccd1 vccd1 _4398_/A sky130_fd_sc_hd__mux2_1
X_7185_ _7191_/A vssd1 vssd1 vccd1 vccd1 _7185_/X sky130_fd_sc_hd__buf_1
X_6136_ _6136_/A vssd1 vssd1 vccd1 vccd1 _6136_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6067_ _8098_/Q _6069_/B vssd1 vssd1 vccd1 vccd1 _6068_/A sky130_fd_sc_hd__and2_2
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _5055_/C _5055_/B _5055_/A vssd1 vssd1 vccd1 vccd1 _5772_/B sky130_fd_sc_hd__nand3b_4
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6622__268 _6624__270/A vssd1 vssd1 vccd1 vccd1 _8028_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6325__198 _6325__198/A vssd1 vssd1 vccd1 vccd1 _7910_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3649_ _7467_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3649_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8666__231 vssd1 vssd1 vccd1 vccd1 _8666__231/HI manufacturerID[3] sky130_fd_sc_hd__conb_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4320_ _8406_/Q _4215_/X _4328_/S vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4251_ _8464_/Q _4229_/X _4251_/S vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4182_ _8258_/Q _4716_/A vssd1 vssd1 vccd1 vccd1 _4666_/D sky130_fd_sc_hd__xnor2_1
XFILLER_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7941_ _8610_/CLK _7941_/D vssd1 vssd1 vccd1 vccd1 _7941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7872_ _8625_/CLK _7872_/D vssd1 vssd1 vccd1 vccd1 _7872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6754_ _6760_/A vssd1 vssd1 vccd1 vccd1 _6754_/X sky130_fd_sc_hd__buf_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3966_ _3965_/X _8590_/Q _3969_/S vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__mux2_1
X_5705_ _5705_/A vssd1 vssd1 vccd1 vccd1 _8030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8424_ _8424_/CLK _8424_/D vssd1 vssd1 vccd1 vccd1 _8424_/Q sky130_fd_sc_hd__dfxtp_1
X_7175__57 _7178__60/A vssd1 vssd1 vccd1 vccd1 _8366_/CLK sky130_fd_sc_hd__inv_2
X_5636_ _8190_/Q vssd1 vssd1 vccd1 vccd1 _5636_/X sky130_fd_sc_hd__clkbuf_2
X_3897_ _5075_/B _5370_/A _3887_/Y vssd1 vssd1 vccd1 vccd1 _3897_/Y sky130_fd_sc_hd__a21oi_1
X_8355_ _8355_/CLK _8355_/D vssd1 vssd1 vccd1 vccd1 _8355_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3434_ _7000_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3434_/X sky130_fd_sc_hd__clkbuf_16
X_5567_ _5416_/X _8115_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5568_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4518_ _4518_/A vssd1 vssd1 vccd1 vccd1 _8332_/D sky130_fd_sc_hd__clkbuf_1
X_5498_ _5498_/A vssd1 vssd1 vccd1 vccd1 _8149_/D sky130_fd_sc_hd__clkbuf_1
X_8286_ _8286_/CLK _8286_/D vssd1 vssd1 vccd1 vccd1 _8286_/Q sky130_fd_sc_hd__dfxtp_1
X_7306_ _8621_/Q _7306_/B _7303_/B vssd1 vssd1 vccd1 vccd1 _7306_/X sky130_fd_sc_hd__or3b_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4449_ _4449_/A vssd1 vssd1 vccd1 vccd1 _8352_/D sky130_fd_sc_hd__clkbuf_1
X_7237_ _8442_/Q _8441_/Q vssd1 vssd1 vccd1 vccd1 _7407_/C sky130_fd_sc_hd__and2_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6119_ _7871_/Q _6126_/B vssd1 vssd1 vccd1 vccd1 _6119_/X sky130_fd_sc_hd__or2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7234__105 _7234__105/A vssd1 vssd1 vccd1 vccd1 _8414_/CLK sky130_fd_sc_hd__inv_2
X_7136__526 _7139__529/A vssd1 vssd1 vccd1 vccd1 _8335_/CLK sky130_fd_sc_hd__inv_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8640__256 vssd1 vssd1 vccd1 vccd1 partID[10] _8640__256/LO sky130_fd_sc_hd__conb_1
X_7471__144 _7471__144/A vssd1 vssd1 vccd1 vccd1 _8483_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3320_ clkbuf_0__3320_/X vssd1 vssd1 vccd1 vccd1 _6813__358/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3251_ clkbuf_0__3251_/X vssd1 vssd1 vccd1 vccd1 _6625_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6571__226 _6572__227/A vssd1 vssd1 vccd1 vccd1 _7986_/CLK sky130_fd_sc_hd__inv_2
X_6470_ _7948_/Q _6464_/X _6452_/X _6469_/X _6459_/X vssd1 vssd1 vccd1 vccd1 _7948_/D
+ sky130_fd_sc_hd__a221o_1
X_5421_ _5420_/X _8182_/Q _5429_/S vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__mux2_1
X_8140_ _8140_/CLK _8140_/D vssd1 vssd1 vccd1 vccd1 _8140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5352_ _8407_/Q _8128_/Q _5352_/S vssd1 vssd1 vccd1 vccd1 _5352_/X sky130_fd_sc_hd__mux2_1
Xoutput203 _6097_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__buf_2
X_8071_ _8071_/CLK _8071_/D vssd1 vssd1 vccd1 vccd1 _8071_/Q sky130_fd_sc_hd__dfxtp_1
X_4303_ _4303_/A vssd1 vssd1 vccd1 vccd1 _8414_/D sky130_fd_sc_hd__clkbuf_1
X_5283_ _8401_/Q _8138_/Q _5283_/S vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__mux2_2
XFILLER_99_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4234_ _4234_/A vssd1 vssd1 vccd1 vccd1 _8471_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3081_ _6347_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3081_/X sky130_fd_sc_hd__clkbuf_16
XINSDIODE2_9 _4212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4165_ _7838_/A _4164_/X _6193_/A vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__a21oi_4
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4096_/A vssd1 vssd1 vccd1 vccd1 _8504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7924_ _7924_/CLK _7924_/D vssd1 vssd1 vccd1 vccd1 _7924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7855_ _7855_/CLK _7855_/D vssd1 vssd1 vccd1 vccd1 _7855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7786_ _7053_/A _7777_/X _7785_/X _6503_/X vssd1 vssd1 vccd1 vccd1 _8616_/D sky130_fd_sc_hd__o211a_1
X_4998_ _4691_/X _4996_/A _4964_/X vssd1 vssd1 vccd1 vccd1 _4998_/Y sky130_fd_sc_hd__o21ai_1
X_3949_ _8570_/Q vssd1 vssd1 vccd1 vccd1 _3949_/X sky130_fd_sc_hd__buf_2
X_6737_ _6737_/A vssd1 vssd1 vccd1 vccd1 _8097_/D sky130_fd_sc_hd__clkbuf_1
X_6668_ _6668_/A vssd1 vssd1 vccd1 vccd1 _6668_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3449_ clkbuf_0__3449_/X vssd1 vssd1 vccd1 vccd1 _7079_/A sky130_fd_sc_hd__clkbuf_4
X_5619_ _8195_/Q vssd1 vssd1 vccd1 vccd1 _5619_/X sky130_fd_sc_hd__buf_2
X_8407_ _8407_/CLK _8407_/D vssd1 vssd1 vccd1 vccd1 _8407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8338_ _8338_/CLK _8338_/D vssd1 vssd1 vccd1 vccd1 _8338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8269_ _8270_/CLK _8269_/D vssd1 vssd1 vccd1 vccd1 _8269_/Q sky130_fd_sc_hd__dfxtp_1
X_6667__290 _6667__290/A vssd1 vssd1 vccd1 vccd1 _8058_/CLK sky130_fd_sc_hd__inv_2
X_6925__377 _6927__379/A vssd1 vssd1 vccd1 vccd1 _8173_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7519__7 _7519__7/A vssd1 vssd1 vccd1 vccd1 _8521_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6635__278 _6637__280/A vssd1 vssd1 vccd1 vccd1 _8038_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5970_ _5970_/A vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _8280_/Q _4874_/X _4822_/X _8242_/Q vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4852_ _4852_/A vssd1 vssd1 vccd1 vccd1 _4853_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7640_ _7640_/A vssd1 vssd1 vccd1 vccd1 _8551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4783_ _4777_/X _4779_/X _4782_/X _4735_/X _4737_/X vssd1 vssd1 vccd1 vccd1 _4783_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7571_ _7566_/X _7567_/Y _7568_/X _7569_/Y _7570_/X vssd1 vssd1 vccd1 vccd1 _7571_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6522_ _6030_/A _7966_/Q _6526_/S vssd1 vssd1 vccd1 vccd1 _6523_/A sky130_fd_sc_hd__mux2_1
X_6453_ _8624_/Q vssd1 vssd1 vccd1 vccd1 _7814_/A sky130_fd_sc_hd__buf_2
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5404_ _5598_/A vssd1 vssd1 vccd1 vccd1 _5404_/X sky130_fd_sc_hd__clkbuf_2
X_8123_ _8123_/CLK _8123_/D vssd1 vssd1 vccd1 vccd1 _8123_/Q sky130_fd_sc_hd__dfxtp_1
X_6384_ _6384_/A _6384_/B vssd1 vssd1 vccd1 vccd1 _6385_/A sky130_fd_sc_hd__or2_1
X_5335_ _5335_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5335_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5266_ _5387_/B _5243_/X _5247_/X _5265_/X vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__a31o_2
X_8054_ _8608_/CLK _8054_/D vssd1 vssd1 vccd1 vccd1 _8054_/Q sky130_fd_sc_hd__dfxtp_1
X_4217_ _4239_/S vssd1 vssd1 vccd1 vccd1 _4230_/S sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0__3450_ clkbuf_0__3450_/X vssd1 vssd1 vccd1 vccd1 _7078__480/A sky130_fd_sc_hd__clkbuf_4
X_5197_ _8521_/Q _8513_/Q _7916_/Q _8529_/Q _5122_/X _5123_/X vssd1 vssd1 vccd1 vccd1
+ _5197_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4148_ _8488_/Q _3940_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4079_ _4079_/A vssd1 vssd1 vccd1 vccd1 _8511_/D sky130_fd_sc_hd__clkbuf_1
X_7907_ _7907_/CLK _7907_/D vssd1 vssd1 vccd1 vccd1 _7907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7838_ _7838_/A _7842_/B _7840_/C vssd1 vssd1 vccd1 vccd1 _7838_/X sky130_fd_sc_hd__and3_1
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7769_ _7771_/A _8605_/Q vssd1 vssd1 vccd1 vccd1 _7770_/A sky130_fd_sc_hd__and2_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3648_ clkbuf_0__3648_/X vssd1 vssd1 vccd1 vccd1 _7466__140/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6980__408 _6980__408/A vssd1 vssd1 vccd1 vccd1 _8212_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ _5120_/A vssd1 vssd1 vccd1 vccd1 _5142_/S sky130_fd_sc_hd__buf_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _8226_/Q _4528_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _5052_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4336_/A vssd1 vssd1 vccd1 vccd1 _4299_/A sky130_fd_sc_hd__buf_2
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5953_ _5953_/A vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _4194_/X _7859_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4904_ _4472_/X _4669_/A _4902_/X _4903_/X vssd1 vssd1 vccd1 vccd1 _8263_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7484__154 _7485__155/A vssd1 vssd1 vccd1 vccd1 _8493_/CLK sky130_fd_sc_hd__inv_2
X_4835_ _8314_/Q _4831_/X _4833_/X _8298_/Q _4834_/X vssd1 vssd1 vccd1 vccd1 _4835_/X
+ sky130_fd_sc_hd__o221a_1
X_7623_ _7623_/A vssd1 vssd1 vccd1 vccd1 _8547_/D sky130_fd_sc_hd__clkbuf_1
X_6989__411 _6993__415/A vssd1 vssd1 vccd1 vccd1 _8217_/CLK sky130_fd_sc_hd__inv_2
X_7554_ _7589_/A _7554_/B _7554_/C vssd1 vssd1 vccd1 vccd1 _7554_/Y sky130_fd_sc_hd__nand3_1
X_4766_ _4671_/X _8267_/Q _4988_/A _4765_/X _4741_/X vssd1 vssd1 vccd1 vccd1 _4766_/X
+ sky130_fd_sc_hd__a221o_1
X_6505_ _6505_/A _6505_/B _7844_/D vssd1 vssd1 vccd1 vccd1 _6550_/A sky130_fd_sc_hd__nand3_4
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4697_ _4834_/A vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6436_ _6474_/A _6436_/B vssd1 vssd1 vccd1 vccd1 _6436_/Y sky130_fd_sc_hd__nor2_1
X_6367_ _7790_/A _7790_/C vssd1 vssd1 vccd1 vccd1 _6371_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3079_ clkbuf_0__3079_/X vssd1 vssd1 vccd1 vccd1 _6338__208/A sky130_fd_sc_hd__clkbuf_4
X_8106_ _8106_/CLK _8106_/D vssd1 vssd1 vccd1 vccd1 _8106_/Q sky130_fd_sc_hd__dfxtp_1
X_5318_ _5233_/X _5316_/X _5317_/X vssd1 vssd1 vccd1 vccd1 _5318_/Y sky130_fd_sc_hd__o21ai_1
X_6330__201 _6331__202/A vssd1 vssd1 vccd1 vccd1 _7913_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6217__190 _6217__190/A vssd1 vssd1 vccd1 vccd1 _7859_/CLK sky130_fd_sc_hd__inv_2
X_6298_ _6298_/A vssd1 vssd1 vccd1 vccd1 _7900_/D sky130_fd_sc_hd__clkbuf_1
X_8037_ _8037_/CLK _8037_/D vssd1 vssd1 vccd1 vccd1 _8037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5249_ _5249_/A vssd1 vssd1 vccd1 vccd1 _5249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8604_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3433_ clkbuf_0__3433_/X vssd1 vssd1 vccd1 vccd1 _6999__420/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4620_ _4620_/A vssd1 vssd1 vccd1 vccd1 _8290_/D sky130_fd_sc_hd__clkbuf_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _8319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4482_ _4534_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _4505_/S sky130_fd_sc_hd__nor2_2
X_7270_ _8431_/Q _7274_/A _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _7373_/A sky130_fd_sc_hd__nand4_1
X_8683__248 vssd1 vssd1 vccd1 vccd1 _8683__248/HI versionID[2] sky130_fd_sc_hd__conb_1
X_6221_ _6647_/A vssd1 vssd1 vccd1 vccd1 _6390_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6152_ _7955_/Q input13/X _6177_/A vssd1 vssd1 vccd1 vccd1 _6152_/X sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5103_ _5112_/B _5103_/B vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__or2_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6073_/X _6076_/X _6079_/X _6082_/X vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5034_ _5034_/A vssd1 vssd1 vccd1 vccd1 _8234_/D sky130_fd_sc_hd__clkbuf_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6985_ _6500_/A _7757_/B _6363_/X _7714_/C vssd1 vssd1 vccd1 vccd1 _8215_/D sky130_fd_sc_hd__o211a_1
X_5936_ _6732_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__and2_1
X_7017__433 _7017__433/A vssd1 vssd1 vccd1 vccd1 _8239_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3080_ clkbuf_0__3080_/X vssd1 vssd1 vccd1 vccd1 _6343__212/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5867_ _5867_/A vssd1 vssd1 vccd1 vccd1 _7910_/D sky130_fd_sc_hd__clkbuf_1
X_7606_ _7603_/Y _7604_/X _7605_/X vssd1 vssd1 vccd1 vccd1 _8543_/D sky130_fd_sc_hd__a21oi_1
XFILLER_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5798_ _7988_/Q _5604_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5799_/A sky130_fd_sc_hd__mux2_1
X_4818_ _8420_/Q _4815_/X _8228_/Q _4817_/X _4699_/X vssd1 vssd1 vccd1 vccd1 _4818_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8586_ _8586_/CLK _8586_/D vssd1 vssd1 vccd1 vccd1 _8586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4749_ _4994_/B _4746_/X _4748_/X vssd1 vssd1 vccd1 vccd1 _4749_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6419_ _8611_/Q vssd1 vssd1 vccd1 vccd1 _6419_/Y sky130_fd_sc_hd__inv_2
X_7399_ _8415_/Q _7399_/B vssd1 vssd1 vccd1 vccd1 _7399_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _6696_/A sky130_fd_sc_hd__buf_6
XFILLER_102_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6337__207 _6340__210/A vssd1 vssd1 vccd1 vccd1 _7919_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7435__115 _7435__115/A vssd1 vssd1 vccd1 vccd1 _8454_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _5147_/A _7757_/B vssd1 vssd1 vccd1 vccd1 _4064_/B sky130_fd_sc_hd__nand2_1
X_5721_ _5721_/A vssd1 vssd1 vccd1 vccd1 _8023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5652_ _5652_/A vssd1 vssd1 vccd1 vccd1 _8061_/D sky130_fd_sc_hd__clkbuf_1
X_8440_ _8440_/CLK _8440_/D vssd1 vssd1 vccd1 vccd1 _8440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5583_ _5412_/X _8108_/Q _5585_/S vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__mux2_1
X_8371_ _8371_/CLK _8371_/D vssd1 vssd1 vccd1 vccd1 _8371_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3450_ _7073_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3450_/X sky130_fd_sc_hd__clkbuf_16
X_4603_ _4472_/X _8297_/Q _4607_/S vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__mux2_1
X_4534_ _4534_/A _5844_/A vssd1 vssd1 vccd1 vccd1 _4550_/S sky130_fd_sc_hd__or2_4
X_7322_ _7590_/A _7281_/X _7299_/Y _7300_/X _7306_/X vssd1 vssd1 vccd1 vccd1 _7327_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7086__486 _7089__489/A vssd1 vssd1 vccd1 vccd1 _8295_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ _4465_/A vssd1 vssd1 vccd1 vccd1 _8348_/D sky130_fd_sc_hd__clkbuf_1
X_7253_ _8626_/Q vssd1 vssd1 vccd1 vccd1 _7324_/A sky130_fd_sc_hd__inv_2
X_4396_ _4396_/A vssd1 vssd1 vccd1 vccd1 _8373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6135_ _6117_/X _6133_/X _6134_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6135_/X sky130_fd_sc_hd__o211a_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6066_/A vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5017_ _5017_/A vssd1 vssd1 vccd1 vccd1 _8241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6899_ _8621_/Q vssd1 vssd1 vccd1 vccd1 _6901_/A sky130_fd_sc_hd__clkinv_2
X_5919_ _8096_/Q _8097_/Q _8098_/Q _8099_/Q vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__and4_2
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3648_ _7461_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3648_/X sky130_fd_sc_hd__clkbuf_16
X_8569_ _8569_/CLK _8569_/D vssd1 vssd1 vccd1 vccd1 _8569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4250_ _4250_/A vssd1 vssd1 vccd1 vccd1 _8465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4181_ _8253_/Q vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7940_ _8610_/CLK _7940_/D vssd1 vssd1 vccd1 vccd1 _7940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7871_ _8625_/CLK _7871_/D vssd1 vssd1 vccd1 vccd1 _7871_/Q sky130_fd_sc_hd__dfxtp_1
X_6822_ _6822_/A vssd1 vssd1 vccd1 vccd1 _6822_/X sky130_fd_sc_hd__buf_1
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3965_ _8574_/Q vssd1 vssd1 vccd1 vccd1 _3965_/X sky130_fd_sc_hd__clkbuf_4
X_5704_ _5598_/X _8030_/Q _5710_/S vssd1 vssd1 vccd1 vccd1 _5705_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3465_ clkbuf_0__3465_/X vssd1 vssd1 vccd1 vccd1 _7158__545/A sky130_fd_sc_hd__clkbuf_4
X_3896_ _3893_/Y _3895_/X _5370_/A vssd1 vssd1 vccd1 vccd1 _3899_/C sky130_fd_sc_hd__a21oi_1
X_8423_ _8423_/CLK _8423_/D vssd1 vssd1 vccd1 vccd1 _8423_/Q sky130_fd_sc_hd__dfxtp_1
X_5635_ _5635_/A vssd1 vssd1 vccd1 vccd1 _8067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3433_ _6994_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3433_/X sky130_fd_sc_hd__clkbuf_16
X_5566_ _5566_/A vssd1 vssd1 vccd1 vccd1 _8116_/D sky130_fd_sc_hd__clkbuf_1
X_8354_ _8354_/CLK _8354_/D vssd1 vssd1 vccd1 vccd1 _8354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4517_ _8332_/Q _4516_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5497_ _8149_/Q _4498_/X _5501_/S vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__mux2_1
X_8285_ _8285_/CLK _8285_/D vssd1 vssd1 vccd1 vccd1 _8285_/Q sky130_fd_sc_hd__dfxtp_1
X_7305_ _8624_/Q vssd1 vssd1 vccd1 vccd1 _7590_/A sky130_fd_sc_hd__clkbuf_4
X_4448_ _4447_/X _8352_/Q _4451_/S vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__mux2_1
X_7236_ _7432_/S vssd1 vssd1 vccd1 vccd1 _7420_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _8380_/Q _4223_/X _4383_/S vssd1 vssd1 vccd1 vccd1 _4380_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7167_ _7173_/A vssd1 vssd1 vccd1 vccd1 _7167_/X sky130_fd_sc_hd__buf_1
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _7946_/Q input4/X _6125_/S vssd1 vssd1 vccd1 vccd1 _6118_/X sky130_fd_sc_hd__mux2_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6058_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7505__171 _7506__172/A vssd1 vssd1 vccd1 vccd1 _8510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3250_ clkbuf_0__3250_/X vssd1 vssd1 vccd1 vccd1 _6596__247/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5420_ _5610_/A vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5351_ _5351_/A _5351_/B _5351_/C vssd1 vssd1 vccd1 vccd1 _5351_/X sky130_fd_sc_hd__or3_1
Xoutput204 _6102_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__buf_2
X_8070_ _8070_/CLK _8070_/D vssd1 vssd1 vccd1 vccd1 _8070_/Q sky130_fd_sc_hd__dfxtp_1
X_4302_ _8414_/Q _4215_/X _4310_/S vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__mux2_1
X_7180__61 _7184__65/A vssd1 vssd1 vccd1 vccd1 _8370_/CLK sky130_fd_sc_hd__inv_2
X_5282_ _5269_/X _5280_/X _5281_/X vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__o21a_1
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _8471_/Q _4232_/X _4239_/S vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3080_ _6341_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3080_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4164_ _6077_/A _6080_/A _4164_/C vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__and3_4
X_4095_ _8504_/Q _3940_/X _4095_/S vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7923_ _7923_/CLK _7923_/D vssd1 vssd1 vccd1 vccd1 _7923_/Q sky130_fd_sc_hd__dfxtp_1
X_6211__185 _6211__185/A vssd1 vssd1 vccd1 vccd1 _7854_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7854_ _7854_/CLK _7854_/D vssd1 vssd1 vccd1 vccd1 _7854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6805_ _6805_/A vssd1 vssd1 vccd1 vccd1 _8146_/D sky130_fd_sc_hd__clkbuf_1
X_7785_ _5978_/A _7778_/X _7777_/A vssd1 vssd1 vccd1 vccd1 _7785_/X sky130_fd_sc_hd__a21bo_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6736_ _8097_/Q _5996_/A _6742_/S vssd1 vssd1 vccd1 vccd1 _6737_/A sky130_fd_sc_hd__mux2_1
X_4997_ _4694_/X _4988_/X _4996_/Y _4964_/X vssd1 vssd1 vccd1 vccd1 _8251_/D sky130_fd_sc_hd__o211a_1
X_3948_ _3948_/A vssd1 vssd1 vccd1 vccd1 _8595_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3448_ clkbuf_0__3448_/X vssd1 vssd1 vccd1 vccd1 _7071__475/A sky130_fd_sc_hd__clkbuf_4
X_3879_ _8201_/Q vssd1 vssd1 vccd1 vccd1 _3983_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8406_ _8406_/CLK _8406_/D vssd1 vssd1 vccd1 vccd1 _8406_/Q sky130_fd_sc_hd__dfxtp_1
X_5618_ _5618_/A vssd1 vssd1 vccd1 vccd1 _8072_/D sky130_fd_sc_hd__clkbuf_1
X_5549_ _8123_/Q _4441_/A _5549_/S vssd1 vssd1 vccd1 vccd1 _5550_/A sky130_fd_sc_hd__mux2_1
X_8337_ _8337_/CLK _8337_/D vssd1 vssd1 vccd1 vccd1 _8337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7142__531 _7144__533/A vssd1 vssd1 vccd1 vccd1 _8340_/CLK sky130_fd_sc_hd__inv_2
X_8268_ _8268_/CLK _8268_/D vssd1 vssd1 vccd1 vccd1 _8268_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3664_ clkbuf_0__3664_/X vssd1 vssd1 vccd1 vccd1 _7728__30/A sky130_fd_sc_hd__clkbuf_4
X_8199_ _8199_/CLK _8199_/D vssd1 vssd1 vccd1 vccd1 _8199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6821__365 _6821__365/A vssd1 vssd1 vccd1 vccd1 _8160_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7004__424 _7005__425/A vssd1 vssd1 vccd1 vccd1 _8230_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8625_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4920_ _4827_/X _4918_/X _4919_/X vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__o21a_1
X_4851_ _7907_/Q _4817_/X _4845_/X _4850_/X vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4782_ _4780_/X _4781_/X _4801_/S vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7570_ _7555_/B _7555_/C _7808_/A vssd1 vssd1 vccd1 vccd1 _7570_/X sky130_fd_sc_hd__a21bo_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7011__428 _7013__430/A vssd1 vssd1 vccd1 vccd1 _8234_/CLK sky130_fd_sc_hd__inv_2
X_6521_ _6521_/A vssd1 vssd1 vccd1 vccd1 _7965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6452_ _6452_/A vssd1 vssd1 vccd1 vccd1 _6452_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5403_ _8194_/Q vssd1 vssd1 vccd1 vccd1 _5598_/A sky130_fd_sc_hd__clkbuf_2
X_8122_ _8122_/CLK _8122_/D vssd1 vssd1 vccd1 vccd1 _8122_/Q sky130_fd_sc_hd__dfxtp_1
X_6383_ _8048_/Q _6403_/A _6382_/X vssd1 vssd1 vccd1 vccd1 _6383_/Y sky130_fd_sc_hd__a21oi_1
X_5334_ _5389_/B _5323_/Y _5326_/Y _5333_/X _5387_/B vssd1 vssd1 vccd1 vccd1 _5335_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_114_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5265_ _5351_/A _5252_/X _5256_/X _5264_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5265_/X
+ sky130_fd_sc_hd__o311a_1
X_8053_ _8608_/CLK _8053_/D vssd1 vssd1 vccd1 vccd1 _8053_/Q sky130_fd_sc_hd__dfxtp_1
X_5196_ _8489_/Q _8473_/Q _8465_/Q _8497_/Q _5324_/S _5101_/X vssd1 vssd1 vccd1 vccd1
+ _5196_/X sky130_fd_sc_hd__mux4_2
X_4216_ _5485_/B _4241_/B vssd1 vssd1 vccd1 vccd1 _4239_/S sky130_fd_sc_hd__nor2_2
X_4147_ _4147_/A vssd1 vssd1 vccd1 vccd1 _8489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7208__84 _7208__84/A vssd1 vssd1 vccd1 vccd1 _8393_/CLK sky130_fd_sc_hd__inv_2
X_4078_ _8511_/Q _3943_/X _4082_/S vssd1 vssd1 vccd1 vccd1 _4079_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7906_ _7906_/CLK _7906_/D vssd1 vssd1 vccd1 vccd1 _7906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7837_ _7837_/A vssd1 vssd1 vccd1 vccd1 _8630_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7768_ _7768_/A vssd1 vssd1 vccd1 vccd1 _8610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6719_ _6719_/A vssd1 vssd1 vccd1 vccd1 _8089_/D sky130_fd_sc_hd__clkbuf_1
X_7699_ _8567_/Q _7687_/X _7698_/X _7684_/A vssd1 vssd1 vccd1 vccd1 _8566_/D sky130_fd_sc_hd__o211a_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6931__382 _6932__383/A vssd1 vssd1 vccd1 vccd1 _8178_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3647_ clkbuf_0__3647_/X vssd1 vssd1 vccd1 vccd1 _7458__133/A sky130_fd_sc_hd__clkbuf_4
X_7521__9 _7521__9/A vssd1 vssd1 vccd1 vccd1 _8523_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6641__283 _6641__283/A vssd1 vssd1 vccd1 vccd1 _8043_/CLK sky130_fd_sc_hd__inv_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__3310_ clkbuf_0__3310_/X vssd1 vssd1 vccd1 vccd1 _6772__330/A sky130_fd_sc_hd__clkbuf_16
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7149__537 _7149__537/A vssd1 vssd1 vccd1 vccd1 _8346_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5050_ _5050_/A vssd1 vssd1 vccd1 vccd1 _8227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4001_ _4001_/A vssd1 vssd1 vccd1 vccd1 _8578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5952_ _7719_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__or2_1
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4903_ _6947_/B vssd1 vssd1 vccd1 vccd1 _4903_/X sky130_fd_sc_hd__clkbuf_2
X_5883_ _5883_/A vssd1 vssd1 vccd1 vccd1 _7860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4834_ _4834_/A vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__clkbuf_2
X_7622_ _7621_/X _7628_/B vssd1 vssd1 vccd1 vccd1 _7623_/A sky130_fd_sc_hd__and2b_1
X_4765_ _4683_/X _4749_/X _4753_/X _4764_/X vssd1 vssd1 vccd1 vccd1 _4765_/X sky130_fd_sc_hd__a31o_2
X_7553_ _7552_/B _7552_/C _7817_/A vssd1 vssd1 vccd1 vccd1 _7553_/Y sky130_fd_sc_hd__a21oi_1
X_6504_ _7958_/Q _6563_/B _6562_/A _6503_/X vssd1 vssd1 vccd1 vccd1 _7958_/D sky130_fd_sc_hd__o211a_1
X_4696_ _4820_/A _4704_/A vssd1 vssd1 vccd1 vccd1 _4834_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _8054_/Q _6403_/X _7055_/B vssd1 vssd1 vccd1 vccd1 _6435_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6366_ _6505_/B _6366_/B _6366_/C _6366_/D vssd1 vssd1 vccd1 vccd1 _7790_/C sky130_fd_sc_hd__or4_1
XFILLER_114_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3078_ clkbuf_0__3078_/X vssd1 vssd1 vccd1 vccd1 _6334__205/A sky130_fd_sc_hd__clkbuf_4
X_5317_ _8392_/Q _5236_/X _5238_/X _8384_/Q _5239_/X vssd1 vssd1 vccd1 vccd1 _5317_/X
+ sky130_fd_sc_hd__o221a_1
X_8105_ _8105_/CLK _8105_/D vssd1 vssd1 vccd1 vccd1 _8105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8036_ _8036_/CLK _8036_/D vssd1 vssd1 vccd1 vccd1 _8036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6297_ _7723_/A _7900_/Q _6297_/S vssd1 vssd1 vccd1 vccd1 _6298_/A sky130_fd_sc_hd__mux2_1
X_6584__237 _6585__238/A vssd1 vssd1 vccd1 vccd1 _7997_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5248_ _5359_/B vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5179_ _5391_/B _5178_/X _5333_/A vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3432_ clkbuf_0__3432_/X vssd1 vssd1 vccd1 vccd1 _6993__415/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6786__341 _6788__343/A vssd1 vssd1 vccd1 vccd1 _8133_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6938__388 _6940__390/A vssd1 vssd1 vccd1 vccd1 _8184_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7202__79 _7203__80/A vssd1 vssd1 vccd1 vccd1 _8388_/CLK sky130_fd_sc_hd__inv_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4450_/X _8319_/Q _4550_/S vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4481_ _8577_/Q vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__buf_2
X_6220_ _6280_/A vssd1 vssd1 vccd1 vccd1 _6647_/A sky130_fd_sc_hd__buf_4
X_6151_ _6136_/X _6148_/X _6150_/X _6139_/X vssd1 vssd1 vccd1 vccd1 _6151_/X sky130_fd_sc_hd__o211a_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5102_ _7927_/Q _8135_/Q _8414_/Q _8162_/Q _5324_/S _5101_/X vssd1 vssd1 vccd1 vccd1
+ _5102_/X sky130_fd_sc_hd__mux4_2
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6101_/A vssd1 vssd1 vccd1 vccd1 _6082_/X sky130_fd_sc_hd__clkbuf_2
X_5033_ _8234_/Q _4528_/X _5035_/S vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__mux2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6984_ _7723_/C vssd1 vssd1 vccd1 vccd1 _7714_/C sky130_fd_sc_hd__clkbuf_1
X_5935_ _5935_/A vssd1 vssd1 vccd1 vccd1 _5935_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5866_ _7910_/Q _5598_/A _5872_/S vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4817_ _4817_/A vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__clkbuf_2
X_7605_ _7603_/A _7667_/B _7683_/A vssd1 vssd1 vccd1 vccd1 _7605_/X sky130_fd_sc_hd__a21bo_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5797_ _5797_/A vssd1 vssd1 vccd1 vccd1 _7989_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3664_ _7542_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3664_/X sky130_fd_sc_hd__clkbuf_16
X_8585_ _8585_/CLK _8585_/D vssd1 vssd1 vccd1 vccd1 _8585_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _4699_/X _4747_/X _4706_/X vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7467_ _7467_/A vssd1 vssd1 vccd1 vccd1 _7467_/X sky130_fd_sc_hd__buf_1
X_4679_ _4684_/B vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6418_ _8629_/Q _6403_/X _6373_/X vssd1 vssd1 vccd1 vccd1 _6422_/B sky130_fd_sc_hd__a21oi_1
X_7398_ _7398_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _8440_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput104 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _6714_/A sky130_fd_sc_hd__buf_6
X_8019_ _8019_/CLK _8019_/D vssd1 vssd1 vccd1 vccd1 _8019_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3415_ clkbuf_0__3415_/X vssd1 vssd1 vccd1 vccd1 _6963__395/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3981_ _3981_/A vssd1 vssd1 vccd1 vccd1 _7757_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0__3481_ clkbuf_0__3481_/X vssd1 vssd1 vccd1 vccd1 _7234__105/A sky130_fd_sc_hd__clkbuf_4
X_5720_ _8023_/Q _5619_/X _5728_/S vssd1 vssd1 vccd1 vccd1 _5721_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8650__215 vssd1 vssd1 vccd1 vccd1 _8650__215/HI core0Index[2] sky130_fd_sc_hd__conb_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7187__67 _7188__68/A vssd1 vssd1 vccd1 vccd1 _8376_/CLK sky130_fd_sc_hd__inv_2
X_5651_ _5601_/X _8061_/Q _5655_/S vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5582_ _5582_/A vssd1 vssd1 vccd1 vccd1 _8109_/D sky130_fd_sc_hd__clkbuf_1
X_8370_ _8370_/CLK _8370_/D vssd1 vssd1 vccd1 vccd1 _8370_/Q sky130_fd_sc_hd__dfxtp_1
X_4602_ _4602_/A vssd1 vssd1 vccd1 vccd1 _8298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4533_ _4533_/A vssd1 vssd1 vccd1 vccd1 _8327_/D sky130_fd_sc_hd__clkbuf_1
X_7321_ _8416_/Q vssd1 vssd1 vccd1 vccd1 _7321_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7252_ _7252_/A _7327_/A _7252_/C vssd1 vssd1 vccd1 vccd1 _7313_/B sky130_fd_sc_hd__and3_1
X_4464_ _4463_/X _8348_/Q _4470_/S vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__mux2_1
X_4395_ _4111_/X _8373_/Q _4401_/S vssd1 vssd1 vccd1 vccd1 _4396_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6134_ _7875_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6134_/X sky130_fd_sc_hd__or2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065_ _8097_/Q _6069_/B vssd1 vssd1 vccd1 vccd1 _6066_/A sky130_fd_sc_hd__and2_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5016_ _8241_/Q _4531_/X _5016_/S vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__mux2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5918_ _6195_/B _5918_/B vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6898_ _8620_/Q _7546_/B vssd1 vssd1 vccd1 vccd1 _7586_/C sky130_fd_sc_hd__xor2_1
XFILLER_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5849_ _5849_/A vssd1 vssd1 vccd1 vccd1 _7918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3647_ _7455_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3647_/X sky130_fd_sc_hd__clkbuf_16
X_8568_ _8568_/CLK _8568_/D vssd1 vssd1 vccd1 vccd1 _8568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8499_ _8499_/CLK _8499_/D vssd1 vssd1 vccd1 vccd1 _8499_/Q sky130_fd_sc_hd__dfxtp_1
X_7106__502 _7109__505/A vssd1 vssd1 vccd1 vccd1 _8311_/CLK sky130_fd_sc_hd__inv_2
X_7497__165 _7497__165/A vssd1 vssd1 vccd1 vccd1 _8504_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6343__212 _6343__212/A vssd1 vssd1 vccd1 vccd1 _7924_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7441__120 _7441__120/A vssd1 vssd1 vccd1 vccd1 _8459_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4180_ _4666_/C _4178_/Y _4179_/X vssd1 vssd1 vccd1 vccd1 _4180_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6799__351 _6799__351/A vssd1 vssd1 vccd1 vccd1 _8143_/CLK sky130_fd_sc_hd__inv_2
X_7870_ _8631_/CLK _7870_/D vssd1 vssd1 vccd1 vccd1 _7870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7092__491 _7094__493/A vssd1 vssd1 vccd1 vccd1 _8300_/CLK sky130_fd_sc_hd__inv_2
X_3964_ _3964_/A vssd1 vssd1 vccd1 vccd1 _8591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5703_ _5703_/A vssd1 vssd1 vccd1 vccd1 _8031_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3464_ clkbuf_0__3464_/X vssd1 vssd1 vccd1 vccd1 _7152__540/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3895_ _8202_/Q _3983_/B _5074_/A vssd1 vssd1 vccd1 vccd1 _3895_/X sky130_fd_sc_hd__a21o_1
X_8422_ _8422_/CLK _8422_/D vssd1 vssd1 vccd1 vccd1 _8422_/Q sky130_fd_sc_hd__dfxtp_1
X_5634_ _8067_/Q _5633_/X _5634_/S vssd1 vssd1 vccd1 vccd1 _5635_/A sky130_fd_sc_hd__mux2_1
X_8353_ _8353_/CLK _8353_/D vssd1 vssd1 vccd1 vccd1 _8353_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3432_ _6988_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3432_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5565_ _5412_/X _8116_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__mux2_1
X_7304_ _7548_/A _7304_/B vssd1 vssd1 vccd1 vccd1 _7304_/Y sky130_fd_sc_hd__nand2_1
X_5496_ _5496_/A vssd1 vssd1 vccd1 vccd1 _8150_/D sky130_fd_sc_hd__clkbuf_1
X_4516_ _8193_/Q vssd1 vssd1 vccd1 vccd1 _4516_/X sky130_fd_sc_hd__clkbuf_4
X_8284_ _8284_/CLK _8284_/D vssd1 vssd1 vccd1 vccd1 _8284_/Q sky130_fd_sc_hd__dfxtp_1
X_4447_ _4447_/A vssd1 vssd1 vccd1 vccd1 _4447_/X sky130_fd_sc_hd__clkbuf_2
X_7235_ _5942_/A _4164_/X _6647_/A vssd1 vssd1 vccd1 vccd1 _7432_/S sky130_fd_sc_hd__a21oi_2
X_7166_ _7479_/A vssd1 vssd1 vccd1 vccd1 _7166_/X sky130_fd_sc_hd__buf_1
X_4378_ _4378_/A vssd1 vssd1 vccd1 vccd1 _8381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6117_ _6136_/A vssd1 vssd1 vccd1 vccd1 _6117_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7097_ _7097_/A vssd1 vssd1 vccd1 vccd1 _7097_/X sky130_fd_sc_hd__buf_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _6048_/A vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _7999_/CLK _7999_/D vssd1 vssd1 vccd1 vccd1 _7999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6679__300 _6679__300/A vssd1 vssd1 vccd1 vccd1 _8068_/CLK sky130_fd_sc_hd__inv_2
X_6605__254 _6606__255/A vssd1 vssd1 vccd1 vccd1 _8014_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5350_ _5305_/A _5348_/X _5349_/X vssd1 vssd1 vccd1 vccd1 _5351_/C sky130_fd_sc_hd__o21a_1
Xoutput205 _6105_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4301_ _4316_/S vssd1 vssd1 vccd1 vccd1 _4310_/S sky130_fd_sc_hd__buf_2
X_6686__304 _6687__305/A vssd1 vssd1 vccd1 vccd1 _8072_/CLK sky130_fd_sc_hd__inv_2
X_5281_ _8393_/Q _5271_/X _5238_/A _8385_/Q _5239_/A vssd1 vssd1 vccd1 vccd1 _5281_/X
+ sky130_fd_sc_hd__o221a_1
X_4232_ _8572_/Q vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__buf_2
X_7020_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7020_/X sky130_fd_sc_hd__buf_1
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4163_ _4259_/A vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4094_ _4094_/A vssd1 vssd1 vccd1 vccd1 _8505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7922_ _7922_/CLK _7922_/D vssd1 vssd1 vccd1 vccd1 _7922_/Q sky130_fd_sc_hd__dfxtp_1
X_8656__221 vssd1 vssd1 vccd1 vccd1 _8656__221/HI core1Index[1] sky130_fd_sc_hd__conb_1
X_7853_ _7853_/CLK _7853_/D vssd1 vssd1 vccd1 vccd1 _7853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6804_ _6714_/A _6492_/C _6804_/S vssd1 vssd1 vccd1 vccd1 _6805_/A sky130_fd_sc_hd__mux2_1
X_7784_ _8615_/Q _7777_/X _7783_/X _6503_/X vssd1 vssd1 vccd1 vccd1 _8615_/D sky130_fd_sc_hd__o211a_1
X_4996_ _4996_/A _4996_/B vssd1 vssd1 vccd1 vccd1 _4996_/Y sky130_fd_sc_hd__nand2_1
X_3947_ _8595_/Q _3946_/X _3950_/S vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__mux2_1
X_6735_ _6735_/A vssd1 vssd1 vccd1 vccd1 _8096_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3447_ clkbuf_0__3447_/X vssd1 vssd1 vccd1 vccd1 _7063__468/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3878_ _8202_/Q vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8405_ _8405_/CLK _8405_/D vssd1 vssd1 vccd1 vccd1 _8405_/Q sky130_fd_sc_hd__dfxtp_1
X_5617_ _5616_/X _8072_/Q _5617_/S vssd1 vssd1 vccd1 vccd1 _5618_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5548_ _5548_/A vssd1 vssd1 vccd1 vccd1 _8124_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3415_ _6941_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3415_/X sky130_fd_sc_hd__clkbuf_16
X_8336_ _8336_/CLK _8336_/D vssd1 vssd1 vccd1 vccd1 _8336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8267_ _8267_/CLK _8267_/D vssd1 vssd1 vccd1 vccd1 _8267_/Q sky130_fd_sc_hd__dfxtp_1
X_5479_ _4444_/X _8157_/Q _5483_/S vssd1 vssd1 vccd1 vccd1 _5480_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8198_ _8198_/CLK _8198_/D vssd1 vssd1 vccd1 vccd1 _8198_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3663_ clkbuf_0__3663_/X vssd1 vssd1 vccd1 vccd1 _7735_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6780__336 _6782__338/A vssd1 vssd1 vccd1 vccd1 _8128_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099__497 _7099__497/A vssd1 vssd1 vccd1 vccd1 _8306_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4850_ _4847_/X _8043_/Q _8027_/Q _4849_/X vssd1 vssd1 vccd1 vccd1 _4850_/X sky130_fd_sc_hd__a22o_1
XFILLER_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4781_ _8230_/Q _8185_/Q _8077_/Q _8422_/Q _4731_/X _4702_/A vssd1 vssd1 vccd1 vccd1
+ _4781_/X sky130_fd_sc_hd__mux4_1
X_6520_ _6028_/A _7965_/Q _6526_/S vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__mux2_1
X_6451_ _6359_/X _6449_/Y _6450_/Y vssd1 vssd1 vccd1 vccd1 _7944_/D sky130_fd_sc_hd__o21ai_1
X_5402_ _5402_/A vssd1 vssd1 vccd1 vccd1 _8187_/D sky130_fd_sc_hd__clkbuf_1
X_6382_ _6396_/A vssd1 vssd1 vccd1 vccd1 _6382_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8121_ _8121_/CLK _8121_/D vssd1 vssd1 vccd1 vccd1 _8121_/Q sky130_fd_sc_hd__dfxtp_1
X_5333_ _5333_/A _5333_/B _5333_/C vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__and3_1
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5264_ _5264_/A _5264_/B _5264_/C vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__or3_1
X_8052_ _8052_/CLK _8052_/D vssd1 vssd1 vccd1 vccd1 _8052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4215_ _8577_/Q vssd1 vssd1 vccd1 vccd1 _4215_/X sky130_fd_sc_hd__clkbuf_2
X_5195_ _3962_/X _5078_/X _5194_/X _5152_/X vssd1 vssd1 vccd1 vccd1 _8212_/D sky130_fd_sc_hd__o211a_1
X_4146_ _8489_/Q _3937_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__mux2_1
X_7454__130 _7454__130/A vssd1 vssd1 vccd1 vccd1 _8469_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4077_/A vssd1 vssd1 vccd1 vccd1 _8512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7905_ _7905_/CLK _7905_/D vssd1 vssd1 vccd1 vccd1 _7905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7836_ _7836_/A _7836_/B _7836_/C vssd1 vssd1 vccd1 vccd1 _7837_/A sky130_fd_sc_hd__and3_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _4979_/A _4986_/B vssd1 vssd1 vccd1 vccd1 _4984_/A sky130_fd_sc_hd__nor2_1
X_7767_ _7771_/A _8604_/Q vssd1 vssd1 vccd1 vccd1 _7768_/A sky130_fd_sc_hd__and2_1
X_6718_ _5978_/A _8089_/Q _6724_/S vssd1 vssd1 vccd1 vccd1 _6719_/A sky130_fd_sc_hd__mux2_1
X_7698_ _8566_/Q _7698_/B vssd1 vssd1 vccd1 vccd1 _7698_/X sky130_fd_sc_hd__or2_1
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6649_ _8261_/Q _8249_/D vssd1 vssd1 vccd1 vccd1 _6650_/A sky130_fd_sc_hd__and2_1
X_8319_ _8319_/CLK _8319_/D vssd1 vssd1 vccd1 vccd1 _8319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3646_ clkbuf_0__3646_/X vssd1 vssd1 vccd1 vccd1 _7454__130/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4000_ _3977_/X _8578_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _4001_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _6008_/B vssd1 vssd1 vccd1 vccd1 _5960_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_80_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ _4671_/X _8263_/Q _4741_/X _4901_/X vssd1 vssd1 vccd1 vccd1 _4902_/X sky130_fd_sc_hd__a211o_1
X_5882_ _4156_/X _7860_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4833_ _4865_/A vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__buf_2
X_7621_ _7619_/Y _7620_/X _7604_/X _7564_/B vssd1 vssd1 vccd1 vccd1 _7621_/X sky130_fd_sc_hd__o22a_1
X_4764_ _4735_/X _4756_/X _4762_/X _4990_/B vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__o211a_1
X_7552_ _8625_/Q _7552_/B _7552_/C vssd1 vssd1 vccd1 vccd1 _7552_/X sky130_fd_sc_hd__and3_1
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6503_ _7771_/A vssd1 vssd1 vccd1 vccd1 _6503_/X sky130_fd_sc_hd__buf_2
X_4695_ _8179_/Q _8171_/Q _7999_/Q _8240_/Q _4691_/X _4694_/X vssd1 vssd1 vccd1 vccd1
+ _4695_/X sky130_fd_sc_hd__mux4_1
X_6434_ _6474_/A vssd1 vssd1 vccd1 vccd1 _6452_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6365_ _7960_/Q vssd1 vssd1 vccd1 vccd1 _7790_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3077_ clkbuf_0__3077_/X vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__clkbuf_4
X_8104_ _8104_/CLK _8104_/D vssd1 vssd1 vccd1 vccd1 _8104_/Q sky130_fd_sc_hd__dfxtp_1
X_5316_ _8368_/Q _8376_/Q _5352_/S vssd1 vssd1 vccd1 vccd1 _5316_/X sky130_fd_sc_hd__mux2_1
X_6296_ _6296_/A vssd1 vssd1 vccd1 vccd1 _7899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5247_ _5247_/A _5247_/B vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__or2_1
X_8035_ _8035_/CLK _8035_/D vssd1 vssd1 vccd1 vccd1 _8035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _8522_/Q _8514_/Q _7917_/Q _8530_/Q _5122_/X _5123_/X vssd1 vssd1 vccd1 vccd1
+ _5178_/X sky130_fd_sc_hd__mux4_1
X_6996__417 _6997__418/A vssd1 vssd1 vccd1 vccd1 _8223_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4129_ _4129_/A vssd1 vssd1 vccd1 vccd1 _8495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7819_ _7817_/Y _7818_/Y _6391_/X vssd1 vssd1 vccd1 vccd1 _8625_/D sky130_fd_sc_hd__a21oi_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7155__542 _7157__544/A vssd1 vssd1 vccd1 vccd1 _8351_/CLK sky130_fd_sc_hd__inv_2
X_7199__76 _7200__77/A vssd1 vssd1 vccd1 vccd1 _8385_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _8343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6150_ _7879_/Q _6175_/A vssd1 vssd1 vccd1 vccd1 _6150_/X sky130_fd_sc_hd__or2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5101_ _5101_/A vssd1 vssd1 vccd1 vccd1 _5101_/X sky130_fd_sc_hd__buf_4
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6173_/A vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__clkbuf_8
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5032_ _5032_/A vssd1 vssd1 vccd1 vccd1 _8235_/D sky130_fd_sc_hd__clkbuf_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8270_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6983_ _6986_/B _6983_/B vssd1 vssd1 vccd1 vccd1 _7723_/C sky130_fd_sc_hd__and2_1
X_5934_ _6714_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__and2_1
X_7056__462 _7058__464/A vssd1 vssd1 vccd1 vccd1 _8271_/CLK sky130_fd_sc_hd__inv_2
X_5865_ _5865_/A vssd1 vssd1 vccd1 vccd1 _7911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3663_ _7541_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3663_/X sky130_fd_sc_hd__clkbuf_16
X_4816_ _4856_/A vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__buf_2
X_7604_ _7647_/A vssd1 vssd1 vccd1 vccd1 _7604_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5796_ _7989_/Q _5601_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5797_/A sky130_fd_sc_hd__mux2_1
X_8584_ _8584_/CLK _8584_/D vssd1 vssd1 vccd1 vccd1 _8584_/Q sky130_fd_sc_hd__dfxtp_1
X_4747_ _8223_/Q _8110_/Q _8006_/Q _7990_/Q _4700_/X _4714_/X vssd1 vssd1 vccd1 vccd1
+ _4747_/X sky130_fd_sc_hd__mux4_1
X_7535_ _7535_/A vssd1 vssd1 vccd1 vccd1 _7535_/X sky130_fd_sc_hd__buf_1
XFILLER_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6590__242 _6591__243/A vssd1 vssd1 vccd1 vccd1 _8002_/CLK sky130_fd_sc_hd__inv_2
X_4678_ _8251_/Q _4806_/B vssd1 vssd1 vccd1 vccd1 _4684_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7397_ _8440_/Q _7384_/A _7360_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7398_/B sky130_fd_sc_hd__o2bb2a_1
X_6417_ _7939_/Q _6410_/X _6416_/Y _6391_/X vssd1 vssd1 vccd1 vccd1 _7939_/D sky130_fd_sc_hd__a211o_1
XFILLER_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7024__439 _7025__440/A vssd1 vssd1 vccd1 vccd1 _8245_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput105 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _6732_/A sky130_fd_sc_hd__clkbuf_8
X_6279_ _8103_/Q _6222_/X _6236_/A _6247_/A _7892_/Q vssd1 vssd1 vccd1 vccd1 _7892_/D
+ sky130_fd_sc_hd__o32a_1
X_8018_ _8018_/CLK _8018_/D vssd1 vssd1 vccd1 vccd1 _8018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3414_ clkbuf_0__3414_/X vssd1 vssd1 vccd1 vccd1 _6937__387/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3276_ clkbuf_0__3276_/X vssd1 vssd1 vccd1 vccd1 _6753__315/A sky130_fd_sc_hd__clkbuf_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8636__252 vssd1 vssd1 vccd1 vccd1 partID[2] _8636__252/LO sky130_fd_sc_hd__conb_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _8215_/Q vssd1 vssd1 vccd1 vccd1 _5147_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3480_ clkbuf_0__3480_/X vssd1 vssd1 vccd1 vccd1 _7436_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5650_ _5650_/A vssd1 vssd1 vccd1 vccd1 _8062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _4469_/X _8298_/Q _4601_/S vssd1 vssd1 vccd1 vccd1 _4602_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5581_ _5408_/X _8109_/Q _5585_/S vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__mux2_1
X_4532_ _8327_/Q _4531_/X _4532_/S vssd1 vssd1 vccd1 vccd1 _4533_/A sky130_fd_sc_hd__mux2_1
X_7320_ _7320_/A vssd1 vssd1 vccd1 vccd1 _8415_/D sky130_fd_sc_hd__clkbuf_1
X_7251_ _8619_/Q _7394_/A _7394_/B vssd1 vssd1 vccd1 vccd1 _7252_/C sky130_fd_sc_hd__nand3b_1
X_4463_ _8193_/Q vssd1 vssd1 vccd1 vccd1 _4463_/X sky130_fd_sc_hd__buf_4
XFILLER_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4394_ _4394_/A vssd1 vssd1 vccd1 vccd1 _8374_/D sky130_fd_sc_hd__clkbuf_1
X_6133_ _7950_/Q input8/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6133_/X sky130_fd_sc_hd__mux2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6064_/A vssd1 vssd1 vccd1 vccd1 _6064_/X sky130_fd_sc_hd__clkbuf_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _8242_/D sky130_fd_sc_hd__clkbuf_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5917_ _8102_/Q _8103_/Q _8100_/Q _8101_/Q vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__and4bb_2
X_6897_ _8556_/Q _6903_/D vssd1 vssd1 vccd1 vccd1 _7546_/B sky130_fd_sc_hd__xnor2_4
X_5848_ _4432_/X _7918_/Q _5854_/S vssd1 vssd1 vccd1 vccd1 _5849_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3646_ _7449_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3646_/X sky130_fd_sc_hd__clkbuf_16
X_5779_ _5779_/A vssd1 vssd1 vccd1 vccd1 _7997_/D sky130_fd_sc_hd__clkbuf_1
X_8567_ _8568_/CLK _8567_/D vssd1 vssd1 vccd1 vccd1 _8567_/Q sky130_fd_sc_hd__dfxtp_1
X_7740__40 _7740__40/A vssd1 vssd1 vccd1 vccd1 _8591_/CLK sky130_fd_sc_hd__inv_2
X_8498_ _8498_/CLK _8498_/D vssd1 vssd1 vccd1 vccd1 _8498_/Q sky130_fd_sc_hd__dfxtp_1
X_7449_ _7473_/A vssd1 vssd1 vccd1 vccd1 _7449_/X sky130_fd_sc_hd__buf_1
XFILLER_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8673__238 vssd1 vssd1 vccd1 vccd1 _8673__238/HI manufacturerID[10] sky130_fd_sc_hd__conb_1
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3259_ clkbuf_0__3259_/X vssd1 vssd1 vccd1 vccd1 _6641__283/A sky130_fd_sc_hd__clkbuf_4
X_6597__248 _6599__250/A vssd1 vssd1 vccd1 vccd1 _8008_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7192__71 _7194__73/A vssd1 vssd1 vccd1 vccd1 _8380_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ _3962_/X _8591_/Q _3969_/S vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5702_ _5593_/X _8031_/Q _5710_/S vssd1 vssd1 vccd1 vccd1 _5703_/A sky130_fd_sc_hd__mux2_1
X_6682_ _6760_/A vssd1 vssd1 vccd1 vccd1 _6682_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3463_ clkbuf_0__3463_/X vssd1 vssd1 vccd1 vccd1 _7146__535/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3894_ _8203_/Q _8198_/Q vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_8421_ _8421_/CLK _8421_/D vssd1 vssd1 vccd1 vccd1 _8421_/Q sky130_fd_sc_hd__dfxtp_1
X_5633_ _8191_/Q vssd1 vssd1 vccd1 vccd1 _5633_/X sky130_fd_sc_hd__buf_2
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5564_ _5564_/A vssd1 vssd1 vccd1 vccd1 _8117_/D sky130_fd_sc_hd__clkbuf_1
X_8352_ _8352_/CLK _8352_/D vssd1 vssd1 vccd1 vccd1 _8352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4515_ _4515_/A vssd1 vssd1 vccd1 vccd1 _8333_/D sky130_fd_sc_hd__clkbuf_1
X_7303_ _7303_/A _7303_/B vssd1 vssd1 vccd1 vccd1 _7304_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5495_ _8150_/Q _4495_/X _5495_/S vssd1 vssd1 vccd1 vccd1 _5496_/A sky130_fd_sc_hd__mux2_1
X_8283_ _8283_/CLK _8283_/D vssd1 vssd1 vccd1 vccd1 _8283_/Q sky130_fd_sc_hd__dfxtp_1
X_4446_ _4446_/A vssd1 vssd1 vccd1 vccd1 _8353_/D sky130_fd_sc_hd__clkbuf_1
X_4377_ _8381_/Q _4220_/X _4383_/S vssd1 vssd1 vccd1 vccd1 _4378_/A sky130_fd_sc_hd__mux2_1
X_7165_ _7165_/A vssd1 vssd1 vccd1 vccd1 _7165_/X sky130_fd_sc_hd__buf_1
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6116_ _6098_/X _6114_/X _6115_/X _6101_/X vssd1 vssd1 vccd1 vccd1 _6116_/X sky130_fd_sc_hd__o211a_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _8089_/Q _6047_/B vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__and2_1
XFILLER_27_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7101__499 _7102__500/A vssd1 vssd1 vccd1 vccd1 _8308_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ _7998_/CLK _7998_/D vssd1 vssd1 vccd1 vccd1 _7998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6949_ _7053_/C vssd1 vssd1 vccd1 vccd1 _6958_/B sky130_fd_sc_hd__clkbuf_1
X_8619_ _8623_/CLK _8619_/D vssd1 vssd1 vccd1 vccd1 _8619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6969__400 _6969__400/A vssd1 vssd1 vccd1 vccd1 _8204_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput206 _6108_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4300_ _5539_/B _5826_/B vssd1 vssd1 vccd1 vccd1 _4316_/S sky130_fd_sc_hd__nor2_2
X_5280_ _8369_/Q _8377_/Q _5345_/S vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _4231_/A vssd1 vssd1 vccd1 vccd1 _8472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _8255_/Q vssd1 vssd1 vccd1 vccd1 _4259_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4093_ _8505_/Q _3937_/X _4095_/S vssd1 vssd1 vccd1 vccd1 _4094_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7921_ _7921_/CLK _7921_/D vssd1 vssd1 vccd1 vccd1 _7921_/Q sky130_fd_sc_hd__dfxtp_1
X_7852_ _7852_/CLK _7852_/D vssd1 vssd1 vccd1 vccd1 _7852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6803_ _6803_/A vssd1 vssd1 vccd1 vccd1 _8145_/D sky130_fd_sc_hd__clkbuf_1
X_7783_ _5980_/A _7778_/X _7777_/A vssd1 vssd1 vccd1 vccd1 _7783_/X sky130_fd_sc_hd__a21bo_1
X_4995_ _4815_/X _4988_/X _4994_/Y _4964_/X vssd1 vssd1 vccd1 vccd1 _8252_/D sky130_fd_sc_hd__o211a_1
X_3946_ _8571_/Q vssd1 vssd1 vccd1 vccd1 _3946_/X sky130_fd_sc_hd__buf_2
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6734_ _8096_/Q _5993_/A _6742_/S vssd1 vssd1 vccd1 vccd1 _6735_/A sky130_fd_sc_hd__mux2_1
X_8404_ _8404_/CLK _8404_/D vssd1 vssd1 vccd1 vccd1 _8404_/Q sky130_fd_sc_hd__dfxtp_1
X_3877_ _5376_/A _3877_/B vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__or2_4
X_5616_ _5616_/A vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5547_ _8124_/Q _4438_/A _5549_/S vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3414_ _6935_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3414_/X sky130_fd_sc_hd__clkbuf_16
X_8335_ _8335_/CLK _8335_/D vssd1 vssd1 vccd1 vccd1 _8335_/Q sky130_fd_sc_hd__dfxtp_1
X_5478_ _5478_/A vssd1 vssd1 vccd1 vccd1 _8158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8266_ _8266_/CLK _8266_/D vssd1 vssd1 vccd1 vccd1 _8266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4429_ _4451_/S vssd1 vssd1 vccd1 vccd1 _4442_/S sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3276_ _6694_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3276_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3662_ clkbuf_0__3662_/X vssd1 vssd1 vccd1 vccd1 _7537__22/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8197_ _8197_/CLK _8197_/D vssd1 vssd1 vccd1 vccd1 _8197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7079_ _7079_/A vssd1 vssd1 vccd1 vccd1 _7079_/X sky130_fd_sc_hd__buf_1
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8679__244 vssd1 vssd1 vccd1 vccd1 _8679__244/HI partID[12] sky130_fd_sc_hd__conb_1
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7119__513 _7119__513/A vssd1 vssd1 vccd1 vccd1 _8322_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _8332_/Q _8117_/Q _8069_/Q _8021_/Q _4731_/X _4729_/X vssd1 vssd1 vccd1 vccd1
+ _4780_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6450_ _7944_/Q _6416_/A _6265_/X vssd1 vssd1 vccd1 vccd1 _6450_/Y sky130_fd_sc_hd__a21oi_1
X_5401_ _5398_/X _8187_/Q _5417_/S vssd1 vssd1 vccd1 vccd1 _5402_/A sky130_fd_sc_hd__mux2_1
X_6356__223 _6356__223/A vssd1 vssd1 vccd1 vccd1 _7935_/CLK sky130_fd_sc_hd__inv_2
X_6381_ _6433_/B _6381_/B vssd1 vssd1 vccd1 vccd1 _6396_/A sky130_fd_sc_hd__or2_1
X_8120_ _8120_/CLK _8120_/D vssd1 vssd1 vccd1 vccd1 _8120_/Q sky130_fd_sc_hd__dfxtp_1
X_5332_ _5274_/X _5330_/X _5331_/X vssd1 vssd1 vccd1 vccd1 _5333_/C sky130_fd_sc_hd__o21ai_1
XFILLER_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5263_ _5294_/A _5261_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _5264_/C sky130_fd_sc_hd__o21a_1
X_8051_ _8608_/CLK _8051_/D vssd1 vssd1 vccd1 vccd1 _8051_/Q sky130_fd_sc_hd__dfxtp_1
X_4214_ _4214_/A vssd1 vssd1 vccd1 vccd1 _8477_/D sky130_fd_sc_hd__clkbuf_1
X_5194_ _8212_/Q _5080_/X _5385_/A _5193_/X _5148_/X vssd1 vssd1 vccd1 vccd1 _5194_/X
+ sky130_fd_sc_hd__a221o_1
X_4145_ _4145_/A vssd1 vssd1 vccd1 vccd1 _8490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4076_ _8512_/Q _3940_/X _4076_/S vssd1 vssd1 vccd1 vccd1 _4077_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7904_ _7904_/CLK _7904_/D vssd1 vssd1 vccd1 vccd1 _7904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7835_ _7714_/A _7778_/A _7826_/A vssd1 vssd1 vccd1 vccd1 _7836_/C sky130_fd_sc_hd__a21o_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7526__13 _7526__13/A vssd1 vssd1 vccd1 vccd1 _8527_/CLK sky130_fd_sc_hd__inv_2
X_4978_ _4985_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4986_/B sky130_fd_sc_hd__nand2_1
X_7766_ _7766_/A vssd1 vssd1 vccd1 vccd1 _8609_/D sky130_fd_sc_hd__clkbuf_1
X_3929_ _8601_/Q _3872_/X _3941_/S vssd1 vssd1 vccd1 vccd1 _3930_/A sky130_fd_sc_hd__mux2_1
X_6717_ _6717_/A vssd1 vssd1 vccd1 vccd1 _8088_/D sky130_fd_sc_hd__clkbuf_1
X_7697_ _8566_/Q _7687_/X _7696_/X _7684_/X vssd1 vssd1 vccd1 vccd1 _8565_/D sky130_fd_sc_hd__o211a_1
XFILLER_109_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6648_ _6663_/B vssd1 vssd1 vccd1 vccd1 _8249_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8318_ _8318_/CLK _8318_/D vssd1 vssd1 vccd1 vccd1 _8318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8249_ _8608_/CLK _8249_/D vssd1 vssd1 vccd1 vccd1 _8249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3645_ clkbuf_0__3645_/X vssd1 vssd1 vccd1 vccd1 _7473_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3259_ _6638_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3259_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7214__89 _7214__89/A vssd1 vssd1 vccd1 vccd1 _8398_/CLK sky130_fd_sc_hd__inv_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5950_ _5950_/A vssd1 vssd1 vccd1 vccd1 _5950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4901_ _4887_/X _4900_/X _4989_/A vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__o21a_1
X_5881_ _5896_/S vssd1 vssd1 vccd1 vccd1 _5890_/S sky130_fd_sc_hd__buf_2
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7620_ _7642_/A vssd1 vssd1 vccd1 vccd1 _7620_/X sky130_fd_sc_hd__clkbuf_2
X_4832_ _4856_/A vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4763_ _4763_/A vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__clkbuf_4
X_7551_ _7551_/A _7551_/B vssd1 vssd1 vccd1 vccd1 _7551_/Y sky130_fd_sc_hd__nand2_1
X_4694_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__buf_4
X_6502_ _7760_/A vssd1 vssd1 vccd1 vccd1 _7771_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6618__265 _6618__265/A vssd1 vssd1 vccd1 vccd1 _8025_/CLK sky130_fd_sc_hd__inv_2
X_6433_ _6433_/A _6433_/B vssd1 vssd1 vccd1 vccd1 _6474_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6364_ _7961_/Q _7962_/Q _6376_/B vssd1 vssd1 vccd1 vccd1 _6433_/A sky130_fd_sc_hd__or3_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3076_ clkbuf_0__3076_/X vssd1 vssd1 vccd1 vccd1 _6325__198/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5315_ _5233_/X _5313_/X _5314_/X vssd1 vssd1 vccd1 vccd1 _5315_/Y sky130_fd_sc_hd__o21ai_1
X_6295_ _7828_/A _7899_/Q _6297_/S vssd1 vssd1 vccd1 vccd1 _6296_/A sky130_fd_sc_hd__mux2_1
X_8103_ _8569_/CLK _8103_/D vssd1 vssd1 vccd1 vccd1 _8103_/Q sky130_fd_sc_hd__dfxtp_1
X_5246_ _5244_/X _5245_/X _5246_/S vssd1 vssd1 vccd1 vccd1 _5247_/B sky130_fd_sc_hd__mux2_1
X_8034_ _8034_/CLK _8034_/D vssd1 vssd1 vccd1 vccd1 _8034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177_ _8490_/Q _8474_/Q _8466_/Q _8498_/Q _5324_/S _5101_/X vssd1 vssd1 vccd1 vccd1
+ _5177_/X sky130_fd_sc_hd__mux4_2
XFILLER_96_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _4127_/X _8495_/Q _4136_/S vssd1 vssd1 vccd1 vccd1 _4129_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4059_ _4059_/A vssd1 vssd1 vccd1 vccd1 _8519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _7818_/A _7818_/B vssd1 vssd1 vccd1 vccd1 _7818_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6793__347 _6794__348/A vssd1 vssd1 vccd1 vccd1 _8139_/CLK sky130_fd_sc_hd__inv_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5100_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5101_/A sky130_fd_sc_hd__clkbuf_2
X_6080_ _6080_/A vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__buf_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5031_ _8235_/Q _4525_/X _5035_/S vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__mux2_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6014_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5864_ _7911_/Q _5593_/A _5872_/S vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3662_ _7535_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3662_/X sky130_fd_sc_hd__clkbuf_16
X_4815_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4815_/X sky130_fd_sc_hd__clkbuf_4
X_7603_ _7603_/A vssd1 vssd1 vccd1 vccd1 _7603_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8583_ _8583_/CLK _8583_/D vssd1 vssd1 vccd1 vccd1 _8583_/Q sky130_fd_sc_hd__dfxtp_2
X_5795_ _5795_/A vssd1 vssd1 vccd1 vccd1 _7990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4746_ _8178_/Q _8170_/Q _7998_/Q _8239_/Q _4691_/X _4694_/X vssd1 vssd1 vccd1 vccd1
+ _4746_/X sky130_fd_sc_hd__mux4_1
X_4677_ _8250_/Q vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__clkbuf_4
X_7396_ _7398_/A _7396_/B vssd1 vssd1 vccd1 vccd1 _8439_/D sky130_fd_sc_hd__nor2_1
X_6416_ _6416_/A _6416_/B _6416_/C vssd1 vssd1 vccd1 vccd1 _6416_/Y sky130_fd_sc_hd__nor3_1
X_6347_ _6353_/A vssd1 vssd1 vccd1 vccd1 _6347_/X sky130_fd_sc_hd__buf_1
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput106 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _6505_/A sky130_fd_sc_hd__buf_8
X_6278_ _8102_/Q _6222_/X _6236_/A _6247_/A _7891_/Q vssd1 vssd1 vccd1 vccd1 _7891_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_102_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8017_ _8017_/CLK _8017_/D vssd1 vssd1 vccd1 vccd1 _8017_/Q sky130_fd_sc_hd__dfxtp_1
X_5229_ _5359_/B vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0__3413_ clkbuf_0__3413_/X vssd1 vssd1 vccd1 vccd1 _6934__385/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6690__307/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6197_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6207__181 _6209__183/A vssd1 vssd1 vccd1 vccd1 _7850_/CLK sky130_fd_sc_hd__inv_2
X_4600_ _4600_/A vssd1 vssd1 vccd1 vccd1 _8299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5580_ _5580_/A vssd1 vssd1 vccd1 vccd1 _8110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4531_ _8188_/Q vssd1 vssd1 vccd1 vccd1 _4531_/X sky130_fd_sc_hd__buf_2
XFILLER_116_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4462_ _4462_/A vssd1 vssd1 vccd1 vccd1 _8349_/D sky130_fd_sc_hd__clkbuf_1
X_7250_ _8620_/Q _7250_/B vssd1 vssd1 vccd1 vccd1 _7327_/A sky130_fd_sc_hd__xor2_1
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4393_ _4104_/X _8374_/Q _4401_/S vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6132_ _6117_/X _6129_/X _6131_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6132_/X sky130_fd_sc_hd__o211a_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6063_ _8096_/Q _6069_/B vssd1 vssd1 vccd1 vccd1 _6064_/A sky130_fd_sc_hd__and2_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5014_ _8242_/Q _4528_/X _5016_/S vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__mux2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5916_ _5916_/A vssd1 vssd1 vccd1 vccd1 _6195_/B sky130_fd_sc_hd__clkbuf_4
X_6896_ _7811_/A _7589_/B _7590_/B _7814_/A _6895_/X vssd1 vssd1 vccd1 vccd1 _6896_/Y
+ sky130_fd_sc_hd__o221ai_1
X_5847_ _5847_/A vssd1 vssd1 vccd1 vccd1 _7919_/D sky130_fd_sc_hd__clkbuf_1
X_5778_ _7997_/Q _5601_/A _5782_/S vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3645_ _7448_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3645_/X sky130_fd_sc_hd__clkbuf_16
X_6817__361 _6819__363/A vssd1 vssd1 vccd1 vccd1 _8156_/CLK sky130_fd_sc_hd__inv_2
X_8566_ _8568_/CLK _8566_/D vssd1 vssd1 vccd1 vccd1 _8566_/Q sky130_fd_sc_hd__dfxtp_1
X_7030__444 _7031__445/A vssd1 vssd1 vccd1 vccd1 _8251_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4729_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__buf_2
X_8497_ _8497_/CLK _8497_/D vssd1 vssd1 vccd1 vccd1 _8497_/Q sky130_fd_sc_hd__dfxtp_1
X_7517_ _7529_/A vssd1 vssd1 vccd1 vccd1 _7517_/X sky130_fd_sc_hd__buf_1
X_7448_ _7448_/A vssd1 vssd1 vccd1 vccd1 _7448_/X sky130_fd_sc_hd__buf_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7379_ _7379_/A _7379_/B vssd1 vssd1 vccd1 vccd1 _7379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _6935_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3258_ clkbuf_0__3258_/X vssd1 vssd1 vccd1 vccd1 _6637__280/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7113__508 _7115__510/A vssd1 vssd1 vccd1 vccd1 _8317_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6350__218 _6351__219/A vssd1 vssd1 vccd1 vccd1 _7930_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5701_ _5716_/S vssd1 vssd1 vccd1 vccd1 _5710_/S sky130_fd_sc_hd__buf_2
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ _8575_/Q vssd1 vssd1 vccd1 vccd1 _3962_/X sky130_fd_sc_hd__buf_2
X_6681_ _6797_/A vssd1 vssd1 vccd1 vccd1 _6681_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3462_ clkbuf_0__3462_/X vssd1 vssd1 vccd1 vccd1 _7140__530/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3893_ _3893_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _3893_/Y sky130_fd_sc_hd__nor2_1
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _8068_/D sky130_fd_sc_hd__clkbuf_1
X_8420_ _8420_/CLK _8420_/D vssd1 vssd1 vccd1 vccd1 _8420_/Q sky130_fd_sc_hd__dfxtp_1
X_5563_ _5408_/X _8117_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5564_/A sky130_fd_sc_hd__mux2_1
X_8351_ _8351_/CLK _8351_/D vssd1 vssd1 vccd1 vccd1 _8351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4514_ _8333_/Q _4513_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__mux2_1
X_7302_ _7266_/A _7280_/C _7308_/C _8437_/Q vssd1 vssd1 vccd1 vccd1 _7303_/B sky130_fd_sc_hd__a31o_1
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5494_ _5494_/A vssd1 vssd1 vccd1 vccd1 _8151_/D sky130_fd_sc_hd__clkbuf_1
X_8282_ _8282_/CLK _8282_/D vssd1 vssd1 vccd1 vccd1 _8282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4445_ _4444_/X _8353_/Q _4451_/S vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__mux2_1
X_4376_ _4376_/A vssd1 vssd1 vccd1 vccd1 _8382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6115_ _7870_/Q _6126_/B vssd1 vssd1 vccd1 vccd1 _6115_/X sky130_fd_sc_hd__or2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6046_/A vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__clkbuf_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _7997_/CLK _7997_/D vssd1 vssd1 vccd1 vccd1 _7997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6948_ _6948_/A vssd1 vssd1 vccd1 vccd1 _8190_/D sky130_fd_sc_hd__clkbuf_1
X_6879_ _7610_/A _7607_/A _7603_/A _8546_/Q vssd1 vssd1 vccd1 vccd1 _6880_/B sky130_fd_sc_hd__a31o_1
X_8618_ _8622_/CLK _8618_/D vssd1 vssd1 vccd1 vccd1 _8618_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6750__312 _6753__315/A vssd1 vssd1 vccd1 vccd1 _8104_/CLK sky130_fd_sc_hd__inv_2
X_8549_ _8630_/CLK _8549_/D vssd1 vssd1 vccd1 vccd1 _8549_/Q sky130_fd_sc_hd__dfxtp_1
X_7069__473 _7069__473/A vssd1 vssd1 vccd1 vccd1 _8282_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6976__405 _6976__405/A vssd1 vssd1 vccd1 vccd1 _8209_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput207 _6113_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_114_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _8472_/Q _4229_/X _4230_/S vssd1 vssd1 vccd1 vccd1 _4231_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4161_ _8256_/Q vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ _4092_/A vssd1 vssd1 vccd1 vccd1 _8506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7920_ _7920_/CLK _7920_/D vssd1 vssd1 vccd1 vccd1 _7920_/Q sky130_fd_sc_hd__dfxtp_1
X_7851_ _7851_/CLK _7851_/D vssd1 vssd1 vccd1 vccd1 _7851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6802_ _6696_/A _6469_/C _6804_/S vssd1 vssd1 vccd1 vccd1 _6803_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7782_ _8614_/Q _7777_/X _7781_/X _6503_/X vssd1 vssd1 vccd1 vccd1 _8614_/D sky130_fd_sc_hd__o211a_1
X_4994_ _4996_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _4994_/Y sky130_fd_sc_hd__nand2_1
X_3945_ _3945_/A vssd1 vssd1 vccd1 vccd1 _8596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6733_ _6748_/S vssd1 vssd1 vccd1 vccd1 _6742_/S sky130_fd_sc_hd__clkbuf_2
X_6664_ _6664_/A vssd1 vssd1 vccd1 vccd1 _8055_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3445_ clkbuf_0__3445_/X vssd1 vssd1 vccd1 vccd1 _7059__465/A sky130_fd_sc_hd__clkbuf_4
X_8403_ _8403_/CLK _8403_/D vssd1 vssd1 vccd1 vccd1 _8403_/Q sky130_fd_sc_hd__dfxtp_1
X_5615_ _5615_/A vssd1 vssd1 vccd1 vccd1 _8073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3876_ _4336_/A _8204_/Q vssd1 vssd1 vccd1 vccd1 _3877_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8334_ _8334_/CLK _8334_/D vssd1 vssd1 vccd1 vccd1 _8334_/Q sky130_fd_sc_hd__dfxtp_1
X_5546_ _5546_/A vssd1 vssd1 vccd1 vccd1 _8125_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3413_ _6929_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3413_/X sky130_fd_sc_hd__clkbuf_16
X_5477_ _4441_/X _8158_/Q _5477_/S vssd1 vssd1 vccd1 vccd1 _5478_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8265_ _8265_/CLK _8265_/D vssd1 vssd1 vccd1 vccd1 _8265_/Q sky130_fd_sc_hd__dfxtp_1
X_7216_ _7222_/A vssd1 vssd1 vccd1 vccd1 _7216_/X sky130_fd_sc_hd__buf_1
X_4428_ _4573_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _4451_/S sky130_fd_sc_hd__or2_2
Xclkbuf_1_0_0__3661_ clkbuf_0__3661_/X vssd1 vssd1 vccd1 vccd1 _7532__18/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3275_ _6688_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3275_/X sky130_fd_sc_hd__clkbuf_16
X_8196_ _8196_/CLK _8196_/D vssd1 vssd1 vccd1 vccd1 _8196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _4111_/X _8389_/Q _4365_/S vssd1 vssd1 vccd1 vccd1 _4360_/A sky130_fd_sc_hd__mux2_1
X_7147_ _7147_/A vssd1 vssd1 vccd1 vccd1 _7147_/X sky130_fd_sc_hd__buf_1
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _6029_/A vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8577_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7043__454 _7044__455/A vssd1 vssd1 vccd1 vccd1 _8261_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_90 _6088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6757__318 _6758__319/A vssd1 vssd1 vccd1 vccd1 _8110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5400_ _5429_/S vssd1 vssd1 vccd1 vccd1 _5417_/S sky130_fd_sc_hd__clkbuf_4
X_6380_ _6501_/B _6499_/B _6384_/B vssd1 vssd1 vccd1 vccd1 _6436_/B sky130_fd_sc_hd__o21ai_2
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5331_ _5254_/X _8156_/Q _7921_/Q _5257_/X _5135_/A vssd1 vssd1 vccd1 vccd1 _5331_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8050_ _8608_/CLK _8050_/D vssd1 vssd1 vccd1 vccd1 _8050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5262_ _5271_/A _8158_/Q _7923_/Q _5359_/B _5134_/A vssd1 vssd1 vccd1 vccd1 _5262_/X
+ sky130_fd_sc_hd__o221a_1
X_5193_ _5087_/X _5180_/X _5184_/X _5192_/X vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__a31o_2
X_4213_ _8477_/Q _4212_/X _4213_/S vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4144_ _8490_/Q _3934_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4075_ _4075_/A vssd1 vssd1 vccd1 vccd1 _8513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7903_ _8568_/CLK _7903_/D vssd1 vssd1 vccd1 vccd1 _7903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7834_ _7834_/A _7842_/C vssd1 vssd1 vccd1 vccd1 _7836_/B sky130_fd_sc_hd__or2_1
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7765_ _7771_/A _8603_/Q vssd1 vssd1 vccd1 vccd1 _7766_/A sky130_fd_sc_hd__and2_1
XFILLER_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6716_ _5976_/A _8088_/Q _6724_/S vssd1 vssd1 vccd1 vccd1 _6717_/A sky130_fd_sc_hd__mux2_1
X_4977_ _4977_/A vssd1 vssd1 vccd1 vccd1 _8258_/D sky130_fd_sc_hd__clkbuf_1
X_3928_ _3950_/S vssd1 vssd1 vccd1 vccd1 _3941_/S sky130_fd_sc_hd__clkbuf_4
X_7696_ _8565_/Q _7698_/B vssd1 vssd1 vccd1 vccd1 _7696_/X sky130_fd_sc_hd__or2_1
XFILLER_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6647_ _6647_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _6663_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0__3428_ clkbuf_0__3428_/X vssd1 vssd1 vccd1 vccd1 _6980__408/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5529_ _8132_/Q _4438_/A _5531_/S vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__mux2_1
X_8317_ _8317_/CLK _8317_/D vssd1 vssd1 vccd1 vccd1 _8317_/Q sky130_fd_sc_hd__dfxtp_1
X_8248_ _8248_/CLK _8248_/D vssd1 vssd1 vccd1 vccd1 _8248_/Q sky130_fd_sc_hd__dfxtp_1
X_8179_ _8179_/CLK _8179_/D vssd1 vssd1 vccd1 vccd1 _8179_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3644_ clkbuf_0__3644_/X vssd1 vssd1 vccd1 vccd1 _7447__125/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3258_ _6632_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3258_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8646__211 vssd1 vssd1 vccd1 vccd1 _8646__211/HI caravel_irq[2] sky130_fd_sc_hd__conb_1
X_6201__176 _6204__179/A vssd1 vssd1 vccd1 vccd1 _7845_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5880_ _5880_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5896_/S sky130_fd_sc_hd__or2_2
X_4900_ _4869_/X _4890_/X _4893_/X _4899_/X _4683_/A vssd1 vssd1 vccd1 vccd1 _4900_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7230__101 _7231__102/A vssd1 vssd1 vccd1 vccd1 _8410_/CLK sky130_fd_sc_hd__inv_2
X_4831_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__buf_2
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4762_ _4758_/X _4759_/X _4761_/X vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7550_ _7550_/A _7550_/B vssd1 vssd1 vccd1 vccd1 _7573_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4693_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__buf_2
X_6501_ _6501_/A _6501_/B vssd1 vssd1 vccd1 vccd1 _6562_/A sky130_fd_sc_hd__nand2_1
X_6432_ _6499_/A vssd1 vssd1 vccd1 vccd1 _6501_/A sky130_fd_sc_hd__clkbuf_2
X_6811__356 _6813__358/A vssd1 vssd1 vccd1 vccd1 _8151_/CLK sky130_fd_sc_hd__inv_2
X_8102_ _8561_/CLK _8102_/D vssd1 vssd1 vccd1 vccd1 _8102_/Q sky130_fd_sc_hd__dfxtp_1
X_6363_ _6403_/A vssd1 vssd1 vccd1 vccd1 _6363_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5314_ _8352_/Q _5220_/X _5238_/X _8502_/Q _5165_/A vssd1 vssd1 vccd1 vccd1 _5314_/X
+ sky130_fd_sc_hd__o221a_1
X_6294_ _6294_/A vssd1 vssd1 vccd1 vccd1 _7898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _8386_/Q _8378_/Q _8370_/Q _8394_/Q _5138_/X _5131_/X vssd1 vssd1 vccd1 vccd1
+ _5245_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8033_ _8033_/CLK _8033_/D vssd1 vssd1 vccd1 vccd1 _8033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5176_ _3959_/X _5078_/X _5175_/X _5152_/X vssd1 vssd1 vccd1 vccd1 _8213_/D sky130_fd_sc_hd__o211a_1
X_4127_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4058_ _3971_/X _8519_/Q _4062_/S vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7817_ _7817_/A _7817_/B vssd1 vssd1 vccd1 vccd1 _7817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7679_ _7682_/A vssd1 vssd1 vccd1 vccd1 _7679_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7162__548 _7162__548/A vssd1 vssd1 vccd1 vccd1 _8357_/CLK sky130_fd_sc_hd__inv_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _8236_/D sky130_fd_sc_hd__clkbuf_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5932_ _6060_/A vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__clkbuf_2
X_6624__270 _6624__270/A vssd1 vssd1 vccd1 vccd1 _8030_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5878_/S vssd1 vssd1 vccd1 vccd1 _5872_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_34_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5794_ _7990_/Q _5598_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3661_ _7529_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3661_/X sky130_fd_sc_hd__clkbuf_16
X_4814_ _8252_/Q vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__clkbuf_1
X_8582_ _8582_/CLK _8582_/D vssd1 vssd1 vccd1 vccd1 _8582_/Q sky130_fd_sc_hd__dfxtp_2
X_7602_ _7664_/B _7580_/X _7599_/X _7601_/X vssd1 vssd1 vccd1 vccd1 _8542_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4745_ _4453_/X _4669_/X _4742_/X _4744_/X vssd1 vssd1 vccd1 vccd1 _8268_/D sky130_fd_sc_hd__o211a_1
X_7752__50 _7752__50/A vssd1 vssd1 vccd1 vccd1 _8601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4676_ _4684_/A vssd1 vssd1 vccd1 vccd1 _4680_/A sky130_fd_sc_hd__clkbuf_2
X_7395_ _8439_/Q _7384_/X _7360_/A _7394_/Y vssd1 vssd1 vccd1 vccd1 _7396_/B sky130_fd_sc_hd__o2bb2a_1
X_6415_ _6413_/Y _6385_/X _6414_/Y _6398_/X _6387_/X vssd1 vssd1 vccd1 vccd1 _6416_/C
+ sky130_fd_sc_hd__o221a_1
X_7063__468 _7063__468/A vssd1 vssd1 vccd1 vccd1 _8277_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8016_ _8016_/CLK _8016_/D vssd1 vssd1 vccd1 vccd1 _8016_/Q sky130_fd_sc_hd__dfxtp_1
Xinput107 wbs_we_i vssd1 vssd1 vccd1 vccd1 _6303_/C sky130_fd_sc_hd__buf_6
X_6277_ _8101_/Q _6222_/X _6236_/A _6272_/X _7890_/Q vssd1 vssd1 vccd1 vccd1 _7890_/D
+ sky130_fd_sc_hd__o32a_1
X_5228_ _5237_/A vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__clkbuf_2
X_5159_ _8600_/Q _8153_/Q _8126_/Q _8584_/Q _5122_/X _5123_/X vssd1 vssd1 vccd1 vccd1
+ _5159_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0_0__3412_ clkbuf_0__3412_/X vssd1 vssd1 vccd1 vccd1 _6927__379/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6687__305/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6567__224 _6568__225/A vssd1 vssd1 vccd1 vccd1 _7984_/CLK sky130_fd_sc_hd__inv_2
X_7474__146 _7477__149/A vssd1 vssd1 vccd1 vccd1 _8485_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7726__28 _7728__30/A vssd1 vssd1 vccd1 vccd1 _8579_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4530_ _4530_/A vssd1 vssd1 vccd1 vccd1 _8328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ _4460_/X _8349_/Q _4470_/S vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6200_ _6212_/A vssd1 vssd1 vccd1 vccd1 _6200_/X sky130_fd_sc_hd__buf_1
X_4392_ _4407_/S vssd1 vssd1 vccd1 vccd1 _4401_/S sky130_fd_sc_hd__buf_2
X_6131_ _7874_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__or2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6062_/A vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5013_ _5013_/A vssd1 vssd1 vccd1 vccd1 _8243_/D sky130_fd_sc_hd__clkbuf_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _6964_/A vssd1 vssd1 vccd1 vccd1 _6964_/X sky130_fd_sc_hd__buf_1
X_5915_ _5915_/A vssd1 vssd1 vccd1 vccd1 _7845_/D sky130_fd_sc_hd__clkbuf_1
X_6895_ _7814_/A _7590_/B _6893_/Y _6894_/X vssd1 vssd1 vccd1 vccd1 _6895_/X sky130_fd_sc_hd__o2bb2a_1
X_5846_ _4427_/X _7919_/Q _5854_/S vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__mux2_1
X_7347__113 _7347__113/A vssd1 vssd1 vccd1 vccd1 _8424_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777_ _5777_/A vssd1 vssd1 vccd1 vccd1 _7998_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3644_ _7442_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3644_/X sky130_fd_sc_hd__clkbuf_16
X_8565_ _8568_/CLK _8565_/D vssd1 vssd1 vccd1 vccd1 _8565_/Q sky130_fd_sc_hd__dfxtp_1
X_4728_ _4756_/S _4726_/X _4727_/X vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__a21o_1
X_8496_ _8496_/CLK _8496_/D vssd1 vssd1 vccd1 vccd1 _8496_/Q sky130_fd_sc_hd__dfxtp_1
X_4659_ _4659_/A vssd1 vssd1 vccd1 vccd1 _8273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7378_ _7386_/A _7378_/B vssd1 vssd1 vccd1 vccd1 _8432_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6329_ _6341_/A vssd1 vssd1 vccd1 vccd1 _6329_/X sky130_fd_sc_hd__buf_1
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3257_ clkbuf_0__3257_/X vssd1 vssd1 vccd1 vccd1 _6668_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8436_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _8592_/D sky130_fd_sc_hd__clkbuf_1
X_5700_ _5700_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5716_/S sky130_fd_sc_hd__or2_2
Xclkbuf_1_1_0__3461_ clkbuf_0__3461_/X vssd1 vssd1 vccd1 vccd1 _7147_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6680_ _7541_/A vssd1 vssd1 vccd1 vccd1 _6680_/X sky130_fd_sc_hd__buf_1
X_3892_ _8199_/Q _8204_/Q vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__and2b_1
X_5631_ _8068_/Q _5630_/X _5634_/S vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__mux2_1
X_5562_ _5562_/A vssd1 vssd1 vccd1 vccd1 _8118_/D sky130_fd_sc_hd__clkbuf_1
X_8350_ _8350_/CLK _8350_/D vssd1 vssd1 vccd1 vccd1 _8350_/Q sky130_fd_sc_hd__dfxtp_1
X_4513_ _8194_/Q vssd1 vssd1 vccd1 vccd1 _4513_/X sky130_fd_sc_hd__clkbuf_4
X_8281_ _8281_/CLK _8281_/D vssd1 vssd1 vccd1 vccd1 _8281_/Q sky130_fd_sc_hd__dfxtp_1
X_7301_ _8437_/Q _7308_/A _7308_/B _7308_/C vssd1 vssd1 vccd1 vccd1 _7303_/A sky130_fd_sc_hd__nand4_1
X_5493_ _8151_/Q _4492_/X _5495_/S vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__mux2_1
X_4444_ _4444_/A vssd1 vssd1 vccd1 vccd1 _4444_/X sky130_fd_sc_hd__clkbuf_2
X_4375_ _8382_/Q _4215_/X _4383_/S vssd1 vssd1 vccd1 vccd1 _4376_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6114_ _7945_/Q input34/X _6125_/S vssd1 vssd1 vccd1 vccd1 _6114_/X sky130_fd_sc_hd__mux2_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _8088_/Q _6047_/B vssd1 vssd1 vccd1 vccd1 _6046_/A sky130_fd_sc_hd__and2_1
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _7996_/CLK _7996_/D vssd1 vssd1 vccd1 vccd1 _7996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6947_ _8564_/Q _6947_/B vssd1 vssd1 vccd1 vccd1 _6948_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3659_ clkbuf_0__3659_/X vssd1 vssd1 vccd1 vccd1 _7521__9/A sky130_fd_sc_hd__clkbuf_4
X_6878_ _6872_/X _6873_/Y _6875_/Y _6877_/X vssd1 vssd1 vccd1 vccd1 _7582_/A sky130_fd_sc_hd__o211a_1
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5829_ _5829_/A vssd1 vssd1 vccd1 vccd1 _7927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8617_ _8617_/CLK _8617_/D vssd1 vssd1 vccd1 vccd1 _8617_/Q sky130_fd_sc_hd__dfxtp_1
X_8548_ _8553_/CLK _8548_/D vssd1 vssd1 vccd1 vccd1 _8548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6637__280 _6637__280/A vssd1 vssd1 vccd1 vccd1 _8040_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8479_ _8479_/CLK _8479_/D vssd1 vssd1 vccd1 vccd1 _8479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3309_ clkbuf_0__3309_/X vssd1 vssd1 vccd1 vccd1 _6785_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7076__478 _7078__480/A vssd1 vssd1 vccd1 vccd1 _8287_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput208 _6116_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_57_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4508_/B _5663_/B _5663_/A vssd1 vssd1 vccd1 vccd1 _5645_/A sky130_fd_sc_hd__or3b_4
XFILLER_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4091_ _8506_/Q _3934_/X _4095_/S vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7850_ _7850_/CLK _7850_/D vssd1 vssd1 vccd1 vccd1 _7850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _6801_/A vssd1 vssd1 vccd1 vccd1 _8144_/D sky130_fd_sc_hd__clkbuf_1
X_7538__23 _7540__25/A vssd1 vssd1 vccd1 vccd1 _8537_/CLK sky130_fd_sc_hd__inv_2
X_7781_ _5982_/A _7778_/X _7777_/A vssd1 vssd1 vccd1 vccd1 _7781_/X sky130_fd_sc_hd__a21bo_1
X_4993_ _4716_/A _4988_/X _4992_/Y _4903_/X vssd1 vssd1 vccd1 vccd1 _8253_/D sky130_fd_sc_hd__o211a_1
X_7487__156 _7488__157/A vssd1 vssd1 vccd1 vccd1 _8495_/CLK sky130_fd_sc_hd__inv_2
X_3944_ _8596_/Q _3943_/X _3950_/S vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__mux2_1
X_6732_ _6732_/A _6732_/B vssd1 vssd1 vccd1 vccd1 _6748_/S sky130_fd_sc_hd__and2_4
X_3875_ _8205_/Q vssd1 vssd1 vccd1 vccd1 _4336_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6663_ _8268_/Q _6663_/B vssd1 vssd1 vccd1 vccd1 _6664_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3444_ clkbuf_0__3444_/X vssd1 vssd1 vccd1 vccd1 _7049__459/A sky130_fd_sc_hd__clkbuf_4
X_8402_ _8402_/CLK _8402_/D vssd1 vssd1 vccd1 vccd1 _8402_/Q sky130_fd_sc_hd__dfxtp_1
X_5614_ _5613_/X _8073_/Q _5617_/S vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3412_ _6923_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3412_/X sky130_fd_sc_hd__clkbuf_16
X_6594_ _6594_/A vssd1 vssd1 vccd1 vccd1 _6594_/X sky130_fd_sc_hd__buf_1
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8333_ _8333_/CLK _8333_/D vssd1 vssd1 vccd1 vccd1 _8333_/Q sky130_fd_sc_hd__dfxtp_1
X_5545_ _8125_/Q _4435_/A _5549_/S vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5476_ _5476_/A vssd1 vssd1 vccd1 vccd1 _8159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7171__54 _7172__55/A vssd1 vssd1 vccd1 vccd1 _8363_/CLK sky130_fd_sc_hd__inv_2
X_8663__228 vssd1 vssd1 vccd1 vccd1 _8663__228/HI manufacturerID[0] sky130_fd_sc_hd__conb_1
X_8264_ _8264_/CLK _8264_/D vssd1 vssd1 vccd1 vccd1 _8264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4427_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3274_ _6682_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3274_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3660_ clkbuf_0__3660_/X vssd1 vssd1 vccd1 vccd1 _7528__15/A sky130_fd_sc_hd__clkbuf_4
X_8195_ _8568_/CLK _8195_/D vssd1 vssd1 vccd1 vccd1 _8195_/Q sky130_fd_sc_hd__dfxtp_4
X_4358_ _4358_/A vssd1 vssd1 vccd1 vccd1 _8390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _8421_/Q _4200_/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4290_/A sky130_fd_sc_hd__mux2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6028_ _6028_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6029_/A sky130_fd_sc_hd__and2_1
XFILLER_104_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7226__99 _7226__99/A vssd1 vssd1 vccd1 vccd1 _8408_/CLK sky130_fd_sc_hd__inv_2
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7979_ _8270_/CLK _7979_/D vssd1 vssd1 vccd1 vccd1 _7979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6982__410 _6982__410/A vssd1 vssd1 vccd1 vccd1 _8214_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_80 _7842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_91 _6088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6321__195 _6321__195/A vssd1 vssd1 vccd1 vccd1 _7907_/CLK sky130_fd_sc_hd__inv_2
X_5330_ _8408_/Q _8129_/Q _5330_/S vssd1 vssd1 vccd1 vccd1 _5330_/X sky130_fd_sc_hd__mux2_1
X_7126__519 _7127__520/A vssd1 vssd1 vccd1 vccd1 _8328_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5261_ _8410_/Q _8131_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__mux2_1
X_7000_ _7000_/A vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__buf_1
X_4212_ _8188_/Q vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__clkbuf_4
X_5192_ _5247_/A _5187_/X _5189_/X _5191_/X _5217_/A vssd1 vssd1 vccd1 vccd1 _5192_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ _4143_/A vssd1 vssd1 vccd1 vccd1 _8491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4074_ _8513_/Q _3937_/X _4076_/S vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7902_ _8441_/CLK _7902_/D vssd1 vssd1 vccd1 vccd1 _7902_/Q sky130_fd_sc_hd__dfxtp_1
X_7833_ _8629_/Q _7840_/C _7832_/X _7763_/A vssd1 vssd1 vccd1 vccd1 _8629_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7764_ _7764_/A vssd1 vssd1 vccd1 vccd1 _8608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6715_ _6730_/S vssd1 vssd1 vccd1 vccd1 _6724_/S sky130_fd_sc_hd__buf_2
X_4976_ _7053_/C _4976_/B _4976_/C vssd1 vssd1 vccd1 vccd1 _4977_/A sky130_fd_sc_hd__and3_1
X_3927_ _5539_/A _5826_/A vssd1 vssd1 vccd1 vccd1 _3950_/S sky130_fd_sc_hd__nor2_2
X_7695_ _8565_/Q _7687_/X _7694_/X _7684_/X vssd1 vssd1 vccd1 vccd1 _8564_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1_0__3427_ clkbuf_0__3427_/X vssd1 vssd1 vccd1 vccd1 _6975__404/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5528_ _5528_/A vssd1 vssd1 vccd1 vccd1 _8133_/D sky130_fd_sc_hd__clkbuf_1
X_8316_ _8316_/CLK _8316_/D vssd1 vssd1 vccd1 vccd1 _8316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5459_ _5416_/X _8167_/Q _5459_/S vssd1 vssd1 vccd1 vccd1 _5460_/A sky130_fd_sc_hd__mux2_1
X_8247_ _8247_/CLK _8247_/D vssd1 vssd1 vccd1 vccd1 _8247_/Q sky130_fd_sc_hd__dfxtp_1
X_8178_ _8178_/CLK _8178_/D vssd1 vssd1 vccd1 vccd1 _8178_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3257_ _6631_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3257_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3643_ clkbuf_0__3643_/X vssd1 vssd1 vccd1 vccd1 _7438__117/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7532__18 _7532__18/A vssd1 vssd1 vccd1 vccd1 _8532_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7438__117 _7438__117/A vssd1 vssd1 vccd1 vccd1 _8456_/CLK sky130_fd_sc_hd__inv_2
X_6763__323 _6763__323/A vssd1 vssd1 vccd1 vccd1 _8115_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4830_ _8282_/Q _4829_/X _4822_/X _8244_/Q vssd1 vssd1 vccd1 vccd1 _4830_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4713_/A _4760_/X _4841_/A vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__a21o_1
X_4692_ _8251_/Q vssd1 vssd1 vccd1 vccd1 _4729_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7480_ _7504_/A vssd1 vssd1 vccd1 vccd1 _7480_/X sky130_fd_sc_hd__buf_1
X_6500_ _6500_/A _7575_/A _7757_/B _6983_/B vssd1 vssd1 vccd1 vccd1 _6563_/B sky130_fd_sc_hd__or4b_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6431_ _7941_/Q _6410_/X _6430_/Y _6423_/X vssd1 vssd1 vccd1 vccd1 _7941_/D sky130_fd_sc_hd__a211o_1
X_7341__108 _7342__109/A vssd1 vssd1 vccd1 vccd1 _8419_/CLK sky130_fd_sc_hd__inv_2
X_6362_ _8144_/Q _6448_/C vssd1 vssd1 vccd1 vccd1 _6403_/A sky130_fd_sc_hd__and2_2
X_5313_ _8400_/Q _8137_/Q _5313_/S vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__mux2_1
X_8101_ _8569_/CLK _8101_/D vssd1 vssd1 vccd1 vccd1 _8101_/Q sky130_fd_sc_hd__dfxtp_1
X_6293_ _7719_/A _7898_/Q _6297_/S vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5244_ _8504_/Q _8402_/Q _8139_/Q _8354_/Q _5123_/A _5140_/X vssd1 vssd1 vccd1 vccd1
+ _5244_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8032_ _8032_/CLK _8032_/D vssd1 vssd1 vccd1 vccd1 _8032_/Q sky130_fd_sc_hd__dfxtp_1
X_5175_ _8213_/Q _5080_/X _5385_/A _5174_/X _5148_/X vssd1 vssd1 vccd1 vccd1 _5175_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4126_ _8572_/Q vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__buf_2
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4057_ _4057_/A vssd1 vssd1 vccd1 vccd1 _8520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7816_ _7814_/Y _7815_/Y _7800_/X vssd1 vssd1 vccd1 vccd1 _8624_/D sky130_fd_sc_hd__a21oi_1
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7747_ _7747_/A vssd1 vssd1 vccd1 vccd1 _7747_/X sky130_fd_sc_hd__buf_1
X_4959_ _4735_/X _4949_/X _4952_/X _4958_/X _4683_/A vssd1 vssd1 vccd1 vccd1 _4959_/X
+ sky130_fd_sc_hd__o311a_1
X_7678_ _8560_/Q _7671_/Y _7677_/X _7601_/X vssd1 vssd1 vccd1 vccd1 _8560_/D sky130_fd_sc_hd__o211a_1
X_8669__234 vssd1 vssd1 vccd1 vccd1 _8669__234/HI manufacturerID[6] sky130_fd_sc_hd__conb_1
XFILLER_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3309_ _6766_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3309_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _5931_/A vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5862_ _5862_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5878_/S sky130_fd_sc_hd__nor2_2
XFILLER_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5793_ _5793_/A vssd1 vssd1 vccd1 vccd1 _7991_/D sky130_fd_sc_hd__clkbuf_1
X_4813_ _4812_/X _8183_/Q _8075_/Q _4665_/X vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_0__3660_ _7523_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3660_/X sky130_fd_sc_hd__clkbuf_16
X_8581_ _8581_/CLK _8581_/D vssd1 vssd1 vccd1 vccd1 _8581_/Q sky130_fd_sc_hd__dfxtp_1
X_7601_ _7628_/B vssd1 vssd1 vccd1 vccd1 _7601_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _6947_/B vssd1 vssd1 vccd1 vccd1 _4744_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4675_ _8252_/Q vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__inv_2
X_7394_ _7394_/A _7394_/B vssd1 vssd1 vccd1 vccd1 _7394_/Y sky130_fd_sc_hd__nand2_1
X_6414_ _8051_/Q _6395_/X _6382_/X vssd1 vssd1 vccd1 vccd1 _6414_/Y sky130_fd_sc_hd__a21oi_1
X_6276_ _8100_/Q _6222_/X _6270_/X _6272_/X _7889_/Q vssd1 vssd1 vccd1 vccd1 _7889_/D
+ sky130_fd_sc_hd__o32a_1
X_8015_ _8015_/CLK _8015_/D vssd1 vssd1 vccd1 vccd1 _8015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5227_ _8322_/Q _8338_/Q _5355_/S vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5158_ _7926_/Q _8134_/Q _8413_/Q _8161_/Q _5313_/S _5110_/X vssd1 vssd1 vccd1 vccd1
+ _5158_/X sky130_fd_sc_hd__mux4_2
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _4109_/A vssd1 vssd1 vccd1 vccd1 _8500_/D sky130_fd_sc_hd__clkbuf_1
X_7139__529 _7139__529/A vssd1 vssd1 vccd1 vccd1 _8338_/CLK sky130_fd_sc_hd__inv_2
X_5089_ _8196_/Q vssd1 vssd1 vccd1 vccd1 _5222_/B sky130_fd_sc_hd__buf_2
XFILLER_112_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6694_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8643__259 vssd1 vssd1 vccd1 vccd1 partID[15] _8643__259/LO sky130_fd_sc_hd__conb_1
XFILLER_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6574__229 _6575__230/A vssd1 vssd1 vccd1 vccd1 _7989_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4460_ _8194_/Q vssd1 vssd1 vccd1 vccd1 _4460_/X sky130_fd_sc_hd__clkbuf_4
X_4391_ _5844_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4407_/S sky130_fd_sc_hd__or2_2
X_6130_ _6149_/A vssd1 vssd1 vccd1 vccd1 _6145_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6061_ _8095_/Q _6069_/B vssd1 vssd1 vccd1 vccd1 _6062_/A sky130_fd_sc_hd__and2_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6214__187 _6217__190/A vssd1 vssd1 vccd1 vccd1 _7856_/CLK sky130_fd_sc_hd__inv_2
X_5012_ _8243_/Q _4525_/X _5016_/S vssd1 vssd1 vccd1 vccd1 _5013_/A sky130_fd_sc_hd__mux2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6776__333 _6776__333/A vssd1 vssd1 vccd1 vccd1 _8125_/CLK sky130_fd_sc_hd__inv_2
X_5914_ _4212_/X _7845_/Q _5914_/S vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__mux2_1
X_6894_ _8625_/Q _7551_/A _7551_/B vssd1 vssd1 vccd1 vccd1 _6894_/X sky130_fd_sc_hd__and3_1
X_5845_ _5860_/S vssd1 vssd1 vccd1 vccd1 _5854_/S sky130_fd_sc_hd__clkbuf_2
X_8633_ _8633_/CLK _8633_/D vssd1 vssd1 vccd1 vccd1 _8633_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5776_ _7998_/Q _5598_/A _5782_/S vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3643_ _7436_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3643_/X sky130_fd_sc_hd__clkbuf_16
X_8564_ _8568_/CLK _8564_/D vssd1 vssd1 vccd1 vccd1 _8564_/Q sky130_fd_sc_hd__dfxtp_1
X_8495_ _8495_/CLK _8495_/D vssd1 vssd1 vccd1 vccd1 _8495_/Q sky130_fd_sc_hd__dfxtp_1
X_4727_ _4841_/A vssd1 vssd1 vccd1 vccd1 _4727_/X sky130_fd_sc_hd__buf_2
XFILLER_108_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4658_ _8273_/Q _4498_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput90 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__buf_4
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4589_ _4450_/X _8303_/Q _4589_/S vssd1 vssd1 vccd1 vccd1 _4590_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7377_ _8432_/Q _7368_/X _7376_/X _7263_/B vssd1 vssd1 vccd1 vccd1 _7378_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6328_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6328_/X sky130_fd_sc_hd__buf_1
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6257_/X _8089_/Q _6253_/X _6255_/X _7878_/Q vssd1 vssd1 vccd1 vccd1 _7878_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6824__367 _6824__367/A vssd1 vssd1 vccd1 vccd1 _8162_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3256_ clkbuf_0__3256_/X vssd1 vssd1 vccd1 vccd1 _6630__275/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7731__32 _7732__33/A vssd1 vssd1 vccd1 vccd1 _8583_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ _3959_/X _8592_/Q _3969_/S vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3460_ clkbuf_0__3460_/X vssd1 vssd1 vccd1 vccd1 _7132__524/A sky130_fd_sc_hd__clkbuf_4
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _8204_/Q _5112_/A vssd1 vssd1 vccd1 vccd1 _3893_/A sky130_fd_sc_hd__and2b_1
X_5630_ _8192_/Q vssd1 vssd1 vccd1 vccd1 _5630_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5561_ _5404_/X _8118_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5562_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4512_ _4512_/A vssd1 vssd1 vccd1 vccd1 _8334_/D sky130_fd_sc_hd__clkbuf_1
X_5492_ _5492_/A vssd1 vssd1 vccd1 vccd1 _8152_/D sky130_fd_sc_hd__clkbuf_1
X_8280_ _8280_/CLK _8280_/D vssd1 vssd1 vccd1 vccd1 _8280_/Q sky130_fd_sc_hd__dfxtp_1
X_7300_ _8625_/Q _7379_/A _7379_/B vssd1 vssd1 vccd1 vccd1 _7300_/X sky130_fd_sc_hd__and3_1
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4443_ _4443_/A vssd1 vssd1 vccd1 vccd1 _8354_/D sky130_fd_sc_hd__clkbuf_1
X_4374_ _4389_/S vssd1 vssd1 vccd1 vccd1 _4383_/S sky130_fd_sc_hd__buf_2
X_6113_ _6098_/X _6110_/X _6112_/X _6101_/X vssd1 vssd1 vccd1 vccd1 _6113_/X sky130_fd_sc_hd__o211a_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6044_/A vssd1 vssd1 vccd1 vccd1 _6044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7995_ _7995_/CLK _7995_/D vssd1 vssd1 vccd1 vccd1 _7995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6946_ _6946_/A vssd1 vssd1 vccd1 vccd1 _8189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3658_ clkbuf_0__3658_/X vssd1 vssd1 vccd1 vccd1 _7513__2/A sky130_fd_sc_hd__clkbuf_4
X_6877_ _8633_/Q _7603_/A vssd1 vssd1 vccd1 vccd1 _6877_/X sky130_fd_sc_hd__xor2_1
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5828_ _7927_/Q _4427_/A _5836_/S vssd1 vssd1 vccd1 vccd1 _5829_/A sky130_fd_sc_hd__mux2_1
X_8616_ _8617_/CLK _8616_/D vssd1 vssd1 vccd1 vccd1 _8616_/Q sky130_fd_sc_hd__dfxtp_2
X_5759_ _5759_/A vssd1 vssd1 vccd1 vccd1 _8006_/D sky130_fd_sc_hd__clkbuf_1
X_8547_ _8553_/CLK _8547_/D vssd1 vssd1 vccd1 vccd1 _8547_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8478_ _8478_/CLK _8478_/D vssd1 vssd1 vccd1 vccd1 _8478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7429_ _8213_/Q _7411_/A _7413_/A _7428_/X _7420_/X vssd1 vssd1 vccd1 vccd1 _8450_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3308_ clkbuf_0__3308_/X vssd1 vssd1 vccd1 vccd1 _6763__323/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7013__430 _7013__430/A vssd1 vssd1 vccd1 vccd1 _8236_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _4090_/A vssd1 vssd1 vccd1 vccd1 _8507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _6281_/A _8144_/Q _6804_/S vssd1 vssd1 vccd1 vccd1 _6801_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7780_ _8613_/Q _7777_/X _7779_/X _6503_/X vssd1 vssd1 vccd1 vccd1 _8613_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4992_ _4996_/A _4992_/B vssd1 vssd1 vccd1 vccd1 _4992_/Y sky130_fd_sc_hd__nand2_1
X_3943_ _8572_/Q vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__buf_2
X_6731_ _6731_/A vssd1 vssd1 vccd1 vccd1 _8095_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3443_ clkbuf_0__3443_/X vssd1 vssd1 vccd1 vccd1 _7041__452/A sky130_fd_sc_hd__clkbuf_4
X_6662_ _6662_/A vssd1 vssd1 vccd1 vccd1 _8054_/D sky130_fd_sc_hd__clkbuf_1
X_3874_ _4027_/B vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__buf_2
X_8401_ _8401_/CLK _8401_/D vssd1 vssd1 vccd1 vccd1 _8401_/Q sky130_fd_sc_hd__dfxtp_1
X_5613_ _5613_/A vssd1 vssd1 vccd1 vccd1 _5613_/X sky130_fd_sc_hd__clkbuf_2
X_8332_ _8332_/CLK _8332_/D vssd1 vssd1 vccd1 vccd1 _8332_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3411_ _6922_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3411_/X sky130_fd_sc_hd__clkbuf_16
X_5544_ _5544_/A vssd1 vssd1 vccd1 vccd1 _8126_/D sky130_fd_sc_hd__clkbuf_1
X_5475_ _4438_/X _8159_/Q _5477_/S vssd1 vssd1 vccd1 vccd1 _5476_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8263_ _8263_/CLK _8263_/D vssd1 vssd1 vccd1 vccd1 _8263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3273_ _6681_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3273_/X sky130_fd_sc_hd__clkbuf_16
X_6333__204 _6334__205/A vssd1 vssd1 vccd1 vccd1 _7916_/CLK sky130_fd_sc_hd__inv_2
X_4426_ _4426_/A vssd1 vssd1 vccd1 vccd1 _8359_/D sky130_fd_sc_hd__clkbuf_1
X_8194_ _8568_/CLK _8194_/D vssd1 vssd1 vccd1 vccd1 _8194_/Q sky130_fd_sc_hd__dfxtp_4
X_4357_ _4104_/X _8390_/Q _4365_/S vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__mux2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4288_/A vssd1 vssd1 vccd1 vccd1 _8422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6036_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7978_ _8270_/CLK _7978_/D vssd1 vssd1 vccd1 vccd1 _7978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6935_/A vssd1 vssd1 vccd1 vccd1 _6929_/X sky130_fd_sc_hd__buf_1
XFILLER_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7082__483 _7083__484/A vssd1 vssd1 vccd1 vccd1 _8292_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_70 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_92 _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_81 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5260_ _8597_/Q _5257_/X _5120_/A _5259_/X vssd1 vssd1 vccd1 vccd1 _5264_/B sky130_fd_sc_hd__o211a_1
XFILLER_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4211_ _4211_/A vssd1 vssd1 vccd1 vccd1 _8478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191_ _5135_/X _5190_/X _5171_/X vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__a21o_1
X_4142_ _8491_/Q _3931_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4143_/A sky130_fd_sc_hd__mux2_1
X_7493__161 _7497__165/A vssd1 vssd1 vccd1 vccd1 _8500_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4073_ _4073_/A vssd1 vssd1 vccd1 vccd1 _8514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7901_ _8441_/CLK _7901_/D vssd1 vssd1 vccd1 vccd1 _7901_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8556_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7832_ _7716_/A _7723_/B _7826_/A vssd1 vssd1 vccd1 vccd1 _7832_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7763_ _7763_/A _8602_/Q vssd1 vssd1 vccd1 vccd1 _7764_/A sky130_fd_sc_hd__and2_1
X_4975_ _8269_/Q _4969_/B _7753_/B _5055_/B vssd1 vssd1 vccd1 vccd1 _4976_/C sky130_fd_sc_hd__a31o_1
X_3926_ _4355_/A vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__clkbuf_4
X_6714_ _6714_/A _6732_/B vssd1 vssd1 vccd1 vccd1 _6730_/S sky130_fd_sc_hd__nand2_2
Xclkbuf_1_1_0__3426_ clkbuf_0__3426_/X vssd1 vssd1 vccd1 vccd1 _7000_/A sky130_fd_sc_hd__clkbuf_4
X_7694_ _8564_/Q _7698_/B vssd1 vssd1 vccd1 vccd1 _7694_/X sky130_fd_sc_hd__or2_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6576_ _6576_/A vssd1 vssd1 vccd1 vccd1 _6576_/X sky130_fd_sc_hd__buf_1
X_5527_ _8133_/Q _4435_/A _5531_/S vssd1 vssd1 vccd1 vccd1 _5528_/A sky130_fd_sc_hd__mux2_1
X_8315_ _8315_/CLK _8315_/D vssd1 vssd1 vccd1 vccd1 _8315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8246_ _8246_/CLK _8246_/D vssd1 vssd1 vccd1 vccd1 _8246_/Q sky130_fd_sc_hd__dfxtp_1
X_5458_ _5458_/A vssd1 vssd1 vccd1 vccd1 _8168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8177_ _8177_/CLK _8177_/D vssd1 vssd1 vccd1 vccd1 _8177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3256_ _6625_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3256_/X sky130_fd_sc_hd__clkbuf_16
X_4409_ _4534_/A _5467_/A vssd1 vssd1 vccd1 vccd1 _4425_/S sky130_fd_sc_hd__or2_4
X_5389_ _5393_/A _5389_/B vssd1 vssd1 vccd1 vccd1 _5389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7128_ _7128_/A vssd1 vssd1 vccd1 vccd1 _7128_/X sky130_fd_sc_hd__buf_1
XFILLER_115_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7132__524 _7132__524/A vssd1 vssd1 vccd1 vccd1 _8333_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _7910_/Q _8030_/Q _8046_/Q _8014_/Q _4955_/S _4702_/A vssd1 vssd1 vccd1 vccd1
+ _4760_/X sky130_fd_sc_hd__mux4_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4691_ _4691_/A vssd1 vssd1 vccd1 vccd1 _4691_/X sky130_fd_sc_hd__buf_4
X_6770__328 _6772__330/A vssd1 vssd1 vccd1 vccd1 _8120_/CLK sky130_fd_sc_hd__inv_2
X_7089__489 _7089__489/A vssd1 vssd1 vccd1 vccd1 _8298_/CLK sky130_fd_sc_hd__inv_2
X_6430_ _6430_/A _6430_/B _6430_/C vssd1 vssd1 vccd1 vccd1 _6430_/Y sky130_fd_sc_hd__nor3_1
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6361_ _6361_/A vssd1 vssd1 vccd1 vccd1 _6448_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_115_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5312_ _5393_/B _5310_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _5312_/Y sky130_fd_sc_hd__o21ai_1
X_8100_ _8569_/CLK _8100_/D vssd1 vssd1 vccd1 vccd1 _8100_/Q sky130_fd_sc_hd__dfxtp_1
X_6292_ _6292_/A vssd1 vssd1 vccd1 vccd1 _7897_/D sky130_fd_sc_hd__clkbuf_1
X_8031_ _8031_/CLK _8031_/D vssd1 vssd1 vccd1 vccd1 _8031_/Q sky130_fd_sc_hd__dfxtp_1
X_5243_ _5391_/B _5231_/X _5241_/X _5389_/B vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__a211o_1
X_5174_ _5087_/X _5157_/X _5161_/X _5173_/X vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__a31o_2
X_4125_ _4125_/A vssd1 vssd1 vccd1 vccd1 _8496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4056_ _3968_/X _8520_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7815_ _7815_/A _7818_/B vssd1 vssd1 vccd1 vccd1 _7815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4958_ _4953_/X _4954_/X _4957_/X _4727_/X vssd1 vssd1 vccd1 vccd1 _4958_/X sky130_fd_sc_hd__a211o_1
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4889_ _8479_/Q _4680_/A _4833_/X _8455_/Q _4687_/A vssd1 vssd1 vccd1 vccd1 _4889_/X
+ sky130_fd_sc_hd__o221a_1
X_7677_ _7677_/A _7682_/B _7677_/C vssd1 vssd1 vccd1 vccd1 _7677_/X sky130_fd_sc_hd__or3_1
X_3909_ _7982_/Q _7981_/Q vssd1 vssd1 vccd1 vccd1 _6499_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6559_ _6505_/A _7778_/A _6195_/C _6448_/C vssd1 vssd1 vccd1 vccd1 _6563_/C sky130_fd_sc_hd__a31o_1
XFILLER_106_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8229_ _8229_/CLK _8229_/D vssd1 vssd1 vccd1 vccd1 _8229_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3308_ _6760_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3308_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7738__38 _7738__38/A vssd1 vssd1 vccd1 vccd1 _8589_/CLK sky130_fd_sc_hd__inv_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7444__122 _7447__125/A vssd1 vssd1 vccd1 vccd1 _8461_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6921__375 _6921__375/A vssd1 vssd1 vccd1 vccd1 _8171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5930_ _6696_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__and2_1
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5861_ _5861_/A vssd1 vssd1 vccd1 vccd1 _7912_/D sky130_fd_sc_hd__clkbuf_1
X_7600_ _7600_/A vssd1 vssd1 vccd1 vccd1 _7628_/B sky130_fd_sc_hd__clkbuf_2
X_5792_ _7991_/Q _5593_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5793_/A sky130_fd_sc_hd__mux2_1
X_4812_ _4812_/A vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__buf_2
X_8580_ _8580_/CLK _8580_/D vssd1 vssd1 vccd1 vccd1 _8580_/Q sky130_fd_sc_hd__dfxtp_1
X_4743_ _4981_/A vssd1 vssd1 vccd1 vccd1 _6947_/B sky130_fd_sc_hd__buf_2
XFILLER_119_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6413_ _8610_/Q vssd1 vssd1 vccd1 vccd1 _6413_/Y sky130_fd_sc_hd__inv_2
X_4674_ _4989_/A vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7393_ _7398_/A _7393_/B vssd1 vssd1 vccd1 vccd1 _8438_/D sky130_fd_sc_hd__nor2_1
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670__292 _6673__295/A vssd1 vssd1 vccd1 vccd1 _8060_/CLK sky130_fd_sc_hd__inv_2
X_6275_ _8099_/Q _6269_/X _6270_/X _6272_/X _7888_/Q vssd1 vssd1 vccd1 vccd1 _7888_/D
+ sky130_fd_sc_hd__o32a_1
X_8014_ _8014_/CLK _8014_/D vssd1 vssd1 vccd1 vccd1 _8014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5226_ _5283_/S vssd1 vssd1 vccd1 vccd1 _5355_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_102_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3410_ clkbuf_0__3410_/X vssd1 vssd1 vccd1 vccd1 _6921__375/A sky130_fd_sc_hd__clkbuf_4
X_5157_ _5095_/X _5154_/X _5156_/X vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _4104_/X _8500_/Q _4124_/S vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5088_ _8197_/Q vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6970_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4039_ _4039_/A vssd1 vssd1 vccd1 vccd1 _8528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ _7735_/A vssd1 vssd1 vccd1 vccd1 _7729_/X sky130_fd_sc_hd__buf_1
XFILLER_40_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7508__174 _7509__175/A vssd1 vssd1 vccd1 vccd1 _8513_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6608__256 _6611__259/A vssd1 vssd1 vccd1 vccd1 _8016_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6689__306 _6690__307/A vssd1 vssd1 vccd1 vccd1 _8074_/CLK sky130_fd_sc_hd__inv_2
X_4390_ _4390_/A vssd1 vssd1 vccd1 vccd1 _8375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6060_/A vssd1 vssd1 vccd1 vccd1 _6069_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5011_ _5011_/A vssd1 vssd1 vccd1 vccd1 _8244_/D sky130_fd_sc_hd__clkbuf_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0__3812_ clkbuf_0__3812_/X vssd1 vssd1 vccd1 vccd1 _7752__50/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6893_ _7551_/A _7551_/B _7817_/A vssd1 vssd1 vccd1 vccd1 _6893_/Y sky130_fd_sc_hd__a21oi_1
X_5913_ _5913_/A vssd1 vssd1 vccd1 vccd1 _7846_/D sky130_fd_sc_hd__clkbuf_1
X_5844_ _5844_/A _5844_/B vssd1 vssd1 vccd1 vccd1 _5860_/S sky130_fd_sc_hd__or2_4
X_8632_ _8633_/CLK _8632_/D vssd1 vssd1 vccd1 vccd1 _8632_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8563_ _8568_/CLK _8563_/D vssd1 vssd1 vccd1 vccd1 _8563_/Q sky130_fd_sc_hd__dfxtp_1
X_5775_ _5775_/A vssd1 vssd1 vccd1 vccd1 _7999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4726_ _7852_/Q _7860_/Q _7935_/Q _8039_/Q _4721_/X _4725_/X vssd1 vssd1 vccd1 vccd1
+ _4726_/X sky130_fd_sc_hd__mux4_1
X_8494_ _8494_/CLK _8494_/D vssd1 vssd1 vccd1 vccd1 _8494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4657_ _4657_/A vssd1 vssd1 vccd1 vccd1 _8274_/D sky130_fd_sc_hd__clkbuf_1
X_7145__534 _7146__535/A vssd1 vssd1 vccd1 vccd1 _8343_/CLK sky130_fd_sc_hd__inv_2
Xinput80 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _5982_/A sky130_fd_sc_hd__buf_4
Xinput91 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _6004_/A sky130_fd_sc_hd__buf_4
X_7376_ _7376_/A vssd1 vssd1 vccd1 vccd1 _7376_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4588_ _4588_/A vssd1 vssd1 vccd1 vccd1 _8304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6258_ _6257_/X _8088_/Q _6253_/X _6255_/X _7877_/Q vssd1 vssd1 vccd1 vccd1 _7877_/D
+ sky130_fd_sc_hd__o32a_1
X_5209_ _5209_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__and2_1
XFILLER_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6189_ _7892_/Q _6088_/B _6176_/A _6188_/X _6101_/A vssd1 vssd1 vccd1 vccd1 _6189_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3255_ clkbuf_0__3255_/X vssd1 vssd1 vccd1 vccd1 _6621__267/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6677__298 _6678__299/A vssd1 vssd1 vccd1 vccd1 _8066_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6580__234 _6581__235/A vssd1 vssd1 vccd1 vccd1 _7994_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _5075_/A _5370_/A vssd1 vssd1 vccd1 vccd1 _3899_/B sky130_fd_sc_hd__and2b_1
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5560_/A vssd1 vssd1 vccd1 vccd1 _8119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4511_ _8334_/Q _4507_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4512_/A sky130_fd_sc_hd__mux2_1
X_7183__64 _7183__64/A vssd1 vssd1 vccd1 vccd1 _8373_/CLK sky130_fd_sc_hd__inv_2
X_5491_ _8152_/Q _4489_/X _5495_/S vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4442_ _4441_/X _8354_/Q _4442_/S vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4373_ _5521_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4389_/S sky130_fd_sc_hd__nor2_2
X_6112_ _7869_/Q _6126_/B vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__or2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _8087_/Q _6047_/B vssd1 vssd1 vccd1 vccd1 _6044_/A sky130_fd_sc_hd__and2_1
XFILLER_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7457__132 _7458__133/A vssd1 vssd1 vccd1 vccd1 _8471_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7994_ _7994_/CLK _7994_/D vssd1 vssd1 vccd1 vccd1 _7994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6945_ _8563_/Q _6947_/B vssd1 vssd1 vccd1 vccd1 _6946_/A sky130_fd_sc_hd__and2_1
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3657_ clkbuf_0__3657_/X vssd1 vssd1 vccd1 vccd1 _7535_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_6876_ _6876_/A vssd1 vssd1 vccd1 vccd1 _7603_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5827_ _5842_/S vssd1 vssd1 vccd1 vccd1 _5836_/S sky130_fd_sc_hd__buf_2
XFILLER_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8615_ _8617_/CLK _8615_/D vssd1 vssd1 vccd1 vccd1 _8615_/Q sky130_fd_sc_hd__dfxtp_1
X_5758_ _8006_/Q _5624_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__mux2_1
X_6934__385 _6934__385/A vssd1 vssd1 vccd1 vccd1 _8181_/CLK sky130_fd_sc_hd__inv_2
X_8546_ _8553_/CLK _8546_/D vssd1 vssd1 vccd1 vccd1 _8546_/Q sky130_fd_sc_hd__dfxtp_1
X_4709_ _4955_/S vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__buf_2
X_8477_ _8477_/CLK _8477_/D vssd1 vssd1 vccd1 vccd1 _8477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5689_ _5689_/A vssd1 vssd1 vccd1 vccd1 _8037_/D sky130_fd_sc_hd__clkbuf_1
X_7428_ _8450_/Q _7430_/B vssd1 vssd1 vccd1 vccd1 _7428_/X sky130_fd_sc_hd__or2_1
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7359_ _7376_/A vssd1 vssd1 vccd1 vccd1 _7360_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3307_ clkbuf_0__3307_/X vssd1 vssd1 vccd1 vccd1 _6759__320/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3322_ clkbuf_0__3322_/X vssd1 vssd1 vccd1 vccd1 _6824__367/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7514__3 _7516__5/A vssd1 vssd1 vccd1 vccd1 _8517_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6730_ _5991_/A _8095_/Q _6730_/S vssd1 vssd1 vccd1 vccd1 _6731_/A sky130_fd_sc_hd__mux2_1
X_4991_ _8254_/Q _4988_/X _4990_/Y _4903_/X vssd1 vssd1 vccd1 vccd1 _8254_/D sky130_fd_sc_hd__o211a_1
X_3942_ _3942_/A vssd1 vssd1 vccd1 vccd1 _8597_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3442_ clkbuf_0__3442_/X vssd1 vssd1 vccd1 vccd1 _7066_/A sky130_fd_sc_hd__clkbuf_4
X_6661_ _8267_/Q _6663_/B vssd1 vssd1 vccd1 vccd1 _6662_/A sky130_fd_sc_hd__and2_1
X_3873_ _8203_/Q vssd1 vssd1 vccd1 vccd1 _4027_/B sky130_fd_sc_hd__clkbuf_1
X_8400_ _8400_/CLK _8400_/D vssd1 vssd1 vccd1 vccd1 _8400_/Q sky130_fd_sc_hd__dfxtp_1
X_5612_ _5612_/A vssd1 vssd1 vccd1 vccd1 _8074_/D sky130_fd_sc_hd__clkbuf_1
X_8331_ _8331_/CLK _8331_/D vssd1 vssd1 vccd1 vccd1 _8331_/Q sky130_fd_sc_hd__dfxtp_1
X_5543_ _8126_/Q _4432_/A _5549_/S vssd1 vssd1 vccd1 vccd1 _5544_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3410_ _6916_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3410_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5474_ _5474_/A vssd1 vssd1 vccd1 vccd1 _8160_/D sky130_fd_sc_hd__clkbuf_1
X_8262_ _8262_/CLK _8262_/D vssd1 vssd1 vccd1 vccd1 _8262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3272_ _6680_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3272_/X sky130_fd_sc_hd__clkbuf_16
X_4425_ _4135_/X _8359_/Q _4425_/S vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__mux2_1
X_8193_ _8568_/CLK _8193_/D vssd1 vssd1 vccd1 vccd1 _8193_/Q sky130_fd_sc_hd__dfxtp_4
X_4356_ _4371_/S vssd1 vssd1 vccd1 vccd1 _4365_/S sky130_fd_sc_hd__buf_2
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _8422_/Q _4197_/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__mux2_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6026_/A vssd1 vssd1 vccd1 vccd1 _6026_/X sky130_fd_sc_hd__clkbuf_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7977_ _8270_/CLK _7977_/D vssd1 vssd1 vccd1 vccd1 _7977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6859_ _8543_/Q vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8529_ _8529_/CLK _8529_/D vssd1 vssd1 vccd1 vccd1 _8529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6789__344 _6790__345/A vssd1 vssd1 vccd1 vccd1 _8136_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_71 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_60 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_93 _8366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_82 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4210_ _8478_/Q _4209_/X _4213_/S vssd1 vssd1 vccd1 vccd1 _4211_/A sky130_fd_sc_hd__mux2_1
X_5190_ _8292_/Q _8276_/Q _8538_/Q _8308_/Q _5341_/S _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5190_/X sky130_fd_sc_hd__mux4_2
XFILLER_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4141_ _4141_/A vssd1 vssd1 vccd1 vccd1 _8492_/D sky130_fd_sc_hd__clkbuf_1
X_4072_ _8514_/Q _3934_/X _4076_/S vssd1 vssd1 vccd1 vccd1 _4073_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7900_ _8631_/CLK _7900_/D vssd1 vssd1 vccd1 vccd1 _7900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7831_ _7564_/A _7840_/C _7830_/X _7763_/A vssd1 vssd1 vccd1 vccd1 _8628_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7762_ _7762_/A vssd1 vssd1 vccd1 vccd1 _8607_/D sky130_fd_sc_hd__clkbuf_1
X_4974_ _5055_/A _4964_/X _4976_/B _4973_/Y vssd1 vssd1 vccd1 vccd1 _8259_/D sky130_fd_sc_hd__a31o_1
X_6713_ _6713_/A vssd1 vssd1 vccd1 vccd1 _8087_/D sky130_fd_sc_hd__clkbuf_1
X_3925_ _4004_/A _5383_/A _5150_/A vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__or3b_4
X_7693_ _8564_/Q _7687_/X _7692_/X _7684_/X vssd1 vssd1 vccd1 vccd1 _8563_/D sky130_fd_sc_hd__o211a_1
X_6644_ _6668_/A vssd1 vssd1 vccd1 vccd1 _6644_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3425_ clkbuf_0__3425_/X vssd1 vssd1 vccd1 vccd1 _6969__400/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5526_ _5526_/A vssd1 vssd1 vccd1 vccd1 _8134_/D sky130_fd_sc_hd__clkbuf_1
X_8314_ _8314_/CLK _8314_/D vssd1 vssd1 vccd1 vccd1 _8314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5457_ _5412_/X _8168_/Q _5459_/S vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__mux2_1
X_8245_ _8245_/CLK _8245_/D vssd1 vssd1 vccd1 vccd1 _8245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7502__169 _7502__169/A vssd1 vssd1 vccd1 vccd1 _8508_/CLK sky130_fd_sc_hd__inv_2
X_4408_ _4408_/A vssd1 vssd1 vccd1 vccd1 _8367_/D sky130_fd_sc_hd__clkbuf_1
X_8176_ _8176_/CLK _8176_/D vssd1 vssd1 vccd1 vccd1 _8176_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3255_ _6619_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3255_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5388_ _8200_/Q _5385_/X _5387_/Y _5374_/X vssd1 vssd1 vccd1 vccd1 _8200_/D sky130_fd_sc_hd__o211a_1
X_4339_ _4104_/X _8398_/Q _4347_/S vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _6009_/A vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8653__218 vssd1 vssd1 vccd1 vccd1 _8653__218/HI core0Index[5] sky130_fd_sc_hd__conb_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _4955_/S vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__clkbuf_4
X_6360_ _6483_/A vssd1 vssd1 vccd1 vccd1 _6416_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5311_ _8360_/Q _5220_/X _5249_/X _8587_/Q _5189_/A vssd1 vssd1 vccd1 vccd1 _5311_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8030_ _8030_/CLK _8030_/D vssd1 vssd1 vccd1 vccd1 _8030_/Q sky130_fd_sc_hd__dfxtp_1
X_6291_ _7716_/A _7897_/Q _6291_/S vssd1 vssd1 vccd1 vccd1 _6292_/A sky130_fd_sc_hd__mux2_1
X_5242_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__buf_2
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5173_ _5247_/A _5164_/X _5167_/X _5172_/X _5217_/A vssd1 vssd1 vccd1 vccd1 _5173_/X
+ sky130_fd_sc_hd__o221a_1
X_4124_ _4123_/X _8496_/Q _4124_/S vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4055_ _4055_/A vssd1 vssd1 vccd1 vccd1 _8521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7814_ _7814_/A _7817_/B vssd1 vssd1 vccd1 vccd1 _7814_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4957_ _8233_/Q _4807_/A _4687_/A _4956_/X vssd1 vssd1 vccd1 vccd1 _4957_/X sky130_fd_sc_hd__o211a_1
X_4888_ _8345_/Q _4829_/X _4822_/X _8058_/Q vssd1 vssd1 vccd1 vccd1 _4888_/X sky130_fd_sc_hd__a22o_1
X_7676_ _8560_/Q _7672_/A _7675_/Y vssd1 vssd1 vccd1 vccd1 _7677_/C sky130_fd_sc_hd__o21a_1
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3908_ _6077_/A _6080_/A vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__and2_1
X_7109__505 _7109__505/A vssd1 vssd1 vccd1 vccd1 _8314_/CLK sky130_fd_sc_hd__inv_2
X_6558_ _7794_/B vssd1 vssd1 vccd1 vccd1 _7778_/A sky130_fd_sc_hd__buf_2
XFILLER_118_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5509_ _8141_/Q _4489_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5510_/A sky130_fd_sc_hd__mux2_1
X_6489_ _7953_/Q _6483_/X _6474_/X _6488_/X _6472_/X vssd1 vssd1 vccd1 vccd1 _7953_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3307_ _6754_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3307_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_79_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8228_ _8228_/CLK _8228_/D vssd1 vssd1 vccd1 vccd1 _8228_/Q sky130_fd_sc_hd__dfxtp_1
X_8159_ _8159_/CLK _8159_/D vssd1 vssd1 vccd1 vccd1 _8159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6346__215 _6346__215/A vssd1 vssd1 vccd1 vccd1 _7927_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7451__127 _7453__129/A vssd1 vssd1 vccd1 vccd1 _8466_/CLK sky130_fd_sc_hd__inv_2
X_6960__392 _6963__395/A vssd1 vssd1 vccd1 vccd1 _8196_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _4450_/X _7912_/Q _5860_/S vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__mux2_1
X_7095__494 _7096__495/A vssd1 vssd1 vccd1 vccd1 _8303_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4812_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5791_ _5806_/S vssd1 vssd1 vccd1 vccd1 _5800_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4742_ _4671_/X _8268_/Q _4988_/A _4739_/X _4741_/X vssd1 vssd1 vccd1 vccd1 _4742_/X
+ sky130_fd_sc_hd__a221o_1
X_7461_ _7467_/A vssd1 vssd1 vccd1 vccd1 _7461_/X sky130_fd_sc_hd__buf_1
X_4673_ _4673_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__clkbuf_2
X_6412_ _7834_/A _6403_/X _6373_/X vssd1 vssd1 vccd1 vccd1 _6416_/B sky130_fd_sc_hd__a21oi_1
X_7392_ _8438_/Q _7384_/X _7360_/A _7250_/B vssd1 vssd1 vccd1 vccd1 _7393_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6274_ _8098_/Q _6269_/X _6270_/X _6272_/X _7887_/Q vssd1 vssd1 vccd1 vccd1 _7887_/D
+ sky130_fd_sc_hd__o32a_1
X_8013_ _8013_/CLK _8013_/D vssd1 vssd1 vccd1 vccd1 _8013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5225_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5305_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _5391_/B _5155_/X _5333_/A vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4107_ _4136_/S vssd1 vssd1 vccd1 vccd1 _4124_/S sky130_fd_sc_hd__clkbuf_4
X_5087_ _5087_/A vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3271_ clkbuf_0__3271_/X vssd1 vssd1 vccd1 vccd1 _6678__299/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4038_ _3968_/X _8528_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4039_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8675__240 vssd1 vssd1 vccd1 vccd1 _8675__240/HI partID[3] sky130_fd_sc_hd__conb_1
XFILLER_71_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6599__250 _6599__250/A vssd1 vssd1 vccd1 vccd1 _8010_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__or2_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7743__42 _7743__42/A vssd1 vssd1 vccd1 vccd1 _8593_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7659_ _7658_/X _7662_/B vssd1 vssd1 vccd1 vccd1 _7660_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput190 _6164_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3469_ clkbuf_0__3469_/X vssd1 vssd1 vccd1 vccd1 _7169__52/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _8244_/Q _4522_/X _5010_/S vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__mux2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0__3811_ clkbuf_0__3811_/X vssd1 vssd1 vccd1 vccd1 _7743__42/A sky130_fd_sc_hd__clkbuf_4
X_8659__224 vssd1 vssd1 vccd1 vccd1 _8659__224/HI core1Index[4] sky130_fd_sc_hd__conb_1
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5912_ _4209_/X _7846_/Q _5914_/S vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__mux2_1
X_6892_ _6886_/B _6886_/C _8551_/Q vssd1 vssd1 vccd1 vccd1 _7551_/B sky130_fd_sc_hd__a21o_1
X_5843_ _5843_/A vssd1 vssd1 vccd1 vccd1 _7920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8631_ _8631_/CLK _8631_/D vssd1 vssd1 vccd1 vccd1 _8631_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8562_ _8568_/CLK _8562_/D vssd1 vssd1 vccd1 vccd1 _8562_/Q sky130_fd_sc_hd__dfxtp_1
X_5774_ _7999_/Q _5593_/A _5782_/S vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4725_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__buf_2
X_8493_ _8493_/CLK _8493_/D vssd1 vssd1 vccd1 vccd1 _8493_/Q sky130_fd_sc_hd__dfxtp_1
X_4656_ _8274_/Q _4495_/X _4656_/S vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__mux2_1
X_4587_ _4447_/X _8304_/Q _4589_/S vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__mux2_1
Xinput81 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _5942_/A sky130_fd_sc_hd__clkbuf_2
Xinput70 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _7842_/A sky130_fd_sc_hd__buf_8
X_7375_ _7386_/A _7375_/B vssd1 vssd1 vccd1 vccd1 _8431_/D sky130_fd_sc_hd__nor2_1
Xinput92 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _7838_/A sky130_fd_sc_hd__buf_8
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6967__398 _6968__399/A vssd1 vssd1 vccd1 vccd1 _8202_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6783__339 _6784__340/A vssd1 vssd1 vccd1 vccd1 _8131_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _6423_/A vssd1 vssd1 vccd1 vccd1 _6257_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5208_ _8590_/Q _8339_/Q _8323_/Q _8363_/Q _5130_/X _5101_/A vssd1 vssd1 vccd1 vccd1
+ _5209_/B sky130_fd_sc_hd__mux4_2
X_6188_ _6188_/A _6188_/B vssd1 vssd1 vccd1 vccd1 _6188_/X sky130_fd_sc_hd__and2_1
X_5139_ _8390_/Q _8382_/Q _8374_/Q _8398_/Q _5138_/X _5131_/X vssd1 vssd1 vccd1 vccd1
+ _5139_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3254_ clkbuf_0__3254_/X vssd1 vssd1 vccd1 vccd1 _6618__265/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6614__261 _6616__263/A vssd1 vssd1 vccd1 vccd1 _8021_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6992__414 _6993__415/A vssd1 vssd1 vccd1 vccd1 _8220_/CLK sky130_fd_sc_hd__inv_2
X_6695__311 _6695__311/A vssd1 vssd1 vccd1 vccd1 _8079_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7168__51 _7169__52/A vssd1 vssd1 vccd1 vccd1 _8360_/CLK sky130_fd_sc_hd__inv_2
X_5490_ _5490_/A vssd1 vssd1 vccd1 vccd1 _8153_/D sky130_fd_sc_hd__clkbuf_1
X_4510_ _4532_/S vssd1 vssd1 vccd1 vccd1 _4523_/S sky130_fd_sc_hd__clkbuf_4
X_4441_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4372_ _4372_/A vssd1 vssd1 vccd1 vccd1 _8383_/D sky130_fd_sc_hd__clkbuf_1
X_6111_ _6149_/A vssd1 vssd1 vccd1 vccd1 _6126_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7091_ _7097_/A vssd1 vssd1 vccd1 vccd1 _7091_/X sky130_fd_sc_hd__buf_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6042_/A vssd1 vssd1 vccd1 vccd1 _6042_/X sky130_fd_sc_hd__clkbuf_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7993_ _7993_/CLK _7993_/D vssd1 vssd1 vccd1 vccd1 _7993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6944_ _6944_/A vssd1 vssd1 vccd1 vccd1 _8188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3656_ clkbuf_0__3656_/X vssd1 vssd1 vccd1 vccd1 _7509__175/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875_ _8632_/Q _7608_/B vssd1 vssd1 vccd1 vccd1 _6875_/Y sky130_fd_sc_hd__xnor2_1
X_8614_ _8617_/CLK _8614_/D vssd1 vssd1 vccd1 vccd1 _8614_/Q sky130_fd_sc_hd__dfxtp_1
X_5826_ _5826_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5842_/S sky130_fd_sc_hd__nor2_2
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5757_ _5757_/A vssd1 vssd1 vccd1 vccd1 _8007_/D sky130_fd_sc_hd__clkbuf_1
X_8545_ _8553_/CLK _8545_/D vssd1 vssd1 vccd1 vccd1 _8545_/Q sky130_fd_sc_hd__dfxtp_1
X_8476_ _8476_/CLK _8476_/D vssd1 vssd1 vccd1 vccd1 _8476_/Q sky130_fd_sc_hd__dfxtp_1
X_4708_ _4994_/B _4695_/X _4707_/X vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__a21o_1
X_5688_ _8037_/Q _5627_/X _5692_/S vssd1 vssd1 vccd1 vccd1 _5689_/A sky130_fd_sc_hd__mux2_1
X_7427_ _8212_/Q _7411_/A _7413_/A _7426_/X _7420_/X vssd1 vssd1 vccd1 vccd1 _8449_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_118_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4639_ _4639_/A vssd1 vssd1 vccd1 vccd1 _8282_/D sky130_fd_sc_hd__clkbuf_1
X_7358_ _7358_/A _7358_/B vssd1 vssd1 vccd1 vccd1 _7376_/A sky130_fd_sc_hd__or2_1
XFILLER_116_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7289_ _7361_/A _7361_/B _6872_/A vssd1 vssd1 vccd1 vccd1 _7289_/Y sky130_fd_sc_hd__a21oi_1
X_6309_ _8416_/Q vssd1 vssd1 vccd1 vccd1 _7407_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6807__353 _6809__355/A vssd1 vssd1 vccd1 vccd1 _8148_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _4996_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4990_/Y sky130_fd_sc_hd__nand2_1
X_3941_ _8597_/Q _3940_/X _3941_/S vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3441_ clkbuf_0__3441_/X vssd1 vssd1 vccd1 vccd1 _7037__450/A sky130_fd_sc_hd__clkbuf_4
X_3872_ _8577_/Q vssd1 vssd1 vccd1 vccd1 _3872_/X sky130_fd_sc_hd__buf_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6660_ _6660_/A vssd1 vssd1 vccd1 vccd1 _8053_/D sky130_fd_sc_hd__clkbuf_1
X_5611_ _5610_/X _8074_/Q _5617_/S vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__mux2_1
X_5542_ _5542_/A vssd1 vssd1 vccd1 vccd1 _8127_/D sky130_fd_sc_hd__clkbuf_1
X_8330_ _8330_/CLK _8330_/D vssd1 vssd1 vccd1 vccd1 _8330_/Q sky130_fd_sc_hd__dfxtp_1
X_5473_ _4435_/X _8160_/Q _5477_/S vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__mux2_1
X_8261_ _8261_/CLK _8261_/D vssd1 vssd1 vccd1 vccd1 _8261_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3271_ _6674_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3271_/X sky130_fd_sc_hd__clkbuf_16
X_4424_ _4424_/A vssd1 vssd1 vccd1 vccd1 _8360_/D sky130_fd_sc_hd__clkbuf_1
X_8192_ _8568_/CLK _8192_/D vssd1 vssd1 vccd1 vccd1 _8192_/Q sky130_fd_sc_hd__dfxtp_4
X_4355_ _4355_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4371_/S sky130_fd_sc_hd__or2_2
XFILLER_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4286_ _4286_/A vssd1 vssd1 vccd1 vccd1 _8423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6025_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6026_/A sky130_fd_sc_hd__and2_1
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6940__390 _6940__390/A vssd1 vssd1 vccd1 vccd1 _8186_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7976_ _8617_/CLK _7976_/D vssd1 vssd1 vccd1 vccd1 _7976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6858_ _8544_/Q vssd1 vssd1 vccd1 vccd1 _7607_/A sky130_fd_sc_hd__clkbuf_2
X_5809_ _5824_/S vssd1 vssd1 vccd1 vccd1 _5818_/S sky130_fd_sc_hd__buf_2
XFILLER_50_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8528_ _8528_/CLK _8528_/D vssd1 vssd1 vccd1 vccd1 _8528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8459_ _8459_/CLK _8459_/D vssd1 vssd1 vccd1 vccd1 _8459_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3469_ _7167_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3469_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_50 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7158__545 _7158__545/A vssd1 vssd1 vccd1 vccd1 _8354_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_61 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_72 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_94 _6303_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_83 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4140_ _8492_/Q _3872_/X _4148_/S vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7102__500 _7102__500/A vssd1 vssd1 vccd1 vccd1 _8309_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _8515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7059__465 _7059__465/A vssd1 vssd1 vccd1 vccd1 _8274_/CLK sky130_fd_sc_hd__inv_2
X_7830_ _7719_/A _7723_/B _7826_/X vssd1 vssd1 vccd1 vccd1 _7830_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7761_ _7763_/A _8249_/Q vssd1 vssd1 vccd1 vccd1 _7762_/A sky130_fd_sc_hd__and2_1
X_4973_ _5772_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _4973_/Y sky130_fd_sc_hd__nor2_1
X_6712_ _7796_/A _8087_/Q _6712_/S vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__mux2_1
X_3924_ _7714_/A _5916_/A _4164_/C _6193_/A vssd1 vssd1 vccd1 vccd1 _5150_/A sky130_fd_sc_hd__a31oi_4
X_7692_ _8563_/Q _7698_/B vssd1 vssd1 vccd1 vccd1 _7692_/X sky130_fd_sc_hd__or2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6593__245 _6593__245/A vssd1 vssd1 vccd1 vccd1 _8005_/CLK sky130_fd_sc_hd__inv_2
X_5525_ _8134_/Q _4432_/A _5531_/S vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__mux2_1
X_8313_ _8313_/CLK _8313_/D vssd1 vssd1 vccd1 vccd1 _8313_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_22_wb_clk_i _6197_/A vssd1 vssd1 vccd1 vccd1 _8608_/CLK sky130_fd_sc_hd__clkbuf_16
X_5456_ _5456_/A vssd1 vssd1 vccd1 vccd1 _8169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8244_ _8244_/CLK _8244_/D vssd1 vssd1 vccd1 vccd1 _8244_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3254_ _6613_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3254_/X sky130_fd_sc_hd__clkbuf_16
X_4407_ _4135_/X _8367_/Q _4407_/S vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8175_ _8175_/CLK _8175_/D vssd1 vssd1 vccd1 vccd1 _8175_/Q sky130_fd_sc_hd__dfxtp_1
X_5387_ _5393_/A _5387_/B vssd1 vssd1 vccd1 vccd1 _5387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4338_ _4353_/S vssd1 vssd1 vccd1 vccd1 _4347_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4269_ _4269_/A vssd1 vssd1 vccd1 vccd1 _8458_/D sky130_fd_sc_hd__clkbuf_1
X_6008_ _6008_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__or2_1
XFILLER_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8639__255 vssd1 vssd1 vccd1 vccd1 partID[8] _8639__255/LO sky130_fd_sc_hd__conb_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7959_ _8452_/CLK _7959_/D vssd1 vssd1 vccd1 vccd1 _7959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5310_ _8320_/Q _8336_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5310_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6290_ _6290_/A vssd1 vssd1 vccd1 vccd1 _7896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5241_ _5233_/X _5235_/X _5240_/X vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5172_ _5135_/X _5170_/X _5171_/X vssd1 vssd1 vccd1 vccd1 _5172_/X sky130_fd_sc_hd__a21o_1
X_4123_ _4441_/A vssd1 vssd1 vccd1 vccd1 _4123_/X sky130_fd_sc_hd__clkbuf_2
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4054_ _3965_/X _8521_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7813_ _7811_/Y _7812_/Y _7800_/X vssd1 vssd1 vccd1 vccd1 _8623_/D sky130_fd_sc_hd__a21oi_1
XFILLER_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6972__401 _6975__404/A vssd1 vssd1 vccd1 vccd1 _8205_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4956_ _8172_/Q _4856_/A _4860_/A _4955_/X vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__o22a_1
X_7033__446 _7034__447/A vssd1 vssd1 vccd1 vccd1 _8253_/CLK sky130_fd_sc_hd__inv_2
X_4887_ _4869_/X _4877_/X _4880_/X _4886_/X _4990_/B vssd1 vssd1 vccd1 vccd1 _4887_/X
+ sky130_fd_sc_hd__o311a_1
X_3907_ _3907_/A _3907_/B _3907_/C _3907_/D vssd1 vssd1 vccd1 vccd1 _6080_/A sky130_fd_sc_hd__nor4_4
X_7675_ _8560_/Q _7672_/A _7681_/A vssd1 vssd1 vccd1 vccd1 _7675_/Y sky130_fd_sc_hd__a21oi_1
X_7522__10 _7519__7/A vssd1 vssd1 vccd1 vccd1 _8524_/CLK sky130_fd_sc_hd__inv_2
X_6557_ _6368_/A _6562_/B _6501_/A vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__o21ai_1
X_5508_ _5508_/A vssd1 vssd1 vccd1 vccd1 _8142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6488_ _7053_/A _6490_/B _6492_/C vssd1 vssd1 vccd1 vccd1 _6488_/X sky130_fd_sc_hd__and3_1
X_5439_ _5412_/X _8176_/Q _5441_/S vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__mux2_1
X_8227_ _8227_/CLK _8227_/D vssd1 vssd1 vccd1 vccd1 _8227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8158_ _8158_/CLK _8158_/D vssd1 vssd1 vccd1 vccd1 _8158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8089_ _8622_/CLK _8089_/D vssd1 vssd1 vccd1 vccd1 _8089_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _8251_/Q vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__inv_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5790_ _5790_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5806_/S sky130_fd_sc_hd__nor2_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4741_/A vssd1 vssd1 vccd1 vccd1 _4741_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4672_ _4672_/A _6647_/B vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__nor2_2
X_6411_ _8630_/Q vssd1 vssd1 vccd1 vccd1 _7834_/A sky130_fd_sc_hd__buf_4
X_7391_ _7398_/A _7391_/B vssd1 vssd1 vccd1 vccd1 _8437_/D sky130_fd_sc_hd__nor2_1
X_6273_ _8097_/Q _6269_/X _6270_/X _6272_/X _7886_/Q vssd1 vssd1 vccd1 vccd1 _7886_/D
+ sky130_fd_sc_hd__o32a_1
X_8012_ _8012_/CLK _8012_/D vssd1 vssd1 vccd1 vccd1 _8012_/Q sky130_fd_sc_hd__dfxtp_1
X_5224_ _5232_/A vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5155_ _8523_/Q _8515_/Q _7918_/Q _8531_/Q _5122_/X _5123_/X vssd1 vssd1 vccd1 vccd1
+ _5155_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4106_ _4573_/A _4241_/B vssd1 vssd1 vccd1 vccd1 _4136_/S sky130_fd_sc_hd__or2_2
X_5086_ _8200_/Q _5144_/B vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__xor2_2
Xclkbuf_1_0_0__3270_ clkbuf_0__3270_/X vssd1 vssd1 vccd1 vccd1 _6672__294/A sky130_fd_sc_hd__clkbuf_4
X_4037_ _4037_/A vssd1 vssd1 vccd1 vccd1 _8529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7115__510 _7115__510/A vssd1 vssd1 vccd1 vccd1 _8319_/CLK sky130_fd_sc_hd__inv_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _5988_/A vssd1 vssd1 vccd1 vccd1 _5988_/X sky130_fd_sc_hd__clkbuf_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4939_ _4934_/X _4935_/X _4938_/X _4992_/B vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__a211o_1
X_7658_ _6835_/B _7642_/X _7647_/X _7546_/B vssd1 vssd1 vccd1 vccd1 _7658_/X sky130_fd_sc_hd__o22a_1
X_7589_ _7589_/A _7589_/B vssd1 vssd1 vccd1 vccd1 _7589_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7165_/A
+ sky130_fd_sc_hd__clkbuf_16
X_6352__220 _6352__220/A vssd1 vssd1 vccd1 vccd1 _7932_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput180 _6127_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput191 _6167_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__buf_2
XFILLER_102_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6979__407 _6982__410/A vssd1 vssd1 vccd1 vccd1 _8211_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3468_ clkbuf_0__3468_/X vssd1 vssd1 vccd1 vccd1 _7173_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7195__74 _7196__75/A vssd1 vssd1 vccd1 vccd1 _8383_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3810_ clkbuf_0__3810_/X vssd1 vssd1 vccd1 vccd1 _7740__40/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _5911_/A vssd1 vssd1 vccd1 vccd1 _7847_/D sky130_fd_sc_hd__clkbuf_1
X_6891_ _6891_/A _6891_/B _6891_/C _6852_/B vssd1 vssd1 vccd1 vccd1 _7551_/A sky130_fd_sc_hd__or4b_1
X_5842_ _7920_/Q _4450_/A _5842_/S vssd1 vssd1 vccd1 vccd1 _5843_/A sky130_fd_sc_hd__mux2_1
X_8630_ _8630_/CLK _8630_/D vssd1 vssd1 vccd1 vccd1 _8630_/Q sky130_fd_sc_hd__dfxtp_1
X_5773_ _5788_/S vssd1 vssd1 vccd1 vccd1 _5782_/S sky130_fd_sc_hd__buf_2
X_8561_ _8561_/CLK _8561_/D vssd1 vssd1 vccd1 vccd1 _8561_/Q sky130_fd_sc_hd__dfxtp_1
X_4724_ _4724_/A vssd1 vssd1 vccd1 vccd1 _4756_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8492_ _8492_/CLK _8492_/D vssd1 vssd1 vccd1 vccd1 _8492_/Q sky130_fd_sc_hd__dfxtp_1
X_4655_ _4655_/A vssd1 vssd1 vccd1 vccd1 _8275_/D sky130_fd_sc_hd__clkbuf_1
X_4586_ _4586_/A vssd1 vssd1 vccd1 vccd1 _8305_/D sky130_fd_sc_hd__clkbuf_1
Xinput60 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _3903_/B sky130_fd_sc_hd__clkbuf_1
Xinput71 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _7812_/A sky130_fd_sc_hd__buf_4
Xinput82 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _5985_/A sky130_fd_sc_hd__clkbuf_2
X_7374_ _8431_/Q _7368_/X _7360_/X _7373_/Y vssd1 vssd1 vccd1 vccd1 _7375_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput93 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _6006_/A sky130_fd_sc_hd__buf_4
XFILLER_103_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6256_ _6249_/X _8087_/Q _6253_/X _6255_/X _7876_/Q vssd1 vssd1 vccd1 vccd1 _7876_/D
+ sky130_fd_sc_hd__o32a_1
X_5207_ _5205_/X _5206_/X _5246_/S vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__mux2_1
X_6187_ _7891_/Q _6175_/X _6176_/X _6186_/X _6101_/A vssd1 vssd1 vccd1 vccd1 _6187_/X
+ sky130_fd_sc_hd__o221a_1
X_5138_ _5258_/S vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__buf_2
XFILLER_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5069_ _5069_/A vssd1 vssd1 vccd1 vccd1 _8219_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3253_ clkbuf_0__3253_/X vssd1 vssd1 vccd1 vccd1 _6611__259/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7046__456 _7050__460/A vssd1 vssd1 vccd1 vccd1 _8263_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3466_ clkbuf_0__3466_/X vssd1 vssd1 vccd1 vccd1 _7162__548/A sky130_fd_sc_hd__clkbuf_16
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4440_/A vssd1 vssd1 vccd1 vccd1 _8355_/D sky130_fd_sc_hd__clkbuf_1
X_4371_ _4135_/X _8383_/Q _4371_/S vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__mux2_1
X_6110_ _7944_/Q input33/X _6125_/S vssd1 vssd1 vccd1 vccd1 _6110_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6041_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6042_/A sky130_fd_sc_hd__and2_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7992_ _7992_/CLK _7992_/D vssd1 vssd1 vccd1 vccd1 _7992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6943_ _8562_/Q _6947_/B vssd1 vssd1 vccd1 vccd1 _6944_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3655_ clkbuf_0__3655_/X vssd1 vssd1 vccd1 vccd1 _7502__169/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6874_ _8544_/Q _6876_/A vssd1 vssd1 vccd1 vccd1 _7608_/B sky130_fd_sc_hd__xor2_4
X_5825_ _5825_/A vssd1 vssd1 vccd1 vccd1 _7928_/D sky130_fd_sc_hd__clkbuf_1
X_8613_ _8617_/CLK _8613_/D vssd1 vssd1 vccd1 vccd1 _8613_/Q sky130_fd_sc_hd__dfxtp_1
X_5756_ _8007_/Q _5619_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5757_/A sky130_fd_sc_hd__mux2_1
X_7464__138 _7466__140/A vssd1 vssd1 vccd1 vccd1 _8477_/CLK sky130_fd_sc_hd__inv_2
X_8544_ _8553_/CLK _8544_/D vssd1 vssd1 vccd1 vccd1 _8544_/Q sky130_fd_sc_hd__dfxtp_2
X_8475_ _8475_/CLK _8475_/D vssd1 vssd1 vccd1 vccd1 _8475_/Q sky130_fd_sc_hd__dfxtp_1
X_4707_ _4699_/X _4703_/X _4706_/X vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__a21o_1
X_5687_ _5687_/A vssd1 vssd1 vccd1 vccd1 _8038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4638_ _4469_/X _8282_/Q _4638_/S vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__mux2_1
X_7426_ _8449_/Q _7430_/B vssd1 vssd1 vccd1 vccd1 _7426_/X sky130_fd_sc_hd__or2_1
XFILLER_118_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7357_ _7371_/A _7357_/B vssd1 vssd1 vccd1 vccd1 _8426_/D sky130_fd_sc_hd__nor2_1
X_4569_ _8312_/Q _4528_/X _4571_/S vssd1 vssd1 vccd1 vccd1 _4570_/A sky130_fd_sc_hd__mux2_1
X_6308_ _6308_/A vssd1 vssd1 vccd1 vccd1 _7902_/D sky130_fd_sc_hd__clkbuf_1
X_7288_ _8631_/Q _7361_/A _7361_/B vssd1 vssd1 vccd1 vccd1 _7288_/X sky130_fd_sc_hd__and3_1
XFILLER_89_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6239_ _6232_/X _7898_/Q _6236_/X _6238_/X _7866_/Q vssd1 vssd1 vccd1 vccd1 _7866_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6759__320 _6759__320/A vssd1 vssd1 vccd1 vccd1 _8112_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ _8573_/Q vssd1 vssd1 vccd1 vccd1 _3940_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3440_ clkbuf_0__3440_/X vssd1 vssd1 vccd1 vccd1 _7028__442/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5610_ _5610_/A vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__buf_2
X_5541_ _8127_/Q _4427_/A _5549_/S vssd1 vssd1 vccd1 vccd1 _5542_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8260_ _8260_/CLK _8260_/D vssd1 vssd1 vccd1 vccd1 _8260_/Q sky130_fd_sc_hd__dfxtp_1
X_5472_ _5472_/A vssd1 vssd1 vccd1 vccd1 _8161_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3270_ _6668_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3270_/X sky130_fd_sc_hd__clkbuf_16
X_4423_ _4131_/X _8360_/Q _4425_/S vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__mux2_1
X_8191_ _8568_/CLK _8191_/D vssd1 vssd1 vccd1 vccd1 _8191_/Q sky130_fd_sc_hd__dfxtp_2
X_4354_ _4354_/A vssd1 vssd1 vccd1 vccd1 _8391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7073_ _7079_/A vssd1 vssd1 vccd1 vccd1 _7073_/X sky130_fd_sc_hd__buf_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _6024_/A vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__clkbuf_1
X_4285_ _8423_/Q _4194_/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7975_ _8617_/CLK _7975_/D vssd1 vssd1 vccd1 vccd1 _7975_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6857_ _8545_/Q vssd1 vssd1 vccd1 vccd1 _7610_/A sky130_fd_sc_hd__buf_2
X_5808_ _5808_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5824_/S sky130_fd_sc_hd__or2_2
XFILLER_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5739_ _5739_/A vssd1 vssd1 vccd1 vccd1 _8015_/D sky130_fd_sc_hd__clkbuf_1
X_8527_ _8527_/CLK _8527_/D vssd1 vssd1 vccd1 vccd1 _8527_/Q sky130_fd_sc_hd__dfxtp_1
X_8458_ _8458_/CLK _8458_/D vssd1 vssd1 vccd1 vccd1 _8458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8389_ _8389_/CLK _8389_/D vssd1 vssd1 vccd1 vccd1 _8389_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3468_ _7166_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3468_/X sky130_fd_sc_hd__clkbuf_16
X_7409_ _8443_/Q _7420_/A _7405_/Y _7408_/X vssd1 vssd1 vccd1 vccd1 _8443_/D sky130_fd_sc_hd__a31o_1
XINSDIODE2_51 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_40 _6182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_84 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_73 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_62 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6917__371 _6921__375/A vssd1 vssd1 vccd1 vccd1 _8167_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _8515_/Q _3931_/X _4076_/S vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6627__272 _6630__275/A vssd1 vssd1 vccd1 vccd1 _8032_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7760_ _7760_/A vssd1 vssd1 vccd1 vccd1 _7763_/A sky130_fd_sc_hd__buf_2
X_4972_ _5055_/A _5055_/B _5055_/C vssd1 vssd1 vccd1 vccd1 _5898_/B sky130_fd_sc_hd__nand3b_4
XFILLER_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6711_ _6711_/A vssd1 vssd1 vccd1 vccd1 _8086_/D sky130_fd_sc_hd__clkbuf_1
X_3923_ _7790_/B _6384_/A _3923_/C _7774_/B vssd1 vssd1 vccd1 vccd1 _4164_/C sky130_fd_sc_hd__nor4_2
X_7691_ _8563_/Q _7687_/X _7690_/X _7684_/X vssd1 vssd1 vccd1 vccd1 _8562_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8312_ _8312_/CLK _8312_/D vssd1 vssd1 vccd1 vccd1 _8312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5524_ _5524_/A vssd1 vssd1 vccd1 vccd1 _8135_/D sky130_fd_sc_hd__clkbuf_1
X_5455_ _5408_/X _8169_/Q _5459_/S vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3322_ _6822_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3322_/X sky130_fd_sc_hd__clkbuf_16
X_8243_ _8243_/CLK _8243_/D vssd1 vssd1 vccd1 vccd1 _8243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3253_ _6607_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3253_/X sky130_fd_sc_hd__clkbuf_16
X_4406_ _4406_/A vssd1 vssd1 vccd1 vccd1 _8368_/D sky130_fd_sc_hd__clkbuf_1
X_8174_ _8174_/CLK _8174_/D vssd1 vssd1 vccd1 vccd1 _8174_/Q sky130_fd_sc_hd__dfxtp_1
X_5386_ _5386_/A vssd1 vssd1 vccd1 vccd1 _5393_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4337_ _4573_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4353_/S sky130_fd_sc_hd__or2_2
X_4268_ _8458_/Q _4197_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4269_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6007_ _6007_/A vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4199_ _4199_/A vssd1 vssd1 vccd1 vccd1 _8482_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _8612_/CLK _7958_/D vssd1 vssd1 vccd1 vccd1 _7958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6909_/A _6909_/B _7593_/A _7688_/A vssd1 vssd1 vccd1 vccd1 _6911_/B sky130_fd_sc_hd__and4_1
X_7889_ _8561_/CLK _7889_/D vssd1 vssd1 vccd1 vccd1 _7889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7164__550 _7164__550/A vssd1 vssd1 vccd1 vccd1 _8359_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _8306_/Q _5236_/X _5238_/X _8290_/Q _5239_/X vssd1 vssd1 vccd1 vccd1 _5240_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7065__470 _7065__470/A vssd1 vssd1 vccd1 vccd1 _8279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _8573_/Q vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__buf_2
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4053_ _4053_/A vssd1 vssd1 vccd1 vccd1 _8522_/D sky130_fd_sc_hd__clkbuf_1
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7812_ _7812_/A _7812_/B vssd1 vssd1 vccd1 vccd1 _7812_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4955_ _7992_/Q _8164_/Q _4955_/S vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3906_ _3906_/A _3906_/B _3906_/C vssd1 vssd1 vccd1 vccd1 _3907_/D sky130_fd_sc_hd__or3_2
X_4886_ _4881_/X _4882_/X _4885_/X _4992_/B vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__a211o_1
X_7674_ _7672_/A _7671_/Y _7673_/X _7601_/X vssd1 vssd1 vccd1 vccd1 _8559_/D sky130_fd_sc_hd__o211a_1
X_6625_ _6625_/A vssd1 vssd1 vccd1 vccd1 _6625_/X sky130_fd_sc_hd__buf_1
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6556_ _6303_/C _7794_/B _6494_/B vssd1 vssd1 vccd1 vccd1 _6562_/B sky130_fd_sc_hd__a21oi_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5507_ _8142_/Q _4486_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5508_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8226_ _8226_/CLK _8226_/D vssd1 vssd1 vccd1 vccd1 _8226_/Q sky130_fd_sc_hd__dfxtp_1
X_6487_ _8616_/Q vssd1 vssd1 vccd1 vccd1 _7053_/A sky130_fd_sc_hd__buf_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5438_ _5438_/A vssd1 vssd1 vccd1 vccd1 _8177_/D sky130_fd_sc_hd__clkbuf_1
X_8157_ _8157_/CLK _8157_/D vssd1 vssd1 vccd1 vccd1 _8157_/Q sky130_fd_sc_hd__dfxtp_1
X_5369_ _8206_/Q _5147_/A _4064_/B _5303_/X vssd1 vssd1 vccd1 vccd1 _8206_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8088_ _8622_/CLK _8088_/D vssd1 vssd1 vccd1 vccd1 _8088_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7039_ _7051_/A vssd1 vssd1 vccd1 vccd1 _7039_/X sky130_fd_sc_hd__buf_1
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4740_ _8269_/Q _6647_/B vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__and2_1
XFILLER_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4671_ _4672_/A vssd1 vssd1 vccd1 vccd1 _4671_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7390_ _8437_/Q _7384_/X _7360_/A _7304_/B vssd1 vssd1 vccd1 vccd1 _7391_/B sky130_fd_sc_hd__o2bb2a_1
X_6410_ _6483_/A vssd1 vssd1 vccd1 vccd1 _6410_/X sky130_fd_sc_hd__clkbuf_2
X_6341_ _6341_/A vssd1 vssd1 vccd1 vccd1 _6341_/X sky130_fd_sc_hd__buf_1
XFILLER_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6272_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6272_/X sky130_fd_sc_hd__clkbuf_2
X_5223_ _5223_/A _5237_/A vssd1 vssd1 vccd1 vccd1 _5232_/A sky130_fd_sc_hd__nand2_1
X_8011_ _8011_/CLK _8011_/D vssd1 vssd1 vccd1 vccd1 _8011_/Q sky130_fd_sc_hd__dfxtp_1
X_5154_ _8491_/Q _8475_/Q _8467_/Q _8499_/Q _5324_/S _5101_/X vssd1 vssd1 vccd1 vccd1
+ _5154_/X sky130_fd_sc_hd__mux4_2
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ _4299_/A _5373_/A _5376_/A vssd1 vssd1 vccd1 vccd1 _4241_/B sky130_fd_sc_hd__nand3_4
XFILLER_111_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5085_ _5085_/A vssd1 vssd1 vccd1 vccd1 _5144_/B sky130_fd_sc_hd__buf_2
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _3965_/X _8529_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__mux2_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7728__30 _7728__30/A vssd1 vssd1 vccd1 vccd1 _8581_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5987_ _5987_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5988_/A sky130_fd_sc_hd__or2_4
X_4938_ _8008_/Q _4807_/A _4723_/A _4937_/X vssd1 vssd1 vccd1 vccd1 _4938_/X sky130_fd_sc_hd__o211a_1
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6753__315 _6753__315/A vssd1 vssd1 vccd1 vccd1 _8107_/CLK sky130_fd_sc_hd__inv_2
X_4869_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7657_ _7657_/A vssd1 vssd1 vccd1 vccd1 _8555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7588_ _7588_/A _7588_/B _7588_/C vssd1 vssd1 vccd1 vccd1 _7588_/X sky130_fd_sc_hd__and3_1
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539_ _6550_/A vssd1 vssd1 vccd1 vccd1 _6548_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput170 _5929_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8209_ _8209_/CLK _8209_/D vssd1 vssd1 vccd1 vccd1 _8209_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput181 _6132_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput192 _6169_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3467_ clkbuf_0__3467_/X vssd1 vssd1 vccd1 vccd1 _7479_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5910_ _4206_/X _7847_/Q _5914_/S vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6890_ _8550_/Q _8549_/Q vssd1 vssd1 vccd1 vccd1 _6891_/B sky130_fd_sc_hd__nand2_1
X_5841_ _5841_/A vssd1 vssd1 vccd1 vccd1 _7921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5772_ _5772_/A _5772_/B vssd1 vssd1 vccd1 vccd1 _5788_/S sky130_fd_sc_hd__nor2_2
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8560_ _8561_/CLK _8560_/D vssd1 vssd1 vccd1 vccd1 _8560_/Q sky130_fd_sc_hd__dfxtp_1
X_8491_ _8491_/CLK _8491_/D vssd1 vssd1 vccd1 vccd1 _8491_/Q sky130_fd_sc_hd__dfxtp_1
X_4723_ _4723_/A _4723_/B vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__and2_1
X_7511_ _7529_/A vssd1 vssd1 vccd1 vccd1 _7511_/X sky130_fd_sc_hd__buf_1
X_7442_ _7442_/A vssd1 vssd1 vccd1 vccd1 _7442_/X sky130_fd_sc_hd__buf_1
X_4654_ _8275_/Q _4492_/X _4656_/S vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4585_ _4444_/X _8305_/Q _4589_/S vssd1 vssd1 vccd1 vccd1 _4586_/A sky130_fd_sc_hd__mux2_1
Xinput50 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _3902_/C sky130_fd_sc_hd__clkbuf_1
Xinput72 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _7809_/A sky130_fd_sc_hd__buf_4
Xinput61 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__clkbuf_1
X_7373_ _7373_/A _7373_/B vssd1 vssd1 vccd1 vccd1 _7373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput94 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _6008_/A sky130_fd_sc_hd__buf_4
Xinput83 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6255_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6255_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5206_ _8387_/Q _8379_/Q _8371_/Q _8395_/Q _5138_/X _5123_/A vssd1 vssd1 vccd1 vccd1
+ _5206_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6186_ _6186_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6186_/X sky130_fd_sc_hd__and2_1
X_5137_ _5135_/X _5136_/X _5264_/A vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3321_ clkbuf_0__3321_/X vssd1 vssd1 vccd1 vccd1 _6819__363/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5068_ _4472_/X _8219_/Q _5072_/S vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7078__480 _7078__480/A vssd1 vssd1 vccd1 vccd1 _8289_/CLK sky130_fd_sc_hd__inv_2
X_4019_ _8535_/Q _3943_/X _4023_/S vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3252_ clkbuf_0__3252_/X vssd1 vssd1 vccd1 vccd1 _6603__252/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7709_ _7709_/A vssd1 vssd1 vccd1 vccd1 _8570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6621__267 _6621__267/A vssd1 vssd1 vccd1 vccd1 _8027_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6324__197 _6325__198/A vssd1 vssd1 vccd1 vccd1 _7909_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4370_/A vssd1 vssd1 vccd1 vccd1 _8384_/D sky130_fd_sc_hd__clkbuf_1
X_8665__230 vssd1 vssd1 vccd1 vccd1 _8665__230/HI manufacturerID[2] sky130_fd_sc_hd__conb_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A vssd1 vssd1 vccd1 vccd1 _6040_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7991_ _7991_/CLK _7991_/D vssd1 vssd1 vccd1 vccd1 _7991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3654_ clkbuf_0__3654_/X vssd1 vssd1 vccd1 vccd1 _7497__165/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8554_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6873_ _7611_/A _7611_/B _6872_/A vssd1 vssd1 vccd1 vccd1 _6873_/Y sky130_fd_sc_hd__a21oi_1
X_5824_ _5616_/X _7928_/Q _5824_/S vssd1 vssd1 vccd1 vccd1 _5825_/A sky130_fd_sc_hd__mux2_1
X_8612_ _8612_/CLK _8612_/D vssd1 vssd1 vccd1 vccd1 _8612_/Q sky130_fd_sc_hd__dfxtp_1
X_5755_ _5770_/S vssd1 vssd1 vccd1 vccd1 _5764_/S sky130_fd_sc_hd__buf_2
X_8543_ _8553_/CLK _8543_/D vssd1 vssd1 vccd1 vccd1 _8543_/Q sky130_fd_sc_hd__dfxtp_1
X_8474_ _8474_/CLK _8474_/D vssd1 vssd1 vccd1 vccd1 _8474_/Q sky130_fd_sc_hd__dfxtp_1
X_5686_ _8038_/Q _5624_/X _5692_/S vssd1 vssd1 vccd1 vccd1 _5687_/A sky130_fd_sc_hd__mux2_1
X_7174__56 _7178__60/A vssd1 vssd1 vccd1 vccd1 _8365_/CLK sky130_fd_sc_hd__inv_2
X_4706_ _4841_/A vssd1 vssd1 vccd1 vccd1 _4706_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4637_ _4637_/A vssd1 vssd1 vccd1 vccd1 _8283_/D sky130_fd_sc_hd__clkbuf_1
X_7425_ _8211_/Q _7411_/A _7413_/X _7424_/X _7420_/X vssd1 vssd1 vccd1 vccd1 _8448_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_116_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4568_ _4568_/A vssd1 vssd1 vccd1 vccd1 _8313_/D sky130_fd_sc_hd__clkbuf_1
X_7356_ _7349_/B _7292_/B _7350_/Y _7352_/X _8426_/Q vssd1 vssd1 vccd1 vccd1 _7357_/B
+ sky130_fd_sc_hd__a32oi_1
X_4499_ _8337_/Q _4498_/X _4505_/S vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__mux2_1
X_6307_ _6306_/X _6307_/B vssd1 vssd1 vccd1 vccd1 _6308_/A sky130_fd_sc_hd__and2b_1
X_7287_ _8426_/Q _8425_/Q _8427_/Q vssd1 vssd1 vccd1 vccd1 _7361_/B sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1_0__3019_ clkbuf_0__3019_/X vssd1 vssd1 vccd1 vccd1 _6216__189/A sky130_fd_sc_hd__clkbuf_4
X_6238_ _6247_/A vssd1 vssd1 vccd1 vccd1 _6238_/X sky130_fd_sc_hd__clkbuf_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _7884_/Q _6159_/X _6163_/X _6168_/X _6157_/X vssd1 vssd1 vccd1 vccd1 _6169_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7052__461 _7059__465/A vssd1 vssd1 vccd1 vccd1 _8268_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6204__179 _6204__179/A vssd1 vssd1 vccd1 vccd1 _7848_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8649__214 vssd1 vssd1 vccd1 vccd1 _8649__214/HI core0Index[1] sky130_fd_sc_hd__conb_1
XFILLER_5_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7233__104 _7234__105/A vssd1 vssd1 vccd1 vccd1 _8413_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5540_ _5555_/S vssd1 vssd1 vccd1 vccd1 _5549_/S sky130_fd_sc_hd__buf_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5471_ _4432_/X _8161_/Q _5477_/S vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__mux2_1
X_6814__359 _6815__360/A vssd1 vssd1 vccd1 vccd1 _8154_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7210_ _7210_/A vssd1 vssd1 vccd1 vccd1 _7210_/X sky130_fd_sc_hd__buf_1
X_4422_ _4422_/A vssd1 vssd1 vccd1 vccd1 _8361_/D sky130_fd_sc_hd__clkbuf_1
X_8190_ _8568_/CLK _8190_/D vssd1 vssd1 vccd1 vccd1 _8190_/Q sky130_fd_sc_hd__dfxtp_1
X_7141_ _7159_/A vssd1 vssd1 vccd1 vccd1 _7141_/X sky130_fd_sc_hd__buf_1
X_4353_ _4135_/X _8391_/Q _4353_/S vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__mux2_1
X_4284_ _4284_/A vssd1 vssd1 vccd1 vccd1 _8424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7072_ _7072_/A vssd1 vssd1 vccd1 vccd1 _7072_/X sky130_fd_sc_hd__buf_1
X_6023_ _6023_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__and2_1
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7470__143 _7472__145/A vssd1 vssd1 vccd1 vccd1 _8482_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7974_ _8608_/CLK _7974_/D vssd1 vssd1 vccd1 vccd1 _7974_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3020_ clkbuf_0__3020_/X vssd1 vssd1 vccd1 vccd1 _6321__195/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6856_ _8549_/Q vssd1 vssd1 vccd1 vccd1 _6861_/A sky130_fd_sc_hd__inv_2
X_5807_ _5807_/A vssd1 vssd1 vccd1 vccd1 _7984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _3999_/A vssd1 vssd1 vccd1 vccd1 _8579_/D sky130_fd_sc_hd__clkbuf_1
X_5738_ _8015_/Q _5619_/X _5746_/S vssd1 vssd1 vccd1 vccd1 _5739_/A sky130_fd_sc_hd__mux2_1
X_8526_ _8526_/CLK _8526_/D vssd1 vssd1 vccd1 vccd1 _8526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5669_/A vssd1 vssd1 vccd1 vccd1 _8046_/D sky130_fd_sc_hd__clkbuf_1
X_8457_ _8457_/CLK _8457_/D vssd1 vssd1 vccd1 vccd1 _8457_/Q sky130_fd_sc_hd__dfxtp_1
X_8388_ _8388_/CLK _8388_/D vssd1 vssd1 vccd1 vccd1 _8388_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3467_ _7165_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3467_/X sky130_fd_sc_hd__clkbuf_16
X_7408_ _7432_/S _7408_/B _7408_/C vssd1 vssd1 vccd1 vccd1 _7408_/X sky130_fd_sc_hd__and3_1
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_41 _6182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_52 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_30 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_85 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_63 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_74 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7343__110 _7343__110/A vssd1 vssd1 vccd1 vccd1 _8421_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924__376 _6927__379/A vssd1 vssd1 vccd1 vccd1 _8172_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4971_ _5808_/A vssd1 vssd1 vccd1 vccd1 _5772_/A sky130_fd_sc_hd__buf_4
X_6710_ _7799_/A _8086_/Q _6712_/S vssd1 vssd1 vccd1 vccd1 _6711_/A sky130_fd_sc_hd__mux2_1
X_3922_ _6505_/B _6366_/B _6366_/C _6366_/D vssd1 vssd1 vccd1 vccd1 _7774_/B sky130_fd_sc_hd__or4_2
X_7690_ _8562_/Q _7698_/B vssd1 vssd1 vccd1 vccd1 _7690_/X sky130_fd_sc_hd__or2_1
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7534__20 _7534__20/A vssd1 vssd1 vccd1 vccd1 _8534_/CLK sky130_fd_sc_hd__inv_2
X_8311_ _8311_/CLK _8311_/D vssd1 vssd1 vccd1 vccd1 _8311_/Q sky130_fd_sc_hd__dfxtp_1
X_5523_ _8135_/Q _4427_/A _5531_/S vssd1 vssd1 vccd1 vccd1 _5524_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5454_ _5454_/A vssd1 vssd1 vccd1 vccd1 _8170_/D sky130_fd_sc_hd__clkbuf_1
X_6634__277 _6636__279/A vssd1 vssd1 vccd1 vccd1 _8037_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3321_ _6816_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3321_/X sky130_fd_sc_hd__clkbuf_16
X_8242_ _8242_/CLK _8242_/D vssd1 vssd1 vccd1 vccd1 _8242_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3252_ _6601_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3252_/X sky130_fd_sc_hd__clkbuf_16
X_4405_ _4131_/X _8368_/Q _4407_/S vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__mux2_1
X_8173_ _8173_/CLK _8173_/D vssd1 vssd1 vccd1 vccd1 _8173_/Q sky130_fd_sc_hd__dfxtp_1
X_5385_ _5385_/A vssd1 vssd1 vccd1 vccd1 _5385_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4336_ _4336_/A _4336_/B _4027_/B vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__or3b_4
X_4267_ _4267_/A vssd1 vssd1 vccd1 vccd1 _8459_/D sky130_fd_sc_hd__clkbuf_1
X_7055_ _7055_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _8270_/D sky130_fd_sc_hd__nor2_1
X_6006_ _6006_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__or2_1
X_4198_ _8482_/Q _4197_/X _4204_/S vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7957_ _8633_/CLK _7957_/D vssd1 vssd1 vccd1 vccd1 _7957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6908_ _7579_/A _7581_/A vssd1 vssd1 vccd1 vccd1 _7688_/A sky130_fd_sc_hd__and2b_2
XFILLER_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7888_ _8569_/CLK _7888_/D vssd1 vssd1 vccd1 vccd1 _7888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6839_ _8552_/Q _8551_/Q vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__and2_1
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8509_ _8509_/CLK _8509_/D vssd1 vssd1 vccd1 vccd1 _8509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7477__149 _7477__149/A vssd1 vssd1 vccd1 vccd1 _8488_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5170_ _8293_/Q _8277_/Q _8539_/Q _8309_/Q _5341_/S _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5170_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4121_ _4121_/A vssd1 vssd1 vccd1 vccd1 _8497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _3962_/X _8522_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__mux2_1
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7811_ _7811_/A _7811_/B vssd1 vssd1 vccd1 vccd1 _7811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4954_ _4855_/X _7984_/Q _4817_/A _8217_/Q _4724_/A vssd1 vssd1 vccd1 vccd1 _4954_/X
+ sky130_fd_sc_hd__o221a_1
X_3905_ _3905_/A _3905_/B _3905_/C _3905_/D vssd1 vssd1 vccd1 vccd1 _3906_/C sky130_fd_sc_hd__or4_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _7906_/Q _4865_/X _4883_/X _4884_/X vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__o211a_1
X_7673_ _7672_/Y _7664_/B _7682_/A _7682_/B vssd1 vssd1 vccd1 vccd1 _7673_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6555_ _7760_/A vssd1 vssd1 vccd1 vccd1 _7836_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5506_ _5506_/A vssd1 vssd1 vccd1 vccd1 _8143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8225_ _8225_/CLK _8225_/D vssd1 vssd1 vccd1 vccd1 _8225_/Q sky130_fd_sc_hd__dfxtp_1
X_6486_ _7952_/Q _6483_/X _6474_/X _6485_/X _6472_/X vssd1 vssd1 vccd1 vccd1 _7952_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5437_ _5408_/X _8177_/Q _5441_/S vssd1 vssd1 vccd1 vccd1 _5438_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8156_ _8156_/CLK _8156_/D vssd1 vssd1 vccd1 vccd1 _8156_/Q sky130_fd_sc_hd__dfxtp_1
X_5368_ _3977_/X _5078_/A _5367_/X _5303_/X vssd1 vssd1 vccd1 vccd1 _8207_/D sky130_fd_sc_hd__o211a_1
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4319_ _4334_/S vssd1 vssd1 vccd1 vccd1 _4328_/S sky130_fd_sc_hd__buf_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5299_ _5294_/X _5295_/X _5171_/X _5298_/X vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__a211o_1
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8087_ _8630_/CLK _8087_/D vssd1 vssd1 vccd1 vccd1 _8087_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7038_ _7072_/A vssd1 vssd1 vccd1 vccd1 _7038_/X sky130_fd_sc_hd__buf_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7483__153 _7483__153/A vssd1 vssd1 vccd1 vccd1 _8492_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4670_ _8270_/Q vssd1 vssd1 vccd1 vccd1 _4672_/A sky130_fd_sc_hd__clkinv_2
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6271_ _8096_/Q _6269_/X _6270_/X _6263_/X _7885_/Q vssd1 vssd1 vccd1 vccd1 _7885_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_102_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _8197_/Q _5222_/B vssd1 vssd1 vccd1 vccd1 _5237_/A sky130_fd_sc_hd__or2_1
X_8010_ _8010_/CLK _8010_/D vssd1 vssd1 vccd1 vccd1 _8010_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3020_ _6218_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3020_/X sky130_fd_sc_hd__clkbuf_16
X_5153_ _3952_/X _5078_/X _5149_/X _5152_/X vssd1 vssd1 vccd1 vccd1 _8214_/D sky130_fd_sc_hd__o211a_1
X_4104_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__buf_2
XFILLER_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5084_ _5112_/A _5112_/B vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__and2_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4035_ _4035_/A vssd1 vssd1 vccd1 vccd1 _8530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5986_ _5986_/A vssd1 vssd1 vccd1 vccd1 _5986_/X sky130_fd_sc_hd__clkbuf_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4937_ _7904_/Q _4856_/X _4845_/A _4936_/X vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4868_ _8175_/Q _4865_/X _4796_/A _4867_/X vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__o211a_1
X_7656_ _7655_/X _7662_/B vssd1 vssd1 vccd1 vccd1 _7657_/A sky130_fd_sc_hd__and2b_1
X_6607_ _6625_/A vssd1 vssd1 vccd1 vccd1 _6607_/X sky130_fd_sc_hd__buf_1
X_4799_ _8331_/Q _8116_/Q _8068_/Q _8020_/Q _4731_/X _4729_/X vssd1 vssd1 vccd1 vccd1
+ _4799_/X sky130_fd_sc_hd__mux4_1
X_7587_ _7588_/B _7588_/C _7588_/A vssd1 vssd1 vccd1 vccd1 _7587_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6538_ _6538_/A vssd1 vssd1 vccd1 vccd1 _7973_/D sky130_fd_sc_hd__clkbuf_1
X_8682__247 vssd1 vssd1 vccd1 vccd1 _8682__247/HI versionID[1] sky130_fd_sc_hd__conb_1
XFILLER_97_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6469_ _7548_/A _6471_/B _6469_/C vssd1 vssd1 vccd1 vccd1 _6469_/X sky130_fd_sc_hd__and3_1
Xoutput160 _5946_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8208_ _8208_/CLK _8208_/D vssd1 vssd1 vccd1 vccd1 _8208_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput171 _5931_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__buf_2
X_8139_ _8139_/CLK _8139_/D vssd1 vssd1 vccd1 vccd1 _8139_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput193 _6171_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput182 _6135_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_48_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7016__432 _7017__433/A vssd1 vssd1 vccd1 vccd1 _8238_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _7921_/Q _4447_/A _5842_/S vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5771_ _5771_/A vssd1 vssd1 vccd1 vccd1 _8000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8490_ _8490_/CLK _8490_/D vssd1 vssd1 vccd1 vccd1 _8490_/Q sky130_fd_sc_hd__dfxtp_1
X_4722_ _7911_/Q _8031_/Q _8047_/Q _8015_/Q _4721_/X _4694_/A vssd1 vssd1 vccd1 vccd1
+ _4723_/B sky130_fd_sc_hd__mux4_1
X_7510_ _7541_/A vssd1 vssd1 vccd1 vccd1 _7510_/X sky130_fd_sc_hd__buf_1
X_4653_ _4653_/A vssd1 vssd1 vccd1 vccd1 _8276_/D sky130_fd_sc_hd__clkbuf_1
Xinput40 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__buf_4
X_6336__206 _6338__208/A vssd1 vssd1 vccd1 vccd1 _7918_/CLK sky130_fd_sc_hd__inv_2
X_4584_ _4584_/A vssd1 vssd1 vccd1 vccd1 _8306_/D sky130_fd_sc_hd__clkbuf_1
Xinput51 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _3905_/B sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _6017_/A sky130_fd_sc_hd__buf_4
Xinput73 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__buf_4
X_7372_ _7387_/A vssd1 vssd1 vccd1 vccd1 _7386_/A sky130_fd_sc_hd__clkbuf_2
Xinput95 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _7714_/A sky130_fd_sc_hd__buf_6
Xinput84 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6254_ _6249_/X _8086_/Q _6253_/X _6247_/X _7875_/Q vssd1 vssd1 vccd1 vccd1 _7875_/D
+ sky130_fd_sc_hd__o32a_1
X_5205_ _8505_/Q _8403_/Q _8140_/Q _8355_/Q _5169_/A _5140_/X vssd1 vssd1 vccd1 vccd1
+ _5205_/X sky130_fd_sc_hd__mux4_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6185_ _7890_/Q _6175_/X _6176_/X _6184_/X _6173_/X vssd1 vssd1 vccd1 vccd1 _6185_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5136_ _8294_/Q _8278_/Q _8540_/Q _8310_/Q _5130_/X _5101_/A vssd1 vssd1 vccd1 vccd1
+ _5136_/X sky130_fd_sc_hd__mux4_2
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3320_ clkbuf_0__3320_/X vssd1 vssd1 vccd1 vccd1 _6815__360/A sky130_fd_sc_hd__clkbuf_4
X_7434__114 _7435__115/A vssd1 vssd1 vccd1 vccd1 _8453_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5067_ _5067_/A vssd1 vssd1 vccd1 vccd1 _8220_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3251_ clkbuf_0__3251_/X vssd1 vssd1 vccd1 vccd1 _6619_/A sky130_fd_sc_hd__clkbuf_4
X_4018_ _4018_/A vssd1 vssd1 vccd1 vccd1 _8536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5969_ _7803_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__or2_1
XFILLER_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7708_ _7842_/A _7716_/B _7714_/C vssd1 vssd1 vccd1 vccd1 _7709_/A sky130_fd_sc_hd__and3_1
XFILLER_32_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7639_ _7638_/X _7649_/B vssd1 vssd1 vccd1 vccd1 _7640_/A sky130_fd_sc_hd__and2b_1
XFILLER_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3449_ clkbuf_0__3449_/X vssd1 vssd1 vccd1 vccd1 _7097_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6589__241 _6591__243/A vssd1 vssd1 vccd1 vccd1 _8001_/CLK sky130_fd_sc_hd__inv_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7990_ _7990_/CLK _7990_/D vssd1 vssd1 vccd1 vccd1 _7990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6941_ _6964_/A vssd1 vssd1 vccd1 vccd1 _6941_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3653_ clkbuf_0__3653_/X vssd1 vssd1 vccd1 vccd1 _7491__160/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6872_ _6872_/A _7611_/A _7611_/B vssd1 vssd1 vccd1 vccd1 _6872_/X sky130_fd_sc_hd__and3_1
Xclkbuf_1_1_0__3584_ clkbuf_0__3584_/X vssd1 vssd1 vccd1 vccd1 _7347__113/A sky130_fd_sc_hd__clkbuf_4
X_5823_ _5823_/A vssd1 vssd1 vccd1 vccd1 _7929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8611_ _8612_/CLK _8611_/D vssd1 vssd1 vccd1 vccd1 _8611_/Q sky130_fd_sc_hd__dfxtp_1
X_8542_ _8553_/CLK _8542_/D vssd1 vssd1 vccd1 vccd1 _8542_/Q sky130_fd_sc_hd__dfxtp_1
X_5754_ _5772_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5770_/S sky130_fd_sc_hd__nor2_2
X_8473_ _8473_/CLK _8473_/D vssd1 vssd1 vccd1 vccd1 _8473_/Q sky130_fd_sc_hd__dfxtp_1
X_5685_ _5685_/A vssd1 vssd1 vccd1 vccd1 _8039_/D sky130_fd_sc_hd__clkbuf_1
X_4705_ _4716_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4841_/A sky130_fd_sc_hd__xnor2_4
X_4636_ _4466_/X _8283_/Q _4638_/S vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__mux2_1
X_7424_ _8448_/Q _7424_/B vssd1 vssd1 vccd1 vccd1 _7424_/X sky130_fd_sc_hd__or2_1
X_7355_ _7387_/A vssd1 vssd1 vccd1 vccd1 _7371_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4567_ _8313_/Q _4525_/X _4571_/S vssd1 vssd1 vccd1 vccd1 _4568_/A sky130_fd_sc_hd__mux2_1
X_6306_ _6306_/A _6306_/B _6306_/C vssd1 vssd1 vccd1 vccd1 _6306_/X sky130_fd_sc_hd__and3_1
XFILLER_1_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4498_ _8572_/Q vssd1 vssd1 vccd1 vccd1 _4498_/X sky130_fd_sc_hd__clkbuf_4
X_7286_ _7834_/A _7286_/B vssd1 vssd1 vccd1 vccd1 _7330_/C sky130_fd_sc_hd__xor2_1
Xclkbuf_1_1_0__3018_ clkbuf_0__3018_/X vssd1 vssd1 vccd1 vccd1 _6209__183/A sky130_fd_sc_hd__clkbuf_4
X_6237_ _6232_/X _7897_/Q _6236_/X _6229_/X _7865_/Q vssd1 vssd1 vccd1 vccd1 _7865_/D
+ sky130_fd_sc_hd__o32a_1
X_6168_ _6168_/A _6172_/B vssd1 vssd1 vccd1 vccd1 _6168_/X sky130_fd_sc_hd__and2_4
XFILLER_97_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5119_ _8492_/Q _8476_/Q _8468_/Q _8500_/Q _5313_/S _5110_/X vssd1 vssd1 vccd1 vccd1
+ _5119_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _7941_/Q input30/X _6106_/S vssd1 vssd1 vccd1 vccd1 _6099_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5470_ _5470_/A vssd1 vssd1 vccd1 vccd1 _8162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4421_ _4127_/X _8361_/Q _4425_/S vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4352_ _4352_/A vssd1 vssd1 vccd1 vccd1 _8392_/D sky130_fd_sc_hd__clkbuf_1
X_4283_ _8424_/Q _4156_/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__mux2_1
X_6022_ _6022_/A vssd1 vssd1 vccd1 vccd1 _6022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7973_ _8608_/CLK _7973_/D vssd1 vssd1 vccd1 vccd1 _7973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6855_ _7564_/A _7626_/A _7626_/B vssd1 vssd1 vccd1 vccd1 _7584_/B sky130_fd_sc_hd__nand3_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5806_ _7984_/Q _5616_/A _5806_/S vssd1 vssd1 vccd1 vccd1 _5807_/A sky130_fd_sc_hd__mux2_1
X_3998_ _3974_/X _8579_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3999_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8525_ _8525_/CLK _8525_/D vssd1 vssd1 vccd1 vccd1 _8525_/Q sky130_fd_sc_hd__dfxtp_1
X_5737_ _5752_/S vssd1 vssd1 vccd1 vccd1 _5746_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8456_ _8456_/CLK _8456_/D vssd1 vssd1 vccd1 vccd1 _8456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _5598_/X _8046_/Q _5674_/S vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__mux2_1
X_7407_ _8443_/Q _7318_/A _7407_/C _7407_/D vssd1 vssd1 vccd1 vccd1 _7408_/C sky130_fd_sc_hd__and4bb_1
X_5599_ _5598_/X _8078_/Q _5608_/S vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3466_ _7159_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3466_/X sky130_fd_sc_hd__clkbuf_16
X_8387_ _8387_/CLK _8387_/D vssd1 vssd1 vccd1 vccd1 _8387_/Q sky130_fd_sc_hd__dfxtp_1
X_4619_ _8290_/Q _4495_/X _4619_/S vssd1 vssd1 vccd1 vccd1 _4620_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7338_ _7436_/A vssd1 vssd1 vccd1 vccd1 _7338_/X sky130_fd_sc_hd__buf_1
X_7269_ _8627_/Q vssd1 vssd1 vccd1 vccd1 _7569_/A sky130_fd_sc_hd__inv_2
XFILLER_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_20 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_31 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_42 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_64 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_86 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_75 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_53 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6210__184 _6211__185/A vssd1 vssd1 vccd1 vccd1 _7853_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6772__330 _6772__330/A vssd1 vssd1 vccd1 vccd1 _8122_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3079_ clkbuf_0__3079_/X vssd1 vssd1 vccd1 vccd1 _6340__210/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8452_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6820__364 _6821__365/A vssd1 vssd1 vccd1 vccd1 _8159_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _4979_/A _4970_/B _4970_/C vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__or3_4
XFILLER_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3921_ _7970_/Q _7971_/Q _7972_/Q _7969_/Q vssd1 vssd1 vccd1 vccd1 _6366_/D sky130_fd_sc_hd__or4b_2
X_5522_ _5537_/S vssd1 vssd1 vccd1 vccd1 _5531_/S sky130_fd_sc_hd__buf_2
X_8310_ _8310_/CLK _8310_/D vssd1 vssd1 vccd1 vccd1 _8310_/Q sky130_fd_sc_hd__dfxtp_1
X_5453_ _5404_/X _8170_/Q _5459_/S vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3320_ _6810_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3320_/X sky130_fd_sc_hd__clkbuf_16
X_8241_ _8241_/CLK _8241_/D vssd1 vssd1 vccd1 vccd1 _8241_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3251_ _6600_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3251_/X sky130_fd_sc_hd__clkbuf_16
X_4404_ _4404_/A vssd1 vssd1 vccd1 vccd1 _8369_/D sky130_fd_sc_hd__clkbuf_1
X_8172_ _8172_/CLK _8172_/D vssd1 vssd1 vccd1 vccd1 _8172_/Q sky130_fd_sc_hd__dfxtp_1
X_5384_ _5384_/A vssd1 vssd1 vccd1 vccd1 _8201_/D sky130_fd_sc_hd__clkbuf_1
X_4335_ _4335_/A vssd1 vssd1 vccd1 vccd1 _8399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7003__423 _7005__425/A vssd1 vssd1 vccd1 vccd1 _8229_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4266_ _8459_/Q _4194_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7054_ _7054_/A vssd1 vssd1 vccd1 vccd1 _8269_/D sky130_fd_sc_hd__clkbuf_1
X_6005_ _6005_/A vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__clkbuf_1
X_4197_ _8193_/Q vssd1 vssd1 vccd1 vccd1 _4197_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7207__83 _7208__84/A vssd1 vssd1 vccd1 vccd1 _8392_/CLK sky130_fd_sc_hd__inv_2
X_7956_ _8617_/CLK _7956_/D vssd1 vssd1 vccd1 vccd1 _7956_/Q sky130_fd_sc_hd__dfxtp_1
X_6907_ _8542_/Q vssd1 vssd1 vccd1 vccd1 _7581_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7887_ _8556_/CLK _7887_/D vssd1 vssd1 vccd1 vccd1 _7887_/Q sky130_fd_sc_hd__dfxtp_1
X_6838_ _8554_/Q vssd1 vssd1 vccd1 vccd1 _6838_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8508_ _8508_/CLK _8508_/D vssd1 vssd1 vccd1 vccd1 _8508_/Q sky130_fd_sc_hd__dfxtp_1
X_7010__427 _7013__430/A vssd1 vssd1 vccd1 vccd1 _8233_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8439_ _8439_/CLK _8439_/D vssd1 vssd1 vccd1 vccd1 _8439_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3449_ _7072_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3449_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6930__381 _6932__383/A vssd1 vssd1 vccd1 vccd1 _8177_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4120_ _4119_/X _8497_/Q _4124_/S vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _4051_/A vssd1 vssd1 vccd1 vccd1 _8523_/D sky130_fd_sc_hd__clkbuf_1
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7810_ _7808_/Y _7809_/Y _7800_/X vssd1 vssd1 vccd1 vccd1 _8622_/D sky130_fd_sc_hd__a21oi_1
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6640__282 _6641__283/A vssd1 vssd1 vccd1 vccd1 _8042_/CLK sky130_fd_sc_hd__inv_2
X_4953_ _4849_/X _8104_/Q _8000_/Q _4822_/A _4845_/A vssd1 vssd1 vccd1 vccd1 _4953_/X
+ sky130_fd_sc_hd__a221o_1
X_7741_ _7747_/A vssd1 vssd1 vccd1 vccd1 _7741_/X sky130_fd_sc_hd__buf_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3904_ _3904_/A _3904_/B input57/X input58/X vssd1 vssd1 vccd1 vccd1 _3906_/B sky130_fd_sc_hd__or4bb_1
X_7672_ _7672_/A vssd1 vssd1 vccd1 vccd1 _7672_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4884_ _4853_/A _8042_/Q _8026_/Q _4874_/A _4861_/A vssd1 vssd1 vccd1 vccd1 _4884_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148__536 _7149__537/A vssd1 vssd1 vccd1 vccd1 _8345_/CLK sky130_fd_sc_hd__inv_2
X_6554_ _6554_/A vssd1 vssd1 vccd1 vccd1 _7980_/D sky130_fd_sc_hd__clkbuf_1
X_5505_ _8143_/Q _4481_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5506_/A sky130_fd_sc_hd__mux2_1
X_6485_ _8617_/Q _6490_/B _6492_/C vssd1 vssd1 vccd1 vccd1 _6485_/X sky130_fd_sc_hd__and3_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5436_ _5436_/A vssd1 vssd1 vccd1 vccd1 _8178_/D sky130_fd_sc_hd__clkbuf_1
X_8224_ _8224_/CLK _8224_/D vssd1 vssd1 vccd1 vccd1 _8224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8155_ _8155_/CLK _8155_/D vssd1 vssd1 vccd1 vccd1 _8155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5367_ _8207_/Q _5081_/A _5386_/A _5366_/X _5148_/A vssd1 vssd1 vccd1 vccd1 _5367_/X
+ sky130_fd_sc_hd__a221o_1
X_4318_ _5539_/B _5503_/B vssd1 vssd1 vccd1 vccd1 _4334_/S sky130_fd_sc_hd__nor2_2
X_5298_ _5294_/A _5296_/X _5297_/X _5165_/A vssd1 vssd1 vccd1 vccd1 _5298_/X sky130_fd_sc_hd__o211a_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8086_ _8630_/CLK _8086_/D vssd1 vssd1 vccd1 vccd1 _8086_/Q sky130_fd_sc_hd__dfxtp_1
X_4249_ _8465_/Q _4226_/X _4251_/S vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _8610_/CLK _7939_/D vssd1 vssd1 vccd1 vccd1 _7939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6583__236 _6585__238/A vssd1 vssd1 vccd1 vccd1 _7996_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7201__78 _7203__80/A vssd1 vssd1 vccd1 vccd1 _8387_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6270_ _6306_/A vssd1 vssd1 vccd1 vccd1 _6270_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _5221_/A _5222_/B vssd1 vssd1 vccd1 vccd1 _5223_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _5377_/A vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4103_ _8577_/Q vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _8198_/Q _8197_/Q _8196_/Q vssd1 vssd1 vccd1 vccd1 _5112_/B sky130_fd_sc_hd__and3_1
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4034_ _3962_/X _8530_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4035_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5985_ _5985_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5986_/A sky130_fd_sc_hd__or2_4
X_7724_ _7724_/A vssd1 vssd1 vccd1 vccd1 _8577_/D sky130_fd_sc_hd__clkbuf_1
X_6937__387 _6937__387/A vssd1 vssd1 vccd1 vccd1 _8183_/CLK sky130_fd_sc_hd__inv_2
X_4936_ _4847_/A _8040_/Q _8024_/Q _4874_/A vssd1 vssd1 vccd1 vccd1 _4936_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4867_ _8236_/Q _4821_/X _4866_/X _4845_/A vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__o22a_1
X_7655_ _7654_/Y _7642_/X _7647_/X _7549_/B vssd1 vssd1 vccd1 vccd1 _7655_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7586_ _7586_/A _7586_/B _7586_/C _7586_/D vssd1 vssd1 vccd1 vccd1 _7593_/C sky130_fd_sc_hd__and4_1
XFILLER_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4798_ _4756_/S _4797_/X _4727_/X vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537_ _8088_/Q _7973_/Q _6537_/S vssd1 vssd1 vccd1 vccd1 _6538_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3249_ clkbuf_0__3249_/X vssd1 vssd1 vccd1 vccd1 _6593__245/A sky130_fd_sc_hd__clkbuf_4
X_6468_ _8621_/Q vssd1 vssd1 vccd1 vccd1 _7548_/A sky130_fd_sc_hd__clkbuf_4
Xoutput161 _6007_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__buf_2
Xoutput150 _5986_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5419_ _8190_/Q vssd1 vssd1 vccd1 vccd1 _5610_/A sky130_fd_sc_hd__clkbuf_2
X_6399_ _6394_/Y _6385_/X _6397_/Y _6398_/X _6387_/X vssd1 vssd1 vccd1 vccd1 _6400_/C
+ sky130_fd_sc_hd__o221a_1
X_8207_ _8207_/CLK _8207_/D vssd1 vssd1 vccd1 vccd1 _8207_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput172 _5935_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__buf_2
X_8138_ _8138_/CLK _8138_/D vssd1 vssd1 vccd1 vccd1 _8138_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput194 _6174_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput183 _6140_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8069_ _8069_/CLK _8069_/D vssd1 vssd1 vccd1 vccd1 _8069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3079_ _6335_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3079_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3465_ clkbuf_0__3465_/X vssd1 vssd1 vccd1 vccd1 _7157__544/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7734__35 _7734__35/A vssd1 vssd1 vccd1 vccd1 _8586_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5770_ _8000_/Q _5642_/X _5770_/S vssd1 vssd1 vccd1 vccd1 _5771_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4721_ _4806_/B vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__buf_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4652_ _8276_/Q _4489_/X _4656_/S vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__mux2_1
X_7186__66 _7188__68/A vssd1 vssd1 vccd1 vccd1 _8375_/CLK sky130_fd_sc_hd__inv_2
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4583_ _4441_/X _8306_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4584_/A sky130_fd_sc_hd__mux2_1
Xinput52 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _3905_/A sky130_fd_sc_hd__clkbuf_1
Xinput41 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _6039_/A sky130_fd_sc_hd__buf_4
Xinput63 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _6019_/A sky130_fd_sc_hd__buf_4
X_7371_ _7371_/A _7371_/B vssd1 vssd1 vccd1 vccd1 _8430_/D sky130_fd_sc_hd__nor2_1
X_6322_ _6322_/A vssd1 vssd1 vccd1 vccd1 _6322_/X sky130_fd_sc_hd__buf_1
Xinput96 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _7716_/A sky130_fd_sc_hd__clkbuf_8
Xinput85 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _5991_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _7803_/A sky130_fd_sc_hd__buf_4
X_6253_ _6306_/A vssd1 vssd1 vccd1 vccd1 _6253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5204_ _5204_/A vssd1 vssd1 vccd1 vccd1 _5351_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6184_ _6184_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__and2_1
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5135_ _5135_/A vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5066_ _4469_/X _8220_/Q _5066_/S vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3250_ clkbuf_0__3250_/X vssd1 vssd1 vccd1 vccd1 _6599__250/A sky130_fd_sc_hd__clkbuf_4
X_4017_ _8536_/Q _3940_/X _4017_/S vssd1 vssd1 vccd1 vccd1 _4018_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _5968_/A vssd1 vssd1 vccd1 vccd1 _5968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919_ _8478_/Q _4680_/A _4856_/X _8454_/Q _4687_/A vssd1 vssd1 vccd1 vccd1 _4919_/X
+ sky130_fd_sc_hd__o221a_1
X_7707_ _7842_/B vssd1 vssd1 vccd1 vccd1 _7716_/B sky130_fd_sc_hd__clkbuf_1
X_5899_ _5914_/S vssd1 vssd1 vccd1 vccd1 _5908_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7638_ _6891_/A _7620_/X _7625_/X _7551_/Y vssd1 vssd1 vccd1 vccd1 _7638_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7569_ _7569_/A _7626_/A _7626_/B vssd1 vssd1 vccd1 vccd1 _7569_/Y sky130_fd_sc_hd__nand3_1
XFILLER_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3448_ clkbuf_0__3448_/X vssd1 vssd1 vccd1 vccd1 _7069__473/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7105__501 _7105__501/A vssd1 vssd1 vccd1 vccd1 _8310_/CLK sky130_fd_sc_hd__inv_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7496__164 _7496__164/A vssd1 vssd1 vccd1 vccd1 _8503_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3652_ clkbuf_0__3652_/X vssd1 vssd1 vccd1 vccd1 _7483__153/A sky130_fd_sc_hd__clkbuf_4
X_6871_ _7607_/A _6876_/A _7610_/A vssd1 vssd1 vccd1 vccd1 _7611_/B sky130_fd_sc_hd__a21o_2
X_6342__211 _6343__212/A vssd1 vssd1 vccd1 vccd1 _7923_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3583_ clkbuf_0__3583_/X vssd1 vssd1 vccd1 vccd1 _7343__110/A sky130_fd_sc_hd__clkbuf_4
X_5822_ _5613_/X _7929_/Q _5824_/S vssd1 vssd1 vccd1 vccd1 _5823_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8610_ _8610_/CLK _8610_/D vssd1 vssd1 vccd1 vccd1 _8610_/Q sky130_fd_sc_hd__dfxtp_1
X_5753_ _5753_/A vssd1 vssd1 vccd1 vccd1 _8008_/D sky130_fd_sc_hd__clkbuf_1
X_8541_ _8553_/CLK _8541_/D vssd1 vssd1 vccd1 vccd1 _8541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4704_ _4704_/A vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__buf_2
X_8472_ _8472_/CLK _8472_/D vssd1 vssd1 vccd1 vccd1 _8472_/Q sky130_fd_sc_hd__dfxtp_1
X_5684_ _8039_/Q _5619_/X _5692_/S vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4635_ _4635_/A vssd1 vssd1 vccd1 vccd1 _8284_/D sky130_fd_sc_hd__clkbuf_1
X_7423_ _8210_/Q _7756_/B _7413_/X _7422_/X _7420_/X vssd1 vssd1 vccd1 vccd1 _8447_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _8314_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8623_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7354_ _7294_/B _7350_/Y _7353_/Y _7336_/X vssd1 vssd1 vccd1 vccd1 _8425_/D sky130_fd_sc_hd__o211a_1
XFILLER_116_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6305_ _6305_/A vssd1 vssd1 vccd1 vccd1 _7901_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3017_ clkbuf_0__3017_/X vssd1 vssd1 vccd1 vccd1 _6205__180/A sky130_fd_sc_hd__clkbuf_4
X_4497_ _4497_/A vssd1 vssd1 vccd1 vccd1 _8338_/D sky130_fd_sc_hd__clkbuf_1
X_7285_ _8428_/Q _7361_/A vssd1 vssd1 vccd1 vccd1 _7286_/B sky130_fd_sc_hd__xor2_2
X_6236_ _6236_/A vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _7883_/Q _6159_/X _6163_/X _6166_/X _6157_/X vssd1 vssd1 vccd1 vccd1 _6167_/X
+ sky130_fd_sc_hd__o221a_1
X_5118_ _5361_/S vssd1 vssd1 vccd1 vccd1 _5313_/S sky130_fd_sc_hd__clkbuf_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6098_ _6136_/A vssd1 vssd1 vccd1 vccd1 _6098_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _8227_/Q _4525_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _5050_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4420_ _4420_/A vssd1 vssd1 vccd1 vccd1 _8362_/D sky130_fd_sc_hd__clkbuf_1
X_7029__443 _7031__445/A vssd1 vssd1 vccd1 vccd1 _8250_/CLK sky130_fd_sc_hd__inv_2
X_4351_ _4131_/X _8392_/Q _4353_/S vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4282_ _4297_/S vssd1 vssd1 vccd1 vccd1 _4291_/S sky130_fd_sc_hd__buf_4
XFILLER_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6021_ _6021_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6022_/A sky130_fd_sc_hd__and2_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7972_ _7972_/CLK _7972_/D vssd1 vssd1 vccd1 vccd1 _7972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6923_ _6935_/A vssd1 vssd1 vccd1 vccd1 _6923_/X sky130_fd_sc_hd__buf_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6604__253 _6606__255/A vssd1 vssd1 vccd1 vccd1 _8013_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6854_ _7626_/A _7626_/B _7564_/A vssd1 vssd1 vccd1 vccd1 _7584_/A sky130_fd_sc_hd__a21o_1
X_6785_ _6785_/A vssd1 vssd1 vccd1 vccd1 _6785_/X sky130_fd_sc_hd__buf_1
X_3997_ _3997_/A vssd1 vssd1 vccd1 vccd1 _8580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5805_ _5805_/A vssd1 vssd1 vccd1 vccd1 _7985_/D sky130_fd_sc_hd__clkbuf_1
X_5736_ _5790_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5752_/S sky130_fd_sc_hd__nor2_2
X_8524_ _8524_/CLK _8524_/D vssd1 vssd1 vccd1 vccd1 _8524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5667_ _5667_/A vssd1 vssd1 vccd1 vccd1 _8047_/D sky130_fd_sc_hd__clkbuf_1
X_8455_ _8455_/CLK _8455_/D vssd1 vssd1 vccd1 vccd1 _8455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4618_ _4618_/A vssd1 vssd1 vccd1 vccd1 _8291_/D sky130_fd_sc_hd__clkbuf_1
X_7406_ _8442_/Q _7401_/X _7405_/Y _7336_/X vssd1 vssd1 vccd1 vccd1 _8442_/D sky130_fd_sc_hd__o211a_1
X_5598_ _5598_/A vssd1 vssd1 vccd1 vccd1 _5598_/X sky130_fd_sc_hd__clkbuf_4
X_8386_ _8386_/CLK _8386_/D vssd1 vssd1 vccd1 vccd1 _8386_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3465_ _7153_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3465_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _8320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7337_ _7321_/Y _7319_/C _7335_/X _7336_/X vssd1 vssd1 vccd1 vccd1 _8416_/D sky130_fd_sc_hd__o211a_1
X_6685__303 _6685__303/A vssd1 vssd1 vccd1 vccd1 _8071_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7268_ _7589_/A _7268_/B vssd1 vssd1 vccd1 vccd1 _7297_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_10 _5101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_43 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6349__217 _6351__219/A vssd1 vssd1 vccd1 vccd1 _7929_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_32 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_76 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_54 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_65 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_87 _3968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8655__220 vssd1 vssd1 vccd1 vccd1 _8655__220/HI core0Index[7] sky130_fd_sc_hd__conb_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7447__125 _7447__125/A vssd1 vssd1 vccd1 vccd1 _8464_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3078_ clkbuf_0__3078_/X vssd1 vssd1 vccd1 vccd1 _6331__202/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7098__496 _7099__497/A vssd1 vssd1 vccd1 vccd1 _8305_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _7977_/Q _7978_/Q _7979_/Q _7980_/Q vssd1 vssd1 vccd1 vccd1 _6366_/C sky130_fd_sc_hd__or4_2
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6570_ _6576_/A vssd1 vssd1 vccd1 vccd1 _6570_/X sky130_fd_sc_hd__buf_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5521_ _5521_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5537_/S sky130_fd_sc_hd__nor2_2
X_8240_ _8240_/CLK _8240_/D vssd1 vssd1 vccd1 vccd1 _8240_/Q sky130_fd_sc_hd__dfxtp_1
X_6673__295 _6673__295/A vssd1 vssd1 vccd1 vccd1 _8063_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5452_ _5452_/A vssd1 vssd1 vccd1 vccd1 _8171_/D sky130_fd_sc_hd__clkbuf_1
X_8171_ _8171_/CLK _8171_/D vssd1 vssd1 vccd1 vccd1 _8171_/Q sky130_fd_sc_hd__dfxtp_1
X_4403_ _4127_/X _8369_/Q _4407_/S vssd1 vssd1 vccd1 vccd1 _4404_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3250_ _6594_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3250_/X sky130_fd_sc_hd__clkbuf_16
X_5383_ _5383_/A _6986_/B _5383_/C vssd1 vssd1 vccd1 vccd1 _5384_/A sky130_fd_sc_hd__and3_1
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4334_ _8399_/Q _4238_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__mux2_1
X_7122_ _7122_/A vssd1 vssd1 vccd1 vccd1 _7122_/X sky130_fd_sc_hd__buf_1
XFILLER_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7053_ _7053_/A _8163_/Q _7053_/C vssd1 vssd1 vccd1 vccd1 _7054_/A sky130_fd_sc_hd__and3_1
X_6004_ _6004_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _6005_/A sky130_fd_sc_hd__or2_1
X_4265_ _4265_/A vssd1 vssd1 vccd1 vccd1 _8460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4196_ _4196_/A vssd1 vssd1 vccd1 vccd1 _8483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7955_ _8091_/CLK _7955_/D vssd1 vssd1 vccd1 vccd1 _7955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6906_ _8541_/Q vssd1 vssd1 vccd1 vccd1 _7579_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7886_ _8569_/CLK _7886_/D vssd1 vssd1 vccd1 vccd1 _7886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6837_ _7798_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6847_/A sky130_fd_sc_hd__nand2_1
X_8507_ _8507_/CLK _8507_/D vssd1 vssd1 vccd1 vccd1 _8507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5719_ _5734_/S vssd1 vssd1 vccd1 vccd1 _5728_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_6_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6699_ _6699_/A vssd1 vssd1 vccd1 vccd1 _8080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7540__25 _7540__25/A vssd1 vssd1 vccd1 vccd1 _8539_/CLK sky130_fd_sc_hd__inv_2
X_8438_ _8631_/CLK _8438_/D vssd1 vssd1 vccd1 vccd1 _8438_/Q sky130_fd_sc_hd__dfxtp_1
X_8369_ _8369_/CLK _8369_/D vssd1 vssd1 vccd1 vccd1 _8369_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3448_ _7066_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3448_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _3959_/X _8523_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4952_ _4845_/X _4950_/X _4951_/X vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4883_ _8010_/Q _4716_/B _4821_/A vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__a21o_1
X_3903_ _3903_/A _3903_/B input69/X vssd1 vssd1 vccd1 vccd1 _3906_/A sky130_fd_sc_hd__or3b_1
X_7671_ _7682_/A _7682_/B vssd1 vssd1 vccd1 vccd1 _7671_/Y sky130_fd_sc_hd__nor2_1
X_6553_ _8095_/Q _7980_/Q _6804_/S vssd1 vssd1 vccd1 vccd1 _6554_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5504_ _5519_/S vssd1 vssd1 vccd1 vccd1 _5513_/S sky130_fd_sc_hd__clkbuf_2
X_6484_ _8146_/Q vssd1 vssd1 vccd1 vccd1 _6492_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5435_ _5404_/X _8178_/Q _5441_/S vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__mux2_1
X_8223_ _8223_/CLK _8223_/D vssd1 vssd1 vccd1 vccd1 _8223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8154_ _8154_/CLK _8154_/D vssd1 vssd1 vccd1 vccd1 _8154_/Q sky130_fd_sc_hd__dfxtp_1
X_5366_ _5387_/B _5344_/X _5351_/X _5365_/X vssd1 vssd1 vccd1 vccd1 _5366_/X sky130_fd_sc_hd__a31o_1
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4317_ _4317_/A vssd1 vssd1 vccd1 vccd1 _8407_/D sky130_fd_sc_hd__clkbuf_1
X_5297_ _8580_/Q _5276_/A _5238_/A _8596_/Q vssd1 vssd1 vccd1 vccd1 _5297_/X sky130_fd_sc_hd__o22a_1
X_8085_ _8625_/CLK _8085_/D vssd1 vssd1 vccd1 vccd1 _8085_/Q sky130_fd_sc_hd__dfxtp_1
X_4248_ _4248_/A vssd1 vssd1 vccd1 vccd1 _8466_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3481_ clkbuf_0__3481_/X vssd1 vssd1 vccd1 vccd1 _7231__102/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4179_ _8253_/Q _4666_/C _4179_/C _8258_/Q vssd1 vssd1 vccd1 vccd1 _4179_/X sky130_fd_sc_hd__and4bb_1
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7938_ _8570_/CLK _7938_/D vssd1 vssd1 vccd1 vccd1 _7938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7869_ _8631_/CLK _7869_/D vssd1 vssd1 vccd1 vccd1 _7869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7490__159 _7491__160/A vssd1 vssd1 vccd1 vccd1 _8498_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995__416 _6997__418/A vssd1 vssd1 vccd1 vccd1 _8222_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _6964_/A sky130_fd_sc_hd__clkbuf_16
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5220_ _5276_/A vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _6986_/B vssd1 vssd1 vccd1 vccd1 _5377_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4102_ _4102_/A vssd1 vssd1 vccd1 vccd1 _8501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5082_ _5216_/A vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4033_ _4033_/A vssd1 vssd1 vccd1 vccd1 _8531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7154__541 _7158__545/A vssd1 vssd1 vccd1 vccd1 _8350_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5984_ _5995_/A vssd1 vssd1 vccd1 vccd1 _5993_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7723_ _7723_/A _7723_/B _7723_/C vssd1 vssd1 vccd1 vccd1 _7724_/A sky130_fd_sc_hd__and3_1
X_4935_ _4815_/X _8032_/Q _7845_/Q _4865_/X _4756_/S vssd1 vssd1 vccd1 vccd1 _4935_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4866_ _4849_/A _8167_/Q _7995_/Q _4847_/A vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__a22o_1
X_7654_ _8555_/Q vssd1 vssd1 vccd1 vccd1 _7654_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4797_ _7849_/Q _7857_/Q _7932_/Q _8036_/Q _4721_/X _4694_/A vssd1 vssd1 vccd1 vccd1
+ _4797_/X sky130_fd_sc_hd__mux4_1
X_7585_ _8621_/Q _7549_/B _6869_/B _7821_/A vssd1 vssd1 vccd1 vccd1 _7586_/D sky130_fd_sc_hd__o22a_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6536_ _6536_/A vssd1 vssd1 vccd1 vccd1 _7972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3248_ clkbuf_0__3248_/X vssd1 vssd1 vccd1 vccd1 _6585__238/A sky130_fd_sc_hd__clkbuf_4
X_6467_ _7947_/Q _6464_/X _6452_/X _6466_/X _6459_/X vssd1 vssd1 vccd1 vccd1 _7947_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput151 _5988_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput140 _5966_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__buf_2
X_5418_ _5418_/A vssd1 vssd1 vccd1 vccd1 _8183_/D sky130_fd_sc_hd__clkbuf_1
X_6398_ _6436_/B vssd1 vssd1 vccd1 vccd1 _6398_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8206_ _8206_/CLK _8206_/D vssd1 vssd1 vccd1 vccd1 _8206_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput173 _5937_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__buf_2
Xoutput162 _6009_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__buf_2
X_8137_ _8137_/CLK _8137_/D vssd1 vssd1 vccd1 vccd1 _8137_/Q sky130_fd_sc_hd__dfxtp_1
X_5349_ _8351_/Q _5276_/X _5249_/A _8501_/Q _5120_/A vssd1 vssd1 vccd1 vccd1 _5349_/X
+ sky130_fd_sc_hd__o221a_1
Xoutput195 _6179_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput184 _6143_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__buf_2
X_8068_ _8068_/CLK _8068_/D vssd1 vssd1 vccd1 vccd1 _8068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3464_ clkbuf_0__3464_/X vssd1 vssd1 vccd1 vccd1 _7149__537/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3078_ _6329_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3078_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7023__438 _7023__438/A vssd1 vssd1 vccd1 vccd1 _8244_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8635__251 vssd1 vssd1 vccd1 vccd1 partID[0] _8635__251/LO sky130_fd_sc_hd__conb_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4720_ _4699_/X _4711_/X _4719_/X vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__a21o_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4651_ _4651_/A vssd1 vssd1 vccd1 vccd1 _8277_/D sky130_fd_sc_hd__clkbuf_1
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _6172_/A sky130_fd_sc_hd__clkbuf_1
X_4582_ _4582_/A vssd1 vssd1 vccd1 vccd1 _8307_/D sky130_fd_sc_hd__clkbuf_1
Xinput53 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _3905_/D sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _6021_/A sky130_fd_sc_hd__buf_4
Xinput42 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _6041_/A sky130_fd_sc_hd__buf_4
X_7370_ _7274_/A _7368_/X _7360_/X _7369_/Y vssd1 vssd1 vccd1 vccd1 _7371_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput97 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _7719_/A sky130_fd_sc_hd__buf_4
Xinput86 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput75 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _7799_/A sky130_fd_sc_hd__buf_4
XFILLER_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6252_ _6249_/X _8085_/Q _6245_/X _6247_/X _7874_/Q vssd1 vssd1 vccd1 vccd1 _7874_/D
+ sky130_fd_sc_hd__o32a_1
X_5203_ _5095_/A _5200_/X _5202_/X vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__a21o_1
X_6183_ _7889_/Q _6175_/X _6176_/X _6182_/X _6173_/X vssd1 vssd1 vccd1 vccd1 _6183_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _5134_/A vssd1 vssd1 vccd1 vccd1 _5135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5065_ _5065_/A vssd1 vssd1 vccd1 vccd1 _8221_/D sky130_fd_sc_hd__clkbuf_1
X_4016_ _4016_/A vssd1 vssd1 vccd1 vccd1 _8537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5967_ _5967_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5968_/A sky130_fd_sc_hd__or2_1
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _8344_/Q _4849_/X _4822_/X _8057_/Q vssd1 vssd1 vccd1 vccd1 _4918_/X sky130_fd_sc_hd__a22o_1
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7706_ _7794_/B vssd1 vssd1 vccd1 vccd1 _7842_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5898_ _5898_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5914_/S sky130_fd_sc_hd__or2_2
X_7637_ _7637_/A vssd1 vssd1 vccd1 vccd1 _8550_/D sky130_fd_sc_hd__clkbuf_1
X_4849_ _4849_/A vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__buf_2
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7568_ _7626_/A _7626_/B _7569_/A vssd1 vssd1 vccd1 vccd1 _7568_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6519_ _6519_/A vssd1 vssd1 vccd1 vccd1 _7964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3447_ clkbuf_0__3447_/X vssd1 vssd1 vccd1 vccd1 _7065__470/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3651_ clkbuf_0__3651_/X vssd1 vssd1 vccd1 vccd1 _7498_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6870_ _7610_/A _7607_/A _6876_/A vssd1 vssd1 vccd1 vccd1 _7611_/A sky130_fd_sc_hd__nand3_4
X_5821_ _5821_/A vssd1 vssd1 vccd1 vccd1 _7930_/D sky130_fd_sc_hd__clkbuf_1
X_8672__237 vssd1 vssd1 vccd1 vccd1 _8672__237/HI manufacturerID[9] sky130_fd_sc_hd__conb_1
XFILLER_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6596__247 _6596__247/A vssd1 vssd1 vccd1 vccd1 _8007_/CLK sky130_fd_sc_hd__inv_2
X_8540_ _8540_/CLK _8540_/D vssd1 vssd1 vccd1 vccd1 _8540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ _8008_/Q _5642_/X _5752_/S vssd1 vssd1 vccd1 vccd1 _5753_/A sky130_fd_sc_hd__mux2_1
X_4703_ _8224_/Q _8111_/Q _8007_/Q _7991_/Q _4700_/X _4702_/X vssd1 vssd1 vccd1 vccd1
+ _4703_/X sky130_fd_sc_hd__mux4_1
X_8471_ _8471_/CLK _8471_/D vssd1 vssd1 vccd1 vccd1 _8471_/Q sky130_fd_sc_hd__dfxtp_1
X_5683_ _5698_/S vssd1 vssd1 vccd1 vccd1 _5692_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_8_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3481_ _7229_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3481_/X sky130_fd_sc_hd__clkbuf_16
X_4634_ _4463_/X _8284_/Q _4638_/S vssd1 vssd1 vccd1 vccd1 _4635_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7422_ _8447_/Q _7424_/B vssd1 vssd1 vccd1 vccd1 _7422_/X sky130_fd_sc_hd__or2_1
XFILLER_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4565_ _8314_/Q _4522_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__mux2_1
X_7353_ _7294_/B _7358_/A _7352_/X vssd1 vssd1 vccd1 vccd1 _7353_/Y sky130_fd_sc_hd__o21bai_1
X_6304_ _6307_/B _6304_/B _6306_/C vssd1 vssd1 vccd1 vccd1 _6305_/A sky130_fd_sc_hd__and3_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3016_ clkbuf_0__3016_/X vssd1 vssd1 vccd1 vccd1 _6212_/A sky130_fd_sc_hd__clkbuf_4
X_4496_ _8338_/Q _4495_/X _4496_/S vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__mux2_1
X_7284_ _8427_/Q _8426_/Q _8425_/Q vssd1 vssd1 vccd1 vccd1 _7361_/A sky130_fd_sc_hd__nand3_2
XFILLER_103_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6235_ _6232_/X _7896_/Q _6225_/X _6229_/X _7864_/Q vssd1 vssd1 vccd1 vccd1 _7864_/D
+ sky130_fd_sc_hd__o32a_1
X_6166_ _6166_/A _6172_/B vssd1 vssd1 vccd1 vccd1 _6166_/X sky130_fd_sc_hd__and2_4
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5258_/S vssd1 vssd1 vccd1 vccd1 _5361_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_85_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6073_/X _6095_/X _6096_/X _6082_/X vssd1 vssd1 vccd1 vccd1 _6097_/X sky130_fd_sc_hd__o211a_1
X_5048_ _5048_/A vssd1 vssd1 vccd1 vccd1 _8228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7100__498 _7102__500/A vssd1 vssd1 vccd1 vccd1 _8307_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4350_ _4350_/A vssd1 vssd1 vccd1 vccd1 _8393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4281_ _5682_/A _5594_/A vssd1 vssd1 vccd1 vccd1 _4297_/S sky130_fd_sc_hd__nor2_2
X_6020_ _6020_/A vssd1 vssd1 vccd1 vccd1 _6020_/X sky130_fd_sc_hd__clkbuf_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7219__93 _7219__93/A vssd1 vssd1 vccd1 vccd1 _8402_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7971_ _7972_/CLK _7971_/D vssd1 vssd1 vccd1 vccd1 _7971_/Q sky130_fd_sc_hd__dfxtp_1
X_6922_ _6970_/A vssd1 vssd1 vccd1 vccd1 _6922_/X sky130_fd_sc_hd__buf_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6853_ _8547_/Q _6842_/C _8548_/Q vssd1 vssd1 vccd1 vccd1 _7626_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5804_ _7985_/Q _5613_/A _5806_/S vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__mux2_1
X_3996_ _3971_/X _8580_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3997_/A sky130_fd_sc_hd__mux2_1
X_5735_ _5735_/A vssd1 vssd1 vccd1 vccd1 _8016_/D sky130_fd_sc_hd__clkbuf_1
X_8523_ _8523_/CLK _8523_/D vssd1 vssd1 vccd1 vccd1 _8523_/Q sky130_fd_sc_hd__dfxtp_1
X_5666_ _5593_/X _8047_/Q _5674_/S vssd1 vssd1 vccd1 vccd1 _5667_/A sky130_fd_sc_hd__mux2_1
X_8454_ _8454_/CLK _8454_/D vssd1 vssd1 vccd1 vccd1 _8454_/Q sky130_fd_sc_hd__dfxtp_1
X_4617_ _8291_/Q _4492_/X _4619_/S vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__mux2_1
X_7405_ _7321_/Y _7318_/A _7407_/C _7408_/B vssd1 vssd1 vccd1 vccd1 _7405_/Y sky130_fd_sc_hd__o31ai_1
X_5597_ _5597_/A vssd1 vssd1 vccd1 vccd1 _8079_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3464_ _7147_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3464_/X sky130_fd_sc_hd__clkbuf_16
X_8385_ _8385_/CLK _8385_/D vssd1 vssd1 vccd1 vccd1 _8385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4548_ _4447_/X _8320_/Q _4550_/S vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7336_ _7420_/A vssd1 vssd1 vccd1 vccd1 _7336_/X sky130_fd_sc_hd__clkbuf_2
X_4479_ _4478_/X _8343_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__mux2_1
X_7267_ _8435_/Q _7267_/B vssd1 vssd1 vccd1 vccd1 _7268_/B sky130_fd_sc_hd__xnor2_2
X_6218_ _6322_/A vssd1 vssd1 vccd1 vccd1 _6218_/X sky130_fd_sc_hd__buf_1
X_7198_ _7210_/A vssd1 vssd1 vccd1 vccd1 _7198_/X sky130_fd_sc_hd__buf_1
XFILLER_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_11 _5162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6149_ _6149_/A vssd1 vssd1 vccd1 vccd1 _6175_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_22 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_33 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_77 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_66 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_44 _6188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_55 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_88 _5162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3077_ clkbuf_0__3077_/X vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6963__395 _6963__395/A vssd1 vssd1 vccd1 vccd1 _8199_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5520_/A vssd1 vssd1 vccd1 vccd1 _8136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5451_ _5398_/X _8171_/Q _5459_/S vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__mux2_1
X_8170_ _8170_/CLK _8170_/D vssd1 vssd1 vccd1 vccd1 _8170_/Q sky130_fd_sc_hd__dfxtp_1
X_4402_ _4402_/A vssd1 vssd1 vccd1 vccd1 _8370_/D sky130_fd_sc_hd__clkbuf_1
X_5382_ _5382_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5383_/C sky130_fd_sc_hd__or2_1
X_4333_ _4333_/A vssd1 vssd1 vccd1 vccd1 _8400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4264_ _8460_/Q _4156_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4265_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6003_ _6003_/A vssd1 vssd1 vccd1 vccd1 _6003_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4195_ _8483_/Q _4194_/X _4204_/S vssd1 vssd1 vccd1 vccd1 _4196_/A sky130_fd_sc_hd__mux2_1
X_8678__243 vssd1 vssd1 vccd1 vccd1 _8678__243/HI partID[9] sky130_fd_sc_hd__conb_1
X_7118__512 _7119__513/A vssd1 vssd1 vccd1 vccd1 _8321_/CLK sky130_fd_sc_hd__inv_2
X_7954_ _8091_/CLK _7954_/D vssd1 vssd1 vccd1 vccd1 _7954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _7793_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _7593_/A sky130_fd_sc_hd__xor2_1
X_7885_ _8556_/CLK _7885_/D vssd1 vssd1 vccd1 vccd1 _7885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6836_ _7588_/B _7588_/C vssd1 vssd1 vccd1 vccd1 _6846_/B sky130_fd_sc_hd__nand2_2
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6767_ _6791_/A vssd1 vssd1 vccd1 vccd1 _6767_/X sky130_fd_sc_hd__buf_1
X_8506_ _8506_/CLK _8506_/D vssd1 vssd1 vccd1 vccd1 _8506_/Q sky130_fd_sc_hd__dfxtp_1
X_5718_ _5790_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5734_/S sky130_fd_sc_hd__nor2_2
X_7525__12 _7526__13/A vssd1 vssd1 vccd1 vccd1 _8526_/CLK sky130_fd_sc_hd__inv_2
X_3979_ _3979_/A vssd1 vssd1 vccd1 vccd1 _8586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3479_ clkbuf_0__3479_/X vssd1 vssd1 vccd1 vccd1 _7224__97/A sky130_fd_sc_hd__clkbuf_4
X_6698_ _7818_/A _8080_/Q _6706_/S vssd1 vssd1 vccd1 vccd1 _6699_/A sky130_fd_sc_hd__mux2_1
X_5649_ _5598_/X _8062_/Q _5655_/S vssd1 vssd1 vccd1 vccd1 _5650_/A sky130_fd_sc_hd__mux2_1
X_6355__222 _6356__223/A vssd1 vssd1 vccd1 vccd1 _7934_/CLK sky130_fd_sc_hd__inv_2
X_8437_ _8439_/CLK _8437_/D vssd1 vssd1 vccd1 vccd1 _8437_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3447_ _7060_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3447_/X sky130_fd_sc_hd__clkbuf_16
X_8368_ _8368_/CLK _8368_/D vssd1 vssd1 vccd1 vccd1 _8368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7319_ _7420_/A _7319_/B _7319_/C vssd1 vssd1 vccd1 vccd1 _7320_/A sky130_fd_sc_hd__and3_1
X_8299_ _8299_/CLK _8299_/D vssd1 vssd1 vccd1 vccd1 _8299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7213__88 _7214__89/A vssd1 vssd1 vccd1 vccd1 _8397_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _8311_/Q _4855_/X _4817_/A _8295_/Q _4834_/X vssd1 vssd1 vccd1 vccd1 _4951_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3902_ _3902_/A _3902_/B _3902_/C _3902_/D vssd1 vssd1 vccd1 vccd1 _3907_/C sky130_fd_sc_hd__or4_2
X_7670_ _7688_/A _7681_/B _7688_/B vssd1 vssd1 vccd1 vccd1 _7682_/B sky130_fd_sc_hd__and3_1
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4882_ _4831_/X _8034_/Q _7847_/Q _4833_/X _4758_/A vssd1 vssd1 vccd1 vccd1 _4882_/X
+ sky130_fd_sc_hd__o221a_1
X_6552_ _6552_/A vssd1 vssd1 vccd1 vccd1 _7979_/D sky130_fd_sc_hd__clkbuf_1
X_5503_ _5521_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _5519_/S sky130_fd_sc_hd__nor2_2
X_6483_ _6483_/A vssd1 vssd1 vccd1 vccd1 _6483_/X sky130_fd_sc_hd__clkbuf_2
X_5434_ _5434_/A vssd1 vssd1 vccd1 vccd1 _8179_/D sky130_fd_sc_hd__clkbuf_1
X_8222_ _8222_/CLK _8222_/D vssd1 vssd1 vccd1 vccd1 _8222_/Q sky130_fd_sc_hd__dfxtp_1
X_8153_ _8153_/CLK _8153_/D vssd1 vssd1 vccd1 vccd1 _8153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7104_ _7122_/A vssd1 vssd1 vccd1 vccd1 _7104_/X sky130_fd_sc_hd__buf_1
X_5365_ _5389_/B _5354_/X _5357_/X _5364_/X _5087_/A vssd1 vssd1 vccd1 vccd1 _5365_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5296_ _8122_/Q _8149_/Q _5361_/S vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__mux2_1
X_4316_ _8407_/Q _4238_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__mux2_1
X_8084_ _8625_/CLK _8084_/D vssd1 vssd1 vccd1 vccd1 _8084_/Q sky130_fd_sc_hd__dfxtp_1
X_4247_ _8466_/Q _4223_/X _4251_/S vssd1 vssd1 vccd1 vccd1 _4248_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3480_ clkbuf_0__3480_/X vssd1 vssd1 vccd1 vccd1 _7442_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4178_ _8258_/Q _4175_/Y _4969_/B vssd1 vssd1 vccd1 vccd1 _4178_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7937_ _8452_/CLK _7937_/D vssd1 vssd1 vccd1 vccd1 _7937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7746__45 _7746__45/A vssd1 vssd1 vccd1 vccd1 _8596_/CLK sky130_fd_sc_hd__inv_2
X_7868_ _8631_/CLK _7868_/D vssd1 vssd1 vccd1 vccd1 _7868_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7799_ _7799_/A _7812_/B vssd1 vssd1 vccd1 vccd1 _7799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6617__264 _6618__265/A vssd1 vssd1 vccd1 vccd1 _8024_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5150_ _5150_/A vssd1 vssd1 vccd1 vccd1 _6986_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4101_ _8501_/Q _3949_/X _4101_/S vssd1 vssd1 vccd1 vccd1 _4102_/A sky130_fd_sc_hd__mux2_1
X_5081_ _5081_/A _7410_/A vssd1 vssd1 vccd1 vccd1 _5216_/A sky130_fd_sc_hd__nor2_1
XFILLER_111_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _3959_/X _8531_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4033_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5983_ _5983_/A vssd1 vssd1 vccd1 vccd1 _5983_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4934_ _4665_/X _7928_/Q _7853_/Q _4812_/X _4861_/X vssd1 vssd1 vccd1 vccd1 _4934_/X
+ sky130_fd_sc_hd__a221o_1
X_7722_ _7722_/A vssd1 vssd1 vccd1 vccd1 _8576_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_19_wb_clk_i _6197_/A vssd1 vssd1 vccd1 vccd1 _8622_/CLK sky130_fd_sc_hd__clkbuf_16
X_6792__346 _6794__348/A vssd1 vssd1 vccd1 vccd1 _8138_/CLK sky130_fd_sc_hd__inv_2
X_4865_ _4865_/A vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__buf_2
X_7653_ _7653_/A vssd1 vssd1 vccd1 vccd1 _8554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4796_ _4796_/A _4796_/B vssd1 vssd1 vccd1 vccd1 _4796_/X sky130_fd_sc_hd__and2_1
X_7584_ _7584_/A _7584_/B vssd1 vssd1 vccd1 vccd1 _7586_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0__3316_ clkbuf_0__3316_/X vssd1 vssd1 vccd1 vccd1 _6799__351/A sky130_fd_sc_hd__clkbuf_4
X_6535_ _8087_/Q _7972_/Q _6537_/S vssd1 vssd1 vccd1 vccd1 _6536_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3247_ clkbuf_0__3247_/X vssd1 vssd1 vccd1 vccd1 _6578__232/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6466_ _7808_/A _6471_/B _6469_/C vssd1 vssd1 vccd1 vccd1 _6466_/X sky130_fd_sc_hd__and3_1
X_8205_ _8205_/CLK _8205_/D vssd1 vssd1 vccd1 vccd1 _8205_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput152 _5990_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput130 _6018_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput141 _5968_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__buf_2
X_5417_ _5416_/X _8183_/Q _5417_/S vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__mux2_1
X_6397_ _8049_/Q _6395_/X _7055_/B vssd1 vssd1 vccd1 vccd1 _6397_/Y sky130_fd_sc_hd__a21oi_1
Xoutput174 _5925_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput163 _5948_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__buf_2
X_8136_ _8136_/CLK _8136_/D vssd1 vssd1 vccd1 vccd1 _8136_/Q sky130_fd_sc_hd__dfxtp_1
X_5348_ _8399_/Q _8136_/Q _5355_/S vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput185 _6146_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8067_ _8067_/CLK _8067_/D vssd1 vssd1 vccd1 vccd1 _8067_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput196 _6181_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__buf_2
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5279_ _5344_/A _5279_/B _5279_/C vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__or3_1
Xclkbuf_0__3077_ _6328_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3077_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3463_ clkbuf_0__3463_/X vssd1 vssd1 vccd1 vccd1 _7144__533/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7466__140 _7466__140/A vssd1 vssd1 vccd1 vccd1 _8479_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4650_ _8277_/Q _4486_/X _4656_/S vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__mux2_1
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__clkbuf_4
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_4
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4581_ _4438_/X _8307_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4582_/A sky130_fd_sc_hd__mux2_1
Xinput54 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _3905_/C sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _6077_/A sky130_fd_sc_hd__buf_2
Xinput76 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _7796_/A sky130_fd_sc_hd__buf_4
Xinput87 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__buf_4
Xinput65 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _6023_/A sky130_fd_sc_hd__buf_4
Xinput98 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _7828_/A sky130_fd_sc_hd__buf_4
XFILLER_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6251_ _6249_/X _8084_/Q _6245_/X _6247_/X _7873_/Q vssd1 vssd1 vccd1 vccd1 _7873_/D
+ sky130_fd_sc_hd__o32a_1
X_5202_ _5121_/X _5201_/X _5171_/X vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__a21o_1
X_6182_ _6182_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__and2_1
XFILLER_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5133_ _5209_/A _5133_/B vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__and2_1
XFILLER_111_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _4466_/X _8221_/Q _5066_/S vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__mux2_1
X_4015_ _8537_/Q _3937_/X _4017_/S vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5966_/A vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5897_ _5897_/A vssd1 vssd1 vccd1 vccd1 _7853_/D sky130_fd_sc_hd__clkbuf_1
X_4917_ _4869_/X _4907_/X _4910_/X _4916_/X _4990_/B vssd1 vssd1 vccd1 vccd1 _4917_/X
+ sky130_fd_sc_hd__o311a_1
X_7705_ _7575_/X _7687_/A _7704_/X _7684_/A vssd1 vssd1 vccd1 vccd1 _8569_/D sky130_fd_sc_hd__o211a_1
X_4848_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4849_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7636_ _7635_/X _7649_/B vssd1 vssd1 vccd1 vccd1 _7637_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4779_ _4756_/S _4778_/X _4727_/X vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__a21o_1
X_7567_ _7566_/B _7566_/C _8626_/Q vssd1 vssd1 vccd1 vccd1 _7567_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7498_ _7498_/A vssd1 vssd1 vccd1 vccd1 _7498_/X sky130_fd_sc_hd__buf_1
X_6518_ _6025_/A _7964_/Q _6526_/S vssd1 vssd1 vccd1 vccd1 _6519_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6449_ _6436_/Y _6446_/X _6448_/X vssd1 vssd1 vccd1 vccd1 _6449_/Y sky130_fd_sc_hd__a21oi_1
X_8119_ _8119_/CLK _8119_/D vssd1 vssd1 vccd1 vccd1 _8119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3650_ clkbuf_0__3650_/X vssd1 vssd1 vccd1 vccd1 _7478__150/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5610_/X _7930_/Q _5824_/S vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7112__507 _7114__509/A vssd1 vssd1 vccd1 vccd1 _8316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5751_ _5751_/A vssd1 vssd1 vccd1 vccd1 _8009_/D sky130_fd_sc_hd__clkbuf_1
X_4702_ _4702_/A vssd1 vssd1 vccd1 vccd1 _4702_/X sky130_fd_sc_hd__buf_2
X_8470_ _8470_/CLK _8470_/D vssd1 vssd1 vccd1 vccd1 _8470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5682_ _5682_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5698_/S sky130_fd_sc_hd__nor2_2
X_7421_ _8209_/Q _7756_/B _7413_/X _7419_/X _7420_/X vssd1 vssd1 vccd1 vccd1 _8446_/D
+ sky130_fd_sc_hd__o311a_1
Xclkbuf_0__3480_ _7228_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3480_/X sky130_fd_sc_hd__clkbuf_16
X_4633_ _4633_/A vssd1 vssd1 vccd1 vccd1 _8285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564_ _4564_/A vssd1 vssd1 vccd1 vccd1 _8315_/D sky130_fd_sc_hd__clkbuf_1
X_7352_ _7384_/A vssd1 vssd1 vccd1 vccd1 _7352_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6303_ _7902_/Q _7901_/Q _6303_/C vssd1 vssd1 vccd1 vccd1 _6306_/C sky130_fd_sc_hd__or3_1
X_7283_ _8629_/Q _7283_/B vssd1 vssd1 vccd1 vccd1 _7331_/C sky130_fd_sc_hd__xor2_1
XFILLER_116_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4495_ _8573_/Q vssd1 vssd1 vccd1 vccd1 _4495_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3015_ clkbuf_0__3015_/X vssd1 vssd1 vccd1 vccd1 _6631_/A sky130_fd_sc_hd__clkbuf_4
X_6234_ _6232_/X _7895_/Q _6225_/X _6229_/X _7863_/Q vssd1 vssd1 vccd1 vccd1 _7863_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6177_/A vssd1 vssd1 vccd1 vccd1 _6172_/B sky130_fd_sc_hd__buf_8
X_5116_ _5095_/X _5102_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__a21o_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _7865_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6096_/X sky130_fd_sc_hd__or2_1
X_5047_ _8228_/Q _4522_/X _5047_/S vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5949_ _7716_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__or2_1
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8599_ _8599_/CLK _8599_/D vssd1 vssd1 vccd1 vccd1 _8599_/Q sky130_fd_sc_hd__dfxtp_1
X_7619_ _8547_/Q vssd1 vssd1 vccd1 vccd1 _7619_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7068__472 _7069__473/A vssd1 vssd1 vccd1 vccd1 _8281_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4280_ _5663_/A _4508_/B _5663_/B vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__or3b_4
XFILLER_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7970_ _8577_/CLK _7970_/D vssd1 vssd1 vccd1 vccd1 _7970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6975__404 _6975__404/A vssd1 vssd1 vccd1 vccd1 _8208_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6852_ _6886_/B _6852_/B vssd1 vssd1 vccd1 vccd1 _7626_/A sky130_fd_sc_hd__nand2_2
XFILLER_35_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7036__449 _7037__450/A vssd1 vssd1 vccd1 vccd1 _8256_/CLK sky130_fd_sc_hd__inv_2
X_5803_ _5803_/A vssd1 vssd1 vccd1 vccd1 _7986_/D sky130_fd_sc_hd__clkbuf_1
X_3995_ _3995_/A vssd1 vssd1 vccd1 vccd1 _8581_/D sky130_fd_sc_hd__clkbuf_1
X_8522_ _8522_/CLK _8522_/D vssd1 vssd1 vccd1 vccd1 _8522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5734_ _8016_/Q _5642_/X _5734_/S vssd1 vssd1 vccd1 vccd1 _5735_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5665_ _5680_/S vssd1 vssd1 vccd1 vccd1 _5674_/S sky130_fd_sc_hd__buf_2
X_8453_ _8453_/CLK _8453_/D vssd1 vssd1 vccd1 vccd1 _8453_/Q sky130_fd_sc_hd__dfxtp_1
X_4616_ _4616_/A vssd1 vssd1 vccd1 vccd1 _8292_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3463_ _7141_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3463_/X sky130_fd_sc_hd__clkbuf_16
X_8384_ _8384_/CLK _8384_/D vssd1 vssd1 vccd1 vccd1 _8384_/Q sky130_fd_sc_hd__dfxtp_1
X_7404_ _7404_/A vssd1 vssd1 vccd1 vccd1 _8441_/D sky130_fd_sc_hd__clkbuf_1
X_5596_ _5593_/X _8079_/Q _5608_/S vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__mux2_1
X_7335_ _7407_/D _7335_/B vssd1 vssd1 vccd1 vccd1 _7335_/X sky130_fd_sc_hd__or2_1
XFILLER_116_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4547_ _4547_/A vssd1 vssd1 vccd1 vccd1 _8321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6611__259 _6611__259/A vssd1 vssd1 vccd1 vccd1 _8019_/CLK sky130_fd_sc_hd__inv_2
X_7266_ _7266_/A _7280_/C _7266_/C vssd1 vssd1 vccd1 vccd1 _7267_/B sky130_fd_sc_hd__and3_1
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4478_ _8188_/Q vssd1 vssd1 vccd1 vccd1 _4478_/X sky130_fd_sc_hd__clkbuf_4
X_7197_ _7448_/A vssd1 vssd1 vccd1 vccd1 _7197_/X sky130_fd_sc_hd__buf_1
XFILLER_100_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6148_ _7954_/Q input12/X _6177_/A vssd1 vssd1 vccd1 vccd1 _6148_/X sky130_fd_sc_hd__mux2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_34 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_12 _6306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_23 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_45 _6188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_67 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_56 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _7861_/Q _6088_/B vssd1 vssd1 vccd1 vccd1 _6079_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_78 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_89 _5205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6692__309 _6693__310/A vssd1 vssd1 vccd1 vccd1 _8077_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3076_ clkbuf_0__3076_/X vssd1 vssd1 vccd1 vccd1 _6327__200/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5450_ _5465_/S vssd1 vssd1 vccd1 vccd1 _5459_/S sky130_fd_sc_hd__buf_2
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4401_ _4123_/X _8370_/Q _4401_/S vssd1 vssd1 vccd1 vccd1 _4402_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5381_ _5381_/A vssd1 vssd1 vccd1 vccd1 _8202_/D sky130_fd_sc_hd__clkbuf_1
X_4332_ _8400_/Q _4235_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ _4278_/S vssd1 vssd1 vccd1 vccd1 _4272_/S sky130_fd_sc_hd__clkbuf_4
X_7051_ _7051_/A vssd1 vssd1 vccd1 vccd1 _7051_/X sky130_fd_sc_hd__buf_1
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6002_ _6002_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__or2_1
X_7042__453 _7044__455/A vssd1 vssd1 vccd1 vccd1 _8260_/CLK sky130_fd_sc_hd__inv_2
X_4194_ _8194_/Q vssd1 vssd1 vccd1 vccd1 _4194_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7953_ _8091_/CLK _7953_/D vssd1 vssd1 vccd1 vccd1 _7953_/Q sky130_fd_sc_hd__dfxtp_1
X_6904_ _8558_/Q _7588_/C _6903_/X vssd1 vssd1 vccd1 vccd1 _6905_/B sky130_fd_sc_hd__a21oi_2
XFILLER_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7884_ _7884_/CLK _7884_/D vssd1 vssd1 vccd1 vccd1 _7884_/Q sky130_fd_sc_hd__dfxtp_1
X_6756__317 _6759__320/A vssd1 vssd1 vccd1 vccd1 _8109_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6835_ _6835_/A _6835_/B _6903_/D vssd1 vssd1 vccd1 vccd1 _7588_/C sky130_fd_sc_hd__or3b_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _6797_/A vssd1 vssd1 vccd1 vccd1 _6766_/X sky130_fd_sc_hd__buf_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3978_ _3977_/X _8586_/Q _3978_/S vssd1 vssd1 vccd1 vccd1 _3979_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3478_ clkbuf_0__3478_/X vssd1 vssd1 vccd1 vccd1 _7221__95/A sky130_fd_sc_hd__clkbuf_4
X_8505_ _8505_/CLK _8505_/D vssd1 vssd1 vccd1 vccd1 _8505_/Q sky130_fd_sc_hd__dfxtp_1
X_5717_ _5717_/A vssd1 vssd1 vccd1 vccd1 _8024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6697_ _6712_/S vssd1 vssd1 vccd1 vccd1 _6706_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _5648_/A vssd1 vssd1 vccd1 vccd1 _8063_/D sky130_fd_sc_hd__clkbuf_1
X_8436_ _8436_/CLK _8436_/D vssd1 vssd1 vccd1 vccd1 _8436_/Q sky130_fd_sc_hd__dfxtp_1
X_5579_ _5404_/X _8110_/Q _5585_/S vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__mux2_1
X_8367_ _8367_/CLK _8367_/D vssd1 vssd1 vccd1 vccd1 _8367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8298_ _8298_/CLK _8298_/D vssd1 vssd1 vccd1 vccd1 _8298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7318_ _7318_/A _7350_/A vssd1 vssd1 vccd1 vccd1 _7319_/C sky130_fd_sc_hd__nand2_1
XFILLER_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7249_ _8438_/Q _7306_/B vssd1 vssd1 vccd1 vccd1 _7250_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7460__135 _7460__135/A vssd1 vssd1 vccd1 vccd1 _8474_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _8279_/Q _4849_/X _4847_/X _8241_/Q vssd1 vssd1 vccd1 vccd1 _4950_/X sky130_fd_sc_hd__a22o_1
X_4881_ _4853_/X _7930_/Q _7855_/Q _4829_/X _4809_/A vssd1 vssd1 vccd1 vccd1 _4881_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3901_ _5382_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5383_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6551_ _8094_/Q _7979_/Q _6804_/S vssd1 vssd1 vccd1 vccd1 _6552_/A sky130_fd_sc_hd__mux2_1
X_5502_ _5502_/A vssd1 vssd1 vccd1 vccd1 _8147_/D sky130_fd_sc_hd__clkbuf_1
X_6482_ _7951_/Q _6464_/X _6474_/X _6481_/X _6472_/X vssd1 vssd1 vccd1 vccd1 _7951_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5433_ _5398_/X _8179_/Q _5441_/S vssd1 vssd1 vccd1 vccd1 _5434_/A sky130_fd_sc_hd__mux2_1
X_8221_ _8221_/CLK _8221_/D vssd1 vssd1 vccd1 vccd1 _8221_/Q sky130_fd_sc_hd__dfxtp_2
X_8152_ _8152_/CLK _8152_/D vssd1 vssd1 vccd1 vccd1 _8152_/Q sky130_fd_sc_hd__dfxtp_1
X_5364_ _5189_/A _5360_/X _5363_/X _5204_/A vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__a211o_1
X_8645__210 vssd1 vssd1 vccd1 vccd1 _8645__210/HI caravel_irq[1] sky130_fd_sc_hd__conb_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4315_ _4315_/A vssd1 vssd1 vccd1 vccd1 _8408_/D sky130_fd_sc_hd__clkbuf_1
X_7103_ _7134_/A vssd1 vssd1 vccd1 vccd1 _7103_/X sky130_fd_sc_hd__buf_1
XFILLER_99_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5295_ _5254_/X _8157_/Q _7922_/Q _5230_/B _5239_/X vssd1 vssd1 vccd1 vccd1 _5295_/X
+ sky130_fd_sc_hd__o221a_1
X_8083_ _8625_/CLK _8083_/D vssd1 vssd1 vccd1 vccd1 _8083_/Q sky130_fd_sc_hd__dfxtp_1
X_4246_ _4246_/A vssd1 vssd1 vccd1 vccd1 _8467_/D sky130_fd_sc_hd__clkbuf_1
X_4177_ _4179_/C vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7936_ _8452_/CLK _7936_/D vssd1 vssd1 vccd1 vccd1 _7936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7867_ _8631_/CLK _7867_/D vssd1 vssd1 vccd1 vccd1 _7867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7798_ _7798_/A _7811_/B vssd1 vssd1 vccd1 vccd1 _7798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6749_ _6749_/A vssd1 vssd1 vccd1 vccd1 _8103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7049__459 _7049__459/A vssd1 vssd1 vccd1 vccd1 _8266_/CLK sky130_fd_sc_hd__inv_2
X_8419_ _8419_/CLK _8419_/D vssd1 vssd1 vccd1 vccd1 _8419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4100_ _4100_/A vssd1 vssd1 vccd1 vccd1 _8502_/D sky130_fd_sc_hd__clkbuf_1
X_5080_ _5081_/A vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4031_ _4031_/A vssd1 vssd1 vccd1 vccd1 _8532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5982_ _5982_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__or2_1
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4933_ _4475_/X _4669_/A _4932_/X _4903_/X vssd1 vssd1 vccd1 vccd1 _8262_/D sky130_fd_sc_hd__o211a_1
X_7721_ _7828_/A _7723_/B _7723_/C vssd1 vssd1 vccd1 vccd1 _7722_/A sky130_fd_sc_hd__and3_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4864_ _4861_/X _4862_/X _4863_/X vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__o21a_1
X_7652_ _7651_/X _7662_/B vssd1 vssd1 vccd1 vccd1 _7653_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4795_ _7908_/Q _8028_/Q _8044_/Q _8012_/Q _4710_/A _4694_/A vssd1 vssd1 vccd1 vccd1
+ _4796_/B sky130_fd_sc_hd__mux4_1
X_7583_ _7548_/A _7549_/B _6869_/X _6864_/Y _7582_/Y vssd1 vssd1 vccd1 vccd1 _7593_/B
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3315_ clkbuf_0__3315_/X vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__clkbuf_4
X_6534_ _6534_/A vssd1 vssd1 vccd1 vccd1 _7971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3246_ clkbuf_0__3246_/X vssd1 vssd1 vccd1 vccd1 _6575__230/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6465_ _8622_/Q vssd1 vssd1 vccd1 vccd1 _7808_/A sky130_fd_sc_hd__clkbuf_4
X_5416_ _5607_/A vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__clkbuf_2
X_8204_ _8204_/CLK _8204_/D vssd1 vssd1 vccd1 vccd1 _8204_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput120 _6013_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__buf_2
Xoutput131 _6020_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput142 _5970_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__buf_2
X_6396_ _6396_/A vssd1 vssd1 vccd1 vccd1 _7055_/B sky130_fd_sc_hd__clkbuf_2
Xoutput153 _5992_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput164 _5950_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__buf_2
Xoutput175 _5927_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__buf_2
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7161__547 _7162__548/A vssd1 vssd1 vccd1 vccd1 _8356_/CLK sky130_fd_sc_hd__inv_2
X_8135_ _8135_/CLK _8135_/D vssd1 vssd1 vccd1 vccd1 _8135_/Q sky130_fd_sc_hd__dfxtp_1
X_5347_ _5269_/X _5345_/X _5346_/X vssd1 vssd1 vccd1 vccd1 _5351_/B sky130_fd_sc_hd__o21a_1
Xoutput186 _6151_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8066_ _8066_/CLK _8066_/D vssd1 vssd1 vccd1 vccd1 _8066_/Q sky130_fd_sc_hd__dfxtp_1
X_5278_ _5274_/X _5275_/X _5277_/X _5142_/S vssd1 vssd1 vccd1 vccd1 _5279_/C sky130_fd_sc_hd__o211a_1
Xoutput197 _6183_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _8573_/Q vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3076_ _6322_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3076_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3462_ clkbuf_0__3462_/X vssd1 vssd1 vccd1 vccd1 _7139__529/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7919_ _7919_/CLK _7919_/D vssd1 vssd1 vccd1 vccd1 _7919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6769__327 _6769__327/A vssd1 vssd1 vccd1 vccd1 _8119_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7062__467 _7063__468/A vssd1 vssd1 vccd1 vccd1 _8276_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7725__27 _7728__30/A vssd1 vssd1 vccd1 vccd1 _8578_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _6180_/A sky130_fd_sc_hd__clkbuf_4
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
X_4580_ _4580_/A vssd1 vssd1 vccd1 vccd1 _8308_/D sky130_fd_sc_hd__clkbuf_1
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
Xinput55 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _3904_/B sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _3907_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _6025_/A sky130_fd_sc_hd__buf_4
Xinput88 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__buf_4
Xinput77 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__buf_4
Xinput99 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _7723_/A sky130_fd_sc_hd__buf_4
X_6250_ _6249_/X _8083_/Q _6245_/X _6247_/X _7872_/Q vssd1 vssd1 vccd1 vccd1 _7872_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5201_ _8598_/Q _8151_/Q _8124_/Q _8582_/Q _5330_/S _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5201_/X sky130_fd_sc_hd__mux4_2
X_6181_ _7888_/Q _6175_/X _6176_/X _6180_/X _6173_/X vssd1 vssd1 vccd1 vccd1 _6181_/X
+ sky130_fd_sc_hd__o221a_1
X_5132_ _8593_/Q _8342_/Q _8326_/Q _8366_/Q _5130_/X _5131_/X vssd1 vssd1 vccd1 vccd1
+ _5133_/B sky130_fd_sc_hd__mux4_1
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5063_ _5063_/A vssd1 vssd1 vccd1 vccd1 _8222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4014_ _4014_/A vssd1 vssd1 vccd1 vccd1 _8538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5965_ _7809_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__or2_1
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5896_ _4212_/X _7853_/Q _5896_/S vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__mux2_1
X_4916_ _4911_/X _4912_/X _4915_/X _4706_/X vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7704_ _8569_/Q _7704_/B vssd1 vssd1 vccd1 vccd1 _7704_/X sky130_fd_sc_hd__or2_1
X_4847_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4847_/X sky130_fd_sc_hd__buf_2
X_7635_ _7634_/Y _7620_/X _7625_/X _6869_/B vssd1 vssd1 vccd1 vccd1 _7635_/X sky130_fd_sc_hd__o22a_1
X_4778_ _7850_/Q _7858_/Q _7933_/Q _8037_/Q _4721_/X _4725_/X vssd1 vssd1 vccd1 vccd1
+ _4778_/X sky130_fd_sc_hd__mux4_1
X_7566_ _8626_/Q _7566_/B _7566_/C vssd1 vssd1 vccd1 vccd1 _7566_/X sky130_fd_sc_hd__and3_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6517_ _6550_/A vssd1 vssd1 vccd1 vccd1 _6526_/S sky130_fd_sc_hd__clkbuf_2
X_6448_ _7817_/A _6481_/C _6448_/C _6474_/A vssd1 vssd1 vccd1 vccd1 _6448_/X sky130_fd_sc_hd__and4_1
XFILLER_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6379_ _6379_/A _6433_/A _7790_/C _6371_/B vssd1 vssd1 vccd1 vccd1 _6384_/B sky130_fd_sc_hd__or4b_1
X_8118_ _8118_/CLK _8118_/D vssd1 vssd1 vccd1 vccd1 _8118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8049_ _8052_/CLK _8049_/D vssd1 vssd1 vccd1 vccd1 _8049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3445_ clkbuf_0__3445_/X vssd1 vssd1 vccd1 vccd1 _7058__464/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7346__112 _7347__113/A vssd1 vssd1 vccd1 vccd1 _8423_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8612_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6669__291 _6672__294/A vssd1 vssd1 vccd1 vccd1 _8059_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5750_ _8009_/Q _5639_/X _5752_/S vssd1 vssd1 vccd1 vccd1 _5751_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4701_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__buf_2
X_5681_ _5681_/A vssd1 vssd1 vccd1 vccd1 _8040_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4632_ _4460_/X _8285_/Q _4638_/S vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__mux2_1
X_7420_ _7420_/A vssd1 vssd1 vccd1 vccd1 _7420_/X sky130_fd_sc_hd__clkbuf_2
X_4563_ _8315_/Q _4519_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__mux2_1
X_7351_ _7407_/D _7335_/B _7350_/B vssd1 vssd1 vccd1 vccd1 _7384_/A sky130_fd_sc_hd__a21o_1
X_4494_ _4494_/A vssd1 vssd1 vccd1 vccd1 _8339_/D sky130_fd_sc_hd__clkbuf_1
X_6302_ _7902_/Q _7901_/Q vssd1 vssd1 vccd1 vccd1 _6304_/B sky130_fd_sc_hd__nand2_1
X_7282_ _7282_/A _7282_/B vssd1 vssd1 vccd1 vccd1 _7283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3014_ clkbuf_0__3014_/X vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__clkbuf_4
X_6233_ _6232_/X _7894_/Q _6225_/X _6229_/X _7862_/Q vssd1 vssd1 vccd1 vccd1 _7862_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _7882_/Q _6159_/X _6160_/X _6163_/X _6157_/X vssd1 vssd1 vccd1 vccd1 _6164_/X
+ sky130_fd_sc_hd__o221a_1
X_5115_ _5391_/B _5111_/X _5344_/A vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__a21o_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _7940_/Q input29/X _6106_/S vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__mux2_1
X_5046_ _5046_/A vssd1 vssd1 vccd1 vccd1 _8229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5948_ _5948_/A vssd1 vssd1 vccd1 vccd1 _5948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5879_ _5879_/A vssd1 vssd1 vccd1 vccd1 _7904_/D sky130_fd_sc_hd__clkbuf_1
X_8598_ _8598_/CLK _8598_/D vssd1 vssd1 vccd1 vccd1 _8598_/Q sky130_fd_sc_hd__dfxtp_1
X_7618_ _7618_/A vssd1 vssd1 vccd1 vccd1 _8546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7549_ _8620_/Q _7549_/B vssd1 vssd1 vccd1 vccd1 _7550_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3428_ clkbuf_0__3428_/X vssd1 vssd1 vccd1 vccd1 _6982__410/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7075__477 _7075__477/A vssd1 vssd1 vccd1 vccd1 _8286_/CLK sky130_fd_sc_hd__inv_2
X_6851_ _8548_/Q _8547_/Q vssd1 vssd1 vccd1 vccd1 _6852_/B sky130_fd_sc_hd__and2_1
X_5802_ _7986_/Q _5610_/A _5806_/S vssd1 vssd1 vccd1 vccd1 _5803_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7537__22 _7537__22/A vssd1 vssd1 vccd1 vccd1 _8536_/CLK sky130_fd_sc_hd__inv_2
X_8521_ _8521_/CLK _8521_/D vssd1 vssd1 vccd1 vccd1 _8521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3994_ _3968_/X _8581_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _5733_/A vssd1 vssd1 vccd1 vccd1 _8017_/D sky130_fd_sc_hd__clkbuf_1
X_5664_ _5808_/A _5862_/B vssd1 vssd1 vccd1 vccd1 _5680_/S sky130_fd_sc_hd__or2_2
X_8452_ _8452_/CLK _8452_/D vssd1 vssd1 vccd1 vccd1 _8452_/Q sky130_fd_sc_hd__dfxtp_1
X_4615_ _8292_/Q _4489_/X _4619_/S vssd1 vssd1 vccd1 vccd1 _4616_/A sky130_fd_sc_hd__mux2_1
X_5595_ _5617_/S vssd1 vssd1 vccd1 vccd1 _5608_/S sky130_fd_sc_hd__buf_2
X_8383_ _8383_/CLK _8383_/D vssd1 vssd1 vccd1 vccd1 _8383_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3462_ _7135_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3462_/X sky130_fd_sc_hd__clkbuf_16
X_7403_ _7401_/X _7432_/S _7403_/C vssd1 vssd1 vccd1 vccd1 _7404_/A sky130_fd_sc_hd__and3b_1
X_4546_ _4444_/X _8321_/Q _4550_/S vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__mux2_1
X_7334_ _8415_/Q _7334_/B _7334_/C _7334_/D vssd1 vssd1 vccd1 vccd1 _7335_/B sky130_fd_sc_hd__and4_1
XFILLER_104_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7170__53 _7172__55/A vssd1 vssd1 vccd1 vccd1 _8362_/CLK sky130_fd_sc_hd__inv_2
X_4477_ _4477_/A vssd1 vssd1 vccd1 vccd1 _8344_/D sky130_fd_sc_hd__clkbuf_1
X_7265_ _8434_/Q _8433_/Q vssd1 vssd1 vccd1 vccd1 _7266_/C sky130_fd_sc_hd__and2_1
X_6147_ _6147_/A vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__buf_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_13 _8364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_35 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_68 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6078_ _6149_/A vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__buf_4
XINSDIODE2_57 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_46 _6188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5029_ _8236_/Q _4522_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_79 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7225__98 _7226__99/A vssd1 vssd1 vccd1 vccd1 _8407_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6579__233 _6581__235/A vssd1 vssd1 vccd1 vccd1 _7993_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8662__227 vssd1 vssd1 vccd1 vccd1 _8662__227/HI core1Index[7] sky130_fd_sc_hd__conb_1
XFILLER_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6219__191 _6219__191/A vssd1 vssd1 vccd1 vccd1 _7860_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4400_ _4400_/A vssd1 vssd1 vccd1 vccd1 _8371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5380_ _5376_/B _5380_/B _6986_/B vssd1 vssd1 vccd1 vccd1 _5381_/A sky130_fd_sc_hd__and3b_1
XFILLER_113_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4331_ _4331_/A vssd1 vssd1 vccd1 vccd1 _8401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _5645_/A _5862_/A vssd1 vssd1 vccd1 vccd1 _4278_/S sky130_fd_sc_hd__nor2_2
X_6001_ _6001_/A vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _4193_/A vssd1 vssd1 vccd1 vccd1 _8484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7952_ _8091_/CLK _7952_/D vssd1 vssd1 vccd1 vccd1 _7952_/Q sky130_fd_sc_hd__dfxtp_1
X_6903_ _8558_/Q _8557_/Q _8556_/Q _6903_/D vssd1 vssd1 vccd1 vccd1 _6903_/X sky130_fd_sc_hd__and4b_1
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7883_ _7884_/CLK _7883_/D vssd1 vssd1 vccd1 vccd1 _7883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _8556_/Q vssd1 vssd1 vccd1 vccd1 _6835_/B sky130_fd_sc_hd__inv_2
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3977_ _8570_/Q vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3477_ clkbuf_0__3477_/X vssd1 vssd1 vccd1 vccd1 _7215__90/A sky130_fd_sc_hd__clkbuf_4
X_8504_ _8504_/CLK _8504_/D vssd1 vssd1 vccd1 vccd1 _8504_/Q sky130_fd_sc_hd__dfxtp_1
X_5716_ _5616_/X _8024_/Q _5716_/S vssd1 vssd1 vccd1 vccd1 _5717_/A sky130_fd_sc_hd__mux2_1
X_8435_ _8436_/CLK _8435_/D vssd1 vssd1 vccd1 vccd1 _8435_/Q sky130_fd_sc_hd__dfxtp_1
X_6696_ _6696_/A _6732_/B vssd1 vssd1 vccd1 vccd1 _6712_/S sky130_fd_sc_hd__nand2_2
X_5647_ _5593_/X _8063_/Q _5655_/S vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__mux2_1
X_6320__194 _6321__195/A vssd1 vssd1 vccd1 vccd1 _7906_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5578_ _5578_/A vssd1 vssd1 vccd1 vccd1 _8111_/D sky130_fd_sc_hd__clkbuf_1
X_8366_ _8366_/CLK _8366_/D vssd1 vssd1 vccd1 vccd1 _8366_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3445_ _7051_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3445_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7125__518 _7127__520/A vssd1 vssd1 vccd1 vccd1 _8327_/CLK sky130_fd_sc_hd__inv_2
X_4529_ _8328_/Q _4528_/X _4532_/S vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7317_ _7399_/B _7350_/A _7430_/B _7318_/A vssd1 vssd1 vccd1 vccd1 _7319_/B sky130_fd_sc_hd__a211o_1
X_8297_ _8297_/CLK _8297_/D vssd1 vssd1 vccd1 vccd1 _8297_/Q sky130_fd_sc_hd__dfxtp_1
X_7248_ _7244_/A _7394_/B _8619_/Q vssd1 vssd1 vccd1 vccd1 _7252_/A sky130_fd_sc_hd__a21bo_1
X_7179_ _7191_/A vssd1 vssd1 vccd1 vccd1 _7179_/X sky130_fd_sc_hd__buf_1
XFILLER_105_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7531__17 _7532__18/A vssd1 vssd1 vccd1 vccd1 _8531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4880_ _8329_/Q _4817_/X _4723_/A _4879_/X vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__o211a_1
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3900_ _8215_/Q _3981_/A vssd1 vssd1 vccd1 vccd1 _5382_/B sky130_fd_sc_hd__and2_1
XFILLER_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6550_ _6550_/A vssd1 vssd1 vccd1 vccd1 _6804_/S sky130_fd_sc_hd__clkbuf_4
X_5501_ _8147_/Q _4504_/X _5501_/S vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6481_ _7793_/A _6490_/B _6481_/C vssd1 vssd1 vccd1 vccd1 _6481_/X sky130_fd_sc_hd__and3_1
X_5432_ _5447_/S vssd1 vssd1 vccd1 vccd1 _5441_/S sky130_fd_sc_hd__buf_2
X_8220_ _8220_/CLK _8220_/D vssd1 vssd1 vccd1 vccd1 _8220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8151_ _8151_/CLK _8151_/D vssd1 vssd1 vccd1 vccd1 _8151_/Q sky130_fd_sc_hd__dfxtp_1
X_5363_ _5274_/X _5361_/X _5362_/X vssd1 vssd1 vccd1 vccd1 _5363_/X sky130_fd_sc_hd__o21a_1
X_4314_ _8408_/Q _4235_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__mux2_1
X_5294_ _5294_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5294_/X sky130_fd_sc_hd__or2_1
X_8082_ _8625_/CLK _8082_/D vssd1 vssd1 vccd1 vccd1 _8082_/Q sky130_fd_sc_hd__dfxtp_1
X_4245_ _8467_/Q _4220_/X _4251_/S vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__mux2_1
X_6762__322 _6763__323/A vssd1 vssd1 vccd1 vccd1 _8114_/CLK sky130_fd_sc_hd__inv_2
X_7437__116 _7438__117/A vssd1 vssd1 vccd1 vccd1 _8455_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4176_ _8257_/Q _8256_/Q _8255_/Q vssd1 vssd1 vccd1 vccd1 _4179_/C sky130_fd_sc_hd__and3_1
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7935_ _7935_/CLK _7935_/D vssd1 vssd1 vccd1 vccd1 _7935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7866_ _8439_/CLK _7866_/D vssd1 vssd1 vccd1 vccd1 _7866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7797_ _7793_/Y _7796_/Y _7757_/A vssd1 vssd1 vccd1 vccd1 _8618_/D sky130_fd_sc_hd__a21oi_1
XFILLER_109_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6914__369 _6915__370/A vssd1 vssd1 vccd1 vccd1 _8165_/CLK sky130_fd_sc_hd__inv_2
X_6748_ _8103_/Q _6008_/A _6748_/S vssd1 vssd1 vccd1 vccd1 _6749_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8418_ _8418_/CLK _8418_/D vssd1 vssd1 vccd1 vccd1 _8418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8349_ _8349_/CLK _8349_/D vssd1 vssd1 vccd1 vccd1 _8349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3428_ _6977_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3428_/X sky130_fd_sc_hd__clkbuf_16
X_7340__107 _7342__109/A vssd1 vssd1 vccd1 vccd1 _8418_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8668__233 vssd1 vssd1 vccd1 vccd1 _8668__233/HI manufacturerID[5] sky130_fd_sc_hd__conb_1
XFILLER_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4030_ _3952_/X _8532_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4031_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ _5981_/A vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4932_ _4671_/X _8262_/Q _4741_/X _4931_/X vssd1 vssd1 vccd1 vccd1 _4932_/X sky130_fd_sc_hd__a211o_1
X_7720_ _7720_/A vssd1 vssd1 vccd1 vccd1 _8575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7651_ _6838_/Y _7642_/X _7647_/X _7548_/B vssd1 vssd1 vccd1 vccd1 _7651_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4863_ _4855_/A _7987_/Q _4865_/A _8220_/Q _4724_/A vssd1 vssd1 vccd1 vccd1 _4863_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4794_ _4713_/X _4791_/X _4793_/X vssd1 vssd1 vccd1 vccd1 _4794_/X sky130_fd_sc_hd__a21o_1
X_7582_ _7582_/A _7582_/B vssd1 vssd1 vccd1 vccd1 _7582_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3314_ clkbuf_0__3314_/X vssd1 vssd1 vccd1 vccd1 _6796__350/A sky130_fd_sc_hd__clkbuf_4
X_6533_ _6041_/A _7971_/Q _6537_/S vssd1 vssd1 vccd1 vccd1 _6534_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3245_ clkbuf_0__3245_/X vssd1 vssd1 vccd1 vccd1 _6594_/A sky130_fd_sc_hd__clkbuf_4
X_6464_ _6483_/A vssd1 vssd1 vccd1 vccd1 _6464_/X sky130_fd_sc_hd__clkbuf_2
Xoutput110 _6033_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__buf_2
X_5415_ _8191_/Q vssd1 vssd1 vccd1 vccd1 _5607_/A sky130_fd_sc_hd__buf_2
X_8203_ _8203_/CLK _8203_/D vssd1 vssd1 vccd1 vccd1 _8203_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput121 _6055_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput132 _6022_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__buf_2
Xoutput143 _5972_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8439_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6395_ _6403_/A vssd1 vssd1 vccd1 vccd1 _6395_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput154 _5994_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput165 _5953_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__buf_2
X_8134_ _8134_/CLK _8134_/D vssd1 vssd1 vccd1 vccd1 _8134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5346_ _8391_/Q _5271_/X _5238_/A _8383_/Q _5239_/A vssd1 vssd1 vccd1 vccd1 _5346_/X
+ sky130_fd_sc_hd__o221a_1
Xoutput176 _6192_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8065_ _8065_/CLK _8065_/D vssd1 vssd1 vccd1 vccd1 _8065_/Q sky130_fd_sc_hd__dfxtp_1
X_5277_ _8361_/Q _5276_/X _5249_/A _8588_/Q vssd1 vssd1 vccd1 vccd1 _5277_/X sky130_fd_sc_hd__o22a_1
Xoutput198 _6185_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput187 _6154_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__buf_2
X_4228_ _4228_/A vssd1 vssd1 vccd1 vccd1 _8473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3461_ clkbuf_0__3461_/X vssd1 vssd1 vccd1 vccd1 _7159_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4159_ _8259_/Q vssd1 vssd1 vccd1 vccd1 _5663_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7918_ _7918_/CLK _7918_/D vssd1 vssd1 vccd1 vccd1 _7918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7849_ _7849_/CLK _7849_/D vssd1 vssd1 vccd1 vccd1 _7849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3659_ clkbuf_0__3659_/X vssd1 vssd1 vccd1 vccd1 _7519__7/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7138__528 _7139__529/A vssd1 vssd1 vccd1 vccd1 _8337_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__3322_ clkbuf_0__3322_/X vssd1 vssd1 vccd1 vccd1 _6915__370/A sky130_fd_sc_hd__clkbuf_16
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _6182_/A sky130_fd_sc_hd__clkbuf_4
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_4
Xinput45 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__clkbuf_1
Xinput56 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__clkbuf_1
Xinput67 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _6028_/A sky130_fd_sc_hd__buf_4
Xinput78 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__buf_4
Xinput89 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__buf_4
X_5200_ _7924_/Q _8132_/Q _8411_/Q _8159_/Q _5313_/S _5110_/X vssd1 vssd1 vccd1 vccd1
+ _5200_/X sky130_fd_sc_hd__mux4_2
X_6180_ _6180_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6180_/X sky130_fd_sc_hd__and2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _5221_/A vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__clkbuf_4
X_8642__258 vssd1 vssd1 vccd1 vccd1 partID[14] _8642__258/LO sky130_fd_sc_hd__conb_1
XFILLER_97_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5062_ _4463_/X _8222_/Q _5066_/S vssd1 vssd1 vccd1 vccd1 _5063_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4013_ _8538_/Q _3934_/X _4017_/S vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5964_ _5964_/A vssd1 vssd1 vccd1 vccd1 _5964_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7703_ _8569_/Q _7687_/A _7702_/X _7684_/A vssd1 vssd1 vccd1 vccd1 _8568_/D sky130_fd_sc_hd__o211a_1
X_5895_ _5895_/A vssd1 vssd1 vccd1 vccd1 _7854_/D sky130_fd_sc_hd__clkbuf_1
X_4915_ _7905_/Q _4838_/X _4913_/X _4914_/X vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _4852_/A vssd1 vssd1 vccd1 vccd1 _4847_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7177__59 _7177__59/A vssd1 vssd1 vccd1 vccd1 _8368_/CLK sky130_fd_sc_hd__inv_2
X_7634_ _8550_/Q vssd1 vssd1 vccd1 vccd1 _7634_/Y sky130_fd_sc_hd__inv_2
X_6573__228 _6575__230/A vssd1 vssd1 vccd1 vccd1 _7988_/CLK sky130_fd_sc_hd__inv_2
X_7565_ _7590_/A _7551_/Y _7562_/X _7563_/Y _7564_/Y vssd1 vssd1 vccd1 vccd1 _7565_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4777_ _4796_/A _4777_/B vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__and2_1
X_6516_ _6516_/A vssd1 vssd1 vccd1 vccd1 _7963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6447_ _8625_/Q vssd1 vssd1 vccd1 vccd1 _7817_/A sky130_fd_sc_hd__clkbuf_4
X_6378_ _7790_/A vssd1 vssd1 vccd1 vccd1 _6379_/A sky130_fd_sc_hd__clkinv_2
X_8117_ _8117_/CLK _8117_/D vssd1 vssd1 vccd1 vccd1 _8117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5329_ _5274_/X _5327_/X _5328_/X vssd1 vssd1 vccd1 vccd1 _5333_/B sky130_fd_sc_hd__o21ai_1
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8048_ _8608_/CLK _8048_/D vssd1 vssd1 vccd1 vccd1 _8048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6213__186 _6217__190/A vssd1 vssd1 vccd1 vccd1 _7855_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3444_ clkbuf_0__3444_/X vssd1 vssd1 vccd1 vccd1 _7050__460/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6775__332 _6776__333/A vssd1 vssd1 vccd1 vccd1 _8124_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7730__31 _7732__33/A vssd1 vssd1 vccd1 vccd1 _8582_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6927__379 _6927__379/A vssd1 vssd1 vccd1 vccd1 _8175_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6823__366 _6824__367/A vssd1 vssd1 vccd1 vccd1 _8161_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4700_ _4955_/S vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__clkbuf_4
X_5680_ _5616_/X _8040_/Q _5680_/S vssd1 vssd1 vccd1 vccd1 _5681_/A sky130_fd_sc_hd__mux2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4631_ _4631_/A vssd1 vssd1 vccd1 vccd1 _8286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4562_ _4562_/A vssd1 vssd1 vccd1 vccd1 _8316_/D sky130_fd_sc_hd__clkbuf_1
X_7350_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7350_/Y sky130_fd_sc_hd__nor2_1
X_4493_ _8339_/Q _4492_/X _4496_/S vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__mux2_1
X_7281_ _7279_/Y _7379_/A _7267_/B vssd1 vssd1 vccd1 vccd1 _7281_/X sky130_fd_sc_hd__a21o_1
X_6301_ _7902_/Q _6299_/X _7760_/A vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__o21a_1
X_6232_ _6423_/A vssd1 vssd1 vccd1 vccd1 _6232_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6176_/A vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5114_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5344_/A sky130_fd_sc_hd__clkbuf_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6073_/X _6091_/X _6093_/X _6082_/X vssd1 vssd1 vccd1 vccd1 _6094_/X sky130_fd_sc_hd__o211a_1
X_5045_ _8229_/Q _4519_/X _5047_/S vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5947_ _7714_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__or2_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5878_ _7904_/Q _5616_/A _5878_/S vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__mux2_1
X_7617_ _7616_/X _7628_/B vssd1 vssd1 vccd1 vccd1 _7618_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4829_ _4874_/A vssd1 vssd1 vccd1 vccd1 _4829_/X sky130_fd_sc_hd__buf_2
X_8597_ _8597_/CLK _8597_/D vssd1 vssd1 vccd1 vccd1 _8597_/Q sky130_fd_sc_hd__dfxtp_1
X_7548_ _7548_/A _7548_/B vssd1 vssd1 vccd1 vccd1 _7550_/A sky130_fd_sc_hd__xnor2_1
XFILLER_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7479_ _7479_/A vssd1 vssd1 vccd1 vccd1 _7479_/X sky130_fd_sc_hd__buf_1
XFILLER_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3427_ clkbuf_0__3427_/X vssd1 vssd1 vccd1 vccd1 _6976__405/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6850_ _6850_/A vssd1 vssd1 vccd1 vccd1 _6886_/B sky130_fd_sc_hd__buf_2
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5801_ _5801_/A vssd1 vssd1 vccd1 vccd1 _7987_/D sky130_fd_sc_hd__clkbuf_1
X_5732_ _8017_/Q _5639_/X _5734_/S vssd1 vssd1 vccd1 vccd1 _5733_/A sky130_fd_sc_hd__mux2_1
X_8520_ _8520_/CLK _8520_/D vssd1 vssd1 vccd1 vccd1 _8520_/Q sky130_fd_sc_hd__dfxtp_1
X_3993_ _3993_/A vssd1 vssd1 vccd1 vccd1 _8582_/D sky130_fd_sc_hd__clkbuf_1
X_8451_ _8604_/CLK _8451_/D vssd1 vssd1 vccd1 vccd1 _8451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5663_ _5663_/A _5663_/B _4508_/B vssd1 vssd1 vccd1 vccd1 _5862_/B sky130_fd_sc_hd__or3b_4
X_8382_ _8382_/CLK _8382_/D vssd1 vssd1 vccd1 vccd1 _8382_/Q sky130_fd_sc_hd__dfxtp_1
X_4614_ _4614_/A vssd1 vssd1 vccd1 vccd1 _8293_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3461_ _7134_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3461_/X sky130_fd_sc_hd__clkbuf_16
X_5594_ _5594_/A _5808_/A vssd1 vssd1 vccd1 vccd1 _5617_/S sky130_fd_sc_hd__or2_2
X_7402_ _7407_/D _7350_/A _7399_/Y _8441_/Q vssd1 vssd1 vccd1 vccd1 _7403_/C sky130_fd_sc_hd__a31o_1
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _8322_/D sky130_fd_sc_hd__clkbuf_1
X_7333_ _7328_/X _7329_/Y _7330_/X _7331_/X _7332_/X vssd1 vssd1 vccd1 vccd1 _7334_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4476_ _4475_/X _8344_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__mux2_1
X_7264_ _8623_/Q vssd1 vssd1 vccd1 vccd1 _7589_/A sky130_fd_sc_hd__inv_2
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6146_ _6136_/X _6144_/X _6145_/X _6139_/X vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__o211a_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_14 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6077_ _6077_/A vssd1 vssd1 vccd1 vccd1 _6149_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_58 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_36 _6160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_47 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5028_ _5028_/A vssd1 vssd1 vccd1 vccd1 _8237_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_69 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7543__26 _7543__26/A vssd1 vssd1 vccd1 vccd1 _8540_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3659_ _7517_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3659_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6332__203 _6334__205/A vssd1 vssd1 vccd1 vccd1 _7915_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4330_ _8401_/Q _4232_/X _4334_/S vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4261_ _5898_/A vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__clkbuf_4
X_6000_ _6000_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__or2_1
X_7081__482 _7084__485/A vssd1 vssd1 vccd1 vccd1 _8291_/CLK sky130_fd_sc_hd__inv_2
X_4192_ _8484_/Q _4156_/X _4204_/S vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7951_ _8622_/CLK _7951_/D vssd1 vssd1 vccd1 vccd1 _7951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6902_ _6885_/X _6896_/Y _7586_/C _6902_/D vssd1 vssd1 vccd1 vccd1 _6909_/B sky130_fd_sc_hd__and4bb_1
X_7882_ _8091_/CLK _7882_/D vssd1 vssd1 vccd1 vccd1 _7882_/Q sky130_fd_sc_hd__dfxtp_1
X_6833_ _8557_/Q vssd1 vssd1 vccd1 vccd1 _6835_/A sky130_fd_sc_hd__inv_2
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3976_ _3976_/A vssd1 vssd1 vccd1 vccd1 _8587_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3476_ clkbuf_0__3476_/X vssd1 vssd1 vccd1 vccd1 _7209__85/A sky130_fd_sc_hd__clkbuf_4
X_5715_ _5715_/A vssd1 vssd1 vccd1 vccd1 _8025_/D sky130_fd_sc_hd__clkbuf_1
X_8503_ _8503_/CLK _8503_/D vssd1 vssd1 vccd1 vccd1 _8503_/Q sky130_fd_sc_hd__dfxtp_1
X_5646_ _5661_/S vssd1 vssd1 vccd1 vccd1 _5655_/S sky130_fd_sc_hd__buf_2
X_8434_ _8441_/CLK _8434_/D vssd1 vssd1 vccd1 vccd1 _8434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5577_ _5398_/X _8111_/Q _5585_/S vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__mux2_1
X_8365_ _8365_/CLK _8365_/D vssd1 vssd1 vccd1 vccd1 _8365_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3444_ _7045_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3444_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4528_ _8189_/Q vssd1 vssd1 vccd1 vccd1 _4528_/X sky130_fd_sc_hd__clkbuf_4
X_8296_ _8296_/CLK _8296_/D vssd1 vssd1 vccd1 vccd1 _8296_/Q sky130_fd_sc_hd__dfxtp_1
X_7316_ _7410_/A _7412_/A vssd1 vssd1 vccd1 vccd1 _7430_/B sky130_fd_sc_hd__nor2_2
X_4459_ _4459_/A vssd1 vssd1 vccd1 vccd1 _8350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7247_ _8438_/Q _7306_/B _8439_/Q vssd1 vssd1 vccd1 vccd1 _7394_/B sky130_fd_sc_hd__a21o_1
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6129_ _7949_/Q input7/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6129_/X sky130_fd_sc_hd__mux2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7019__435 _7019__435/A vssd1 vssd1 vccd1 vccd1 _8241_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5500_ _5500_/A vssd1 vssd1 vccd1 vccd1 _8148_/D sky130_fd_sc_hd__clkbuf_1
X_6339__209 _6340__210/A vssd1 vssd1 vccd1 vccd1 _7921_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ _8618_/Q vssd1 vssd1 vccd1 vccd1 _7793_/A sky130_fd_sc_hd__buf_2
X_5431_ _5898_/A _5772_/B vssd1 vssd1 vccd1 vccd1 _5447_/S sky130_fd_sc_hd__or2_2
X_8150_ _8150_/CLK _8150_/D vssd1 vssd1 vccd1 vccd1 _8150_/Q sky130_fd_sc_hd__dfxtp_1
X_5362_ _8493_/Q _5271_/X _5238_/A _8485_/Q _5239_/A vssd1 vssd1 vccd1 vccd1 _5362_/X
+ sky130_fd_sc_hd__o221a_1
X_4313_ _4313_/A vssd1 vssd1 vccd1 vccd1 _8409_/D sky130_fd_sc_hd__clkbuf_1
X_8081_ _8625_/CLK _8081_/D vssd1 vssd1 vccd1 vccd1 _8081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5293_ _8409_/Q _8130_/Q _5361_/S vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__mux2_1
X_7032_ _7032_/A vssd1 vssd1 vccd1 vccd1 _7032_/X sky130_fd_sc_hd__buf_1
X_4244_ _4244_/A vssd1 vssd1 vccd1 vccd1 _8468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4175_ _8253_/Q vssd1 vssd1 vccd1 vccd1 _4175_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7934_ _7934_/CLK _7934_/D vssd1 vssd1 vccd1 vccd1 _7934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7865_ _8436_/CLK _7865_/D vssd1 vssd1 vccd1 vccd1 _7865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7131__523 _7132__524/A vssd1 vssd1 vccd1 vccd1 _8332_/CLK sky130_fd_sc_hd__inv_2
X_6816_ _6822_/A vssd1 vssd1 vccd1 vccd1 _6816_/X sky130_fd_sc_hd__buf_1
XFILLER_51_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7796_ _7796_/A _7812_/B vssd1 vssd1 vccd1 vccd1 _7796_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7203__80 _7203__80/A vssd1 vssd1 vccd1 vccd1 _8389_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6747_ _6747_/A vssd1 vssd1 vccd1 vccd1 _8102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3959_ _8576_/Q vssd1 vssd1 vccd1 vccd1 _3959_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3459_ clkbuf_0__3459_/X vssd1 vssd1 vccd1 vccd1 _7127__520/A sky130_fd_sc_hd__clkbuf_4
X_5629_ _5629_/A vssd1 vssd1 vccd1 vccd1 _8069_/D sky130_fd_sc_hd__clkbuf_1
X_8417_ _8417_/CLK _8417_/D vssd1 vssd1 vccd1 vccd1 _8417_/Q sky130_fd_sc_hd__dfxtp_1
X_7088__488 _7089__489/A vssd1 vssd1 vccd1 vccd1 _8297_/CLK sky130_fd_sc_hd__inv_2
X_8348_ _8348_/CLK _8348_/D vssd1 vssd1 vccd1 vccd1 _8348_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3427_ _6971_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3427_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8279_ _8279_/CLK _8279_/D vssd1 vssd1 vccd1 vccd1 _8279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7737__37 _7738__38/A vssd1 vssd1 vccd1 vccd1 _8588_/CLK sky130_fd_sc_hd__inv_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7499__166 _7503__170/A vssd1 vssd1 vccd1 vccd1 _8505_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7512__1 _7513__2/A vssd1 vssd1 vccd1 vccd1 _8515_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__or2_1
XFILLER_18_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4931_ _4917_/X _4930_/X _4989_/A vssd1 vssd1 vccd1 vccd1 _4931_/X sky130_fd_sc_hd__o21a_1
X_4862_ _4812_/A _8107_/Q _8003_/Q _4822_/A vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__a22o_1
X_7650_ _7650_/A vssd1 vssd1 vccd1 vccd1 _8553_/D sky130_fd_sc_hd__clkbuf_1
X_6601_ _6625_/A vssd1 vssd1 vccd1 vccd1 _6601_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3313_ clkbuf_0__3313_/X vssd1 vssd1 vccd1 vccd1 _6788__343/A sky130_fd_sc_hd__clkbuf_4
X_4793_ _4758_/X _4792_/X _4706_/X vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__a21o_1
X_7581_ _7581_/A _7579_/A vssd1 vssd1 vccd1 vccd1 _7581_/X sky130_fd_sc_hd__or2b_1
X_6532_ _6532_/A vssd1 vssd1 vccd1 vccd1 _7970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7443__121 _7443__121/A vssd1 vssd1 vccd1 vccd1 _8460_/CLK sky130_fd_sc_hd__inv_2
X_6463_ _7946_/Q _6410_/X _6452_/X _6462_/X _6459_/X vssd1 vssd1 vccd1 vccd1 _7946_/D
+ sky130_fd_sc_hd__a221o_1
X_5414_ _5414_/A vssd1 vssd1 vccd1 vccd1 _8184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8202_ _8202_/CLK _8202_/D vssd1 vssd1 vccd1 vccd1 _8202_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput122 _6057_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput111 _6035_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__buf_2
X_8133_ _8133_/CLK _8133_/D vssd1 vssd1 vccd1 vccd1 _8133_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput133 _6024_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__buf_2
X_6394_ _8608_/Q vssd1 vssd1 vccd1 vccd1 _6394_/Y sky130_fd_sc_hd__inv_2
Xoutput155 _5997_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput144 _5975_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput166 _5955_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__buf_2
X_5345_ _8367_/Q _8375_/Q _5345_/S vssd1 vssd1 vccd1 vccd1 _5345_/X sky130_fd_sc_hd__mux2_1
Xoutput177 _6083_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__buf_2
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8064_ _8064_/CLK _8064_/D vssd1 vssd1 vccd1 vccd1 _8064_/Q sky130_fd_sc_hd__dfxtp_1
X_5276_ _5276_/A vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__clkbuf_2
Xoutput199 _6089_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput188 _6086_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__buf_2
X_4227_ _8473_/Q _4226_/X _4230_/S vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3460_ clkbuf_0__3460_/X vssd1 vssd1 vccd1 vccd1 _7133__525/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4158_ _8257_/Q vssd1 vssd1 vccd1 vccd1 _5663_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4089_ _8507_/Q _3931_/X _4095_/S vssd1 vssd1 vccd1 vccd1 _4090_/A sky130_fd_sc_hd__mux2_1
X_6920__374 _6920__374/A vssd1 vssd1 vccd1 vccd1 _8170_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7917_ _7917_/CLK _7917_/D vssd1 vssd1 vccd1 vccd1 _7917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7848_ _7848_/CLK _7848_/D vssd1 vssd1 vccd1 vccd1 _7848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7779_ _5985_/A _7778_/X _7777_/A vssd1 vssd1 vccd1 vccd1 _7779_/X sky130_fd_sc_hd__a21bo_1
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6630__275 _6630__275/A vssd1 vssd1 vccd1 vccd1 _8035_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3658_ clkbuf_0__3658_/X vssd1 vssd1 vccd1 vccd1 _7516__5/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_4
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _6184_/A sky130_fd_sc_hd__clkbuf_4
Xinput35 caravel_wb_error_i vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _3902_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_116_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7507__173 _7509__175/A vssd1 vssd1 vccd1 vccd1 _8512_/CLK sky130_fd_sc_hd__inv_2
Xinput57 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _6030_/A sky130_fd_sc_hd__buf_4
Xinput79 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _5980_/A sky130_fd_sc_hd__buf_4
XFILLER_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5130_ _5258_/S vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__buf_2
X_5061_ _5061_/A vssd1 vssd1 vccd1 vccd1 _8223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4012_ _4012_/A vssd1 vssd1 vccd1 vccd1 _8539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5963_ _7812_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__or2_1
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4914_ _4853_/A _8041_/Q _8025_/Q _4874_/A _4860_/A vssd1 vssd1 vccd1 vccd1 _4914_/X
+ sky130_fd_sc_hd__a221o_1
X_7702_ _8568_/Q _7704_/B vssd1 vssd1 vccd1 vccd1 _7702_/X sky130_fd_sc_hd__or2_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5894_ _4209_/X _7854_/Q _5896_/S vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4845_ _4845_/A vssd1 vssd1 vccd1 vccd1 _4845_/X sky130_fd_sc_hd__clkbuf_2
X_7633_ _7633_/A vssd1 vssd1 vccd1 vccd1 _8549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4776_ _7909_/Q _8029_/Q _8045_/Q _8013_/Q _4721_/X _4694_/A vssd1 vssd1 vccd1 vccd1
+ _4777_/B sky130_fd_sc_hd__mux4_1
X_7564_ _7564_/A _7564_/B vssd1 vssd1 vccd1 vccd1 _7564_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6515_ _6023_/A _7963_/Q _6515_/S vssd1 vssd1 vccd1 vccd1 _6516_/A sky130_fd_sc_hd__mux2_1
X_6446_ _6481_/C _8249_/Q _6448_/C _7055_/B vssd1 vssd1 vccd1 vccd1 _6446_/X sky130_fd_sc_hd__a31o_1
X_6377_ _6377_/A _6381_/B vssd1 vssd1 vccd1 vccd1 _6499_/B sky130_fd_sc_hd__or2_1
X_8116_ _8116_/CLK _8116_/D vssd1 vssd1 vccd1 vccd1 _8116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5328_ _8579_/Q _5276_/A _5257_/X _8595_/Q _5120_/A vssd1 vssd1 vccd1 vccd1 _5328_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8047_ _8047_/CLK _8047_/D vssd1 vssd1 vccd1 vccd1 _8047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5259_ _8581_/Q _5103_/B _5258_/X _5232_/A vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3443_ clkbuf_0__3443_/X vssd1 vssd1 vccd1 vccd1 _7044__455/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7144__533 _7144__533/A vssd1 vssd1 vccd1 vccd1 _8342_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4453_/X _8286_/Q _4638_/S vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__mux2_1
X_6676__297 _6678__299/A vssd1 vssd1 vccd1 vccd1 _8065_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4561_ _8316_/Q _4516_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__mux2_1
X_6300_ _6300_/A vssd1 vssd1 vccd1 vccd1 _7760_/A sky130_fd_sc_hd__buf_2
X_7182__63 _7183__64/A vssd1 vssd1 vccd1 vccd1 _8372_/CLK sky130_fd_sc_hd__inv_2
X_4492_ _8574_/Q vssd1 vssd1 vccd1 vccd1 _4492_/X sky130_fd_sc_hd__buf_2
X_7280_ _8433_/Q _7282_/B _7280_/C vssd1 vssd1 vccd1 vccd1 _7379_/A sky130_fd_sc_hd__nand3_2
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6231_ _6647_/A vssd1 vssd1 vccd1 vccd1 _6423_/A sky130_fd_sc_hd__clkbuf_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7957_/Q _6195_/C _7794_/B vssd1 vssd1 vccd1 vccd1 _6176_/A sky130_fd_sc_hd__a21bo_2
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5113_ _5144_/B _5125_/B vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__or2_2
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _7864_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6093_/X sky130_fd_sc_hd__or2_1
X_5044_ _5044_/A vssd1 vssd1 vccd1 vccd1 _8230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5946_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5877_ _5877_/A vssd1 vssd1 vccd1 vccd1 _7905_/D sky130_fd_sc_hd__clkbuf_1
X_4828_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__clkbuf_2
X_7616_ _7615_/Y _7667_/B _7604_/X _7563_/B vssd1 vssd1 vccd1 vccd1 _7616_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8596_ _8596_/CLK _8596_/D vssd1 vssd1 vccd1 vccd1 _8596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4759_ _7851_/Q _7859_/Q _7934_/Q _8038_/Q _4691_/A _4725_/X vssd1 vssd1 vccd1 vccd1
+ _4759_/X sky130_fd_sc_hd__mux4_2
X_7547_ _7793_/A _6846_/B _7546_/Y vssd1 vssd1 vccd1 vccd1 _7573_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6429_ _6427_/Y _6385_/A _6428_/Y _6398_/X _6387_/A vssd1 vssd1 vccd1 vccd1 _6430_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8569_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7456__131 _7458__133/A vssd1 vssd1 vccd1 vccd1 _8470_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3426_ clkbuf_0__3426_/X vssd1 vssd1 vccd1 vccd1 _6977_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6933__384 _6934__385/A vssd1 vssd1 vccd1 vccd1 _8180_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6643__285 _6643__285/A vssd1 vssd1 vccd1 vccd1 _8045_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _7987_/Q _5607_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5801_/A sky130_fd_sc_hd__mux2_1
X_3992_ _3965_/X _8582_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _5731_/A vssd1 vssd1 vccd1 vccd1 _8018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5662_ _5662_/A vssd1 vssd1 vccd1 vccd1 _8056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8450_ _8604_/CLK _8450_/D vssd1 vssd1 vccd1 vccd1 _8450_/Q sky130_fd_sc_hd__dfxtp_1
X_8381_ _8381_/CLK _8381_/D vssd1 vssd1 vccd1 vccd1 _8381_/Q sky130_fd_sc_hd__dfxtp_1
X_5593_ _5593_/A vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__buf_2
X_4613_ _8293_/Q _4486_/X _4619_/S vssd1 vssd1 vccd1 vccd1 _4614_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3460_ _7128_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3460_/X sky130_fd_sc_hd__clkbuf_16
X_7401_ _8441_/Q _7408_/B vssd1 vssd1 vccd1 vccd1 _7401_/X sky130_fd_sc_hd__and2_1
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4544_ _4441_/X _8322_/Q _4544_/S vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__mux2_1
X_7332_ _7590_/A _7281_/X _7268_/B _8623_/Q vssd1 vssd1 vccd1 vccd1 _7332_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7263_ _7324_/A _7263_/B vssd1 vssd1 vccd1 vccd1 _7297_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ _8189_/Q vssd1 vssd1 vccd1 vccd1 _4475_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6145_ _7878_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__or2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_15 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6076_ _7936_/Q input3/X _6188_/B vssd1 vssd1 vccd1 vccd1 _6076_/X sky130_fd_sc_hd__mux2_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_37 _6160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_59 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_48 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5027_ _8237_/Q _4519_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_26 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5929_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3658_ _7511_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3658_/X sky130_fd_sc_hd__clkbuf_16
X_8579_ _8579_/CLK _8579_/D vssd1 vssd1 vccd1 vccd1 _8579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6586__239 _6587__240/A vssd1 vssd1 vccd1 vccd1 _7999_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6788__343 _6788__343/A vssd1 vssd1 vccd1 vccd1 _8135_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4260_ _4454_/A _4970_/B _4970_/C vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__or3_2
XFILLER_113_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4213_/S vssd1 vssd1 vccd1 vccd1 _4204_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7950_ _8091_/CLK _7950_/D vssd1 vssd1 vccd1 vccd1 _7950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6901_ _6901_/A _7549_/B vssd1 vssd1 vccd1 vccd1 _6902_/D sky130_fd_sc_hd__xnor2_1
X_7881_ _8091_/CLK _7881_/D vssd1 vssd1 vccd1 vccd1 _7881_/Q sky130_fd_sc_hd__dfxtp_1
X_6832_ _8556_/Q _6903_/D _8557_/Q vssd1 vssd1 vccd1 vccd1 _7588_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3975_ _3974_/X _8587_/Q _3978_/S vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__mux2_1
X_6694_ _6694_/A vssd1 vssd1 vccd1 vccd1 _6694_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3475_ clkbuf_0__3475_/X vssd1 vssd1 vccd1 vccd1 _7203__80/A sky130_fd_sc_hd__clkbuf_4
X_5714_ _5613_/X _8025_/Q _5716_/S vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__mux2_1
X_8502_ _8502_/CLK _8502_/D vssd1 vssd1 vccd1 vccd1 _8502_/Q sky130_fd_sc_hd__dfxtp_1
X_5645_ _5645_/A _5808_/A vssd1 vssd1 vccd1 vccd1 _5661_/S sky130_fd_sc_hd__or2_2
X_8433_ _8436_/CLK _8433_/D vssd1 vssd1 vccd1 vccd1 _8433_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3443_ _7039_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3443_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8364_ _8364_/CLK _8364_/D vssd1 vssd1 vccd1 vccd1 _8364_/Q sky130_fd_sc_hd__dfxtp_2
X_5576_ _5591_/S vssd1 vssd1 vccd1 vccd1 _5585_/S sky130_fd_sc_hd__buf_2
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4527_ _4527_/A vssd1 vssd1 vccd1 vccd1 _8329_/D sky130_fd_sc_hd__clkbuf_1
X_8295_ _8295_/CLK _8295_/D vssd1 vssd1 vccd1 vccd1 _8295_/Q sky130_fd_sc_hd__dfxtp_1
X_7315_ _8616_/Q _7358_/A vssd1 vssd1 vccd1 vccd1 _7412_/A sky130_fd_sc_hd__nand2_1
X_4458_ _4453_/X _8350_/Q _4470_/S vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__mux2_1
X_7246_ _8618_/Q _7246_/B vssd1 vssd1 vccd1 vccd1 _7334_/B sky130_fd_sc_hd__xor2_1
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4389_ _8375_/Q _4238_/X _4389_/S vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6128_ _6147_/A vssd1 vssd1 vccd1 vccd1 _6144_/S sky130_fd_sc_hd__clkbuf_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7501__168 _7502__169/A vssd1 vssd1 vccd1 vccd1 _8507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3260_ clkbuf_0__3260_/X vssd1 vssd1 vccd1 vccd1 _6646__287/A sky130_fd_sc_hd__clkbuf_4
X_5430_ _5430_/A vssd1 vssd1 vccd1 vccd1 _8180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5361_ _8461_/Q _8469_/Q _5361_/S vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4312_ _8409_/Q _4232_/X _4316_/S vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__mux2_1
X_5292_ _5233_/X _5290_/X _5291_/X vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__o21a_1
X_8080_ _8631_/CLK _8080_/D vssd1 vssd1 vccd1 vccd1 _8080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4243_ _8468_/Q _4215_/X _4251_/S vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _8259_/Q _8254_/Q vssd1 vssd1 vccd1 vccd1 _4666_/C sky130_fd_sc_hd__xnor2_1
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7933_ _7933_/CLK _7933_/D vssd1 vssd1 vccd1 vccd1 _7933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8652__217 vssd1 vssd1 vccd1 vccd1 _8652__217/HI core0Index[4] sky130_fd_sc_hd__conb_1
X_7864_ _8436_/CLK _7864_/D vssd1 vssd1 vccd1 vccd1 _7864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7795_ _7818_/B vssd1 vssd1 vccd1 vccd1 _7812_/B sky130_fd_sc_hd__clkbuf_2
X_6746_ _8102_/Q _6006_/A _6748_/S vssd1 vssd1 vccd1 vccd1 _6747_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3458_ clkbuf_0__3458_/X vssd1 vssd1 vccd1 vccd1 _7121__515/A sky130_fd_sc_hd__clkbuf_4
X_3958_ _3958_/A vssd1 vssd1 vccd1 vccd1 _8593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3889_ _8203_/Q _8202_/Q _8201_/Q vssd1 vssd1 vccd1 vccd1 _5370_/A sky130_fd_sc_hd__and3_1
X_5628_ _8069_/Q _5627_/X _5634_/S vssd1 vssd1 vccd1 vccd1 _5629_/A sky130_fd_sc_hd__mux2_1
X_8416_ _8452_/CLK _8416_/D vssd1 vssd1 vccd1 vccd1 _8416_/Q sky130_fd_sc_hd__dfxtp_1
X_5559_ _5398_/X _8119_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__mux2_1
X_8347_ _8347_/CLK _8347_/D vssd1 vssd1 vccd1 vccd1 _8347_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3812_ clkbuf_0__3812_/X vssd1 vssd1 vccd1 vccd1 _7751__49/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3426_ _6970_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3426_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8278_ _8278_/CLK _8278_/D vssd1 vssd1 vccd1 vccd1 _8278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7229_ _7442_/A vssd1 vssd1 vccd1 vccd1 _7229_/X sky130_fd_sc_hd__buf_1
X_7025__440 _7025__440/A vssd1 vssd1 vccd1 vccd1 _8246_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7108__504 _7109__505/A vssd1 vssd1 vccd1 vccd1 _8313_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6345__214 _6346__215/A vssd1 vssd1 vccd1 vccd1 _7926_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _4869_/X _4920_/X _4923_/X _4929_/X _4683_/A vssd1 vssd1 vccd1 vccd1 _4930_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_17_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7189__69 _7190__70/A vssd1 vssd1 vccd1 vccd1 _8378_/CLK sky130_fd_sc_hd__inv_2
X_4861_ _4861_/A vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__clkbuf_2
X_6600_ _6631_/A vssd1 vssd1 vccd1 vccd1 _6600_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3312_ clkbuf_0__3312_/X vssd1 vssd1 vccd1 vccd1 _6784__340/A sky130_fd_sc_hd__clkbuf_4
X_4792_ _8221_/Q _8108_/Q _8004_/Q _7988_/Q _4691_/A _4725_/X vssd1 vssd1 vccd1 vccd1
+ _4792_/X sky130_fd_sc_hd__mux4_1
X_7580_ _7664_/B _7573_/X _7578_/X _7664_/C vssd1 vssd1 vccd1 vccd1 _7580_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3466_ clkbuf_0__3466_/X vssd1 vssd1 vccd1 vccd1 _7164__550/A sky130_fd_sc_hd__clkbuf_16
X_6531_ _6039_/A _7970_/Q _6537_/S vssd1 vssd1 vccd1 vccd1 _6532_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6462_ _7811_/A _6471_/B _6469_/C vssd1 vssd1 vccd1 vccd1 _6462_/X sky130_fd_sc_hd__and3_1
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5413_ _5412_/X _8184_/Q _5417_/S vssd1 vssd1 vccd1 vccd1 _5414_/A sky130_fd_sc_hd__mux2_1
X_6393_ _8632_/Q _6363_/X _6373_/X vssd1 vssd1 vccd1 vccd1 _6400_/B sky130_fd_sc_hd__a21oi_1
X_8201_ _8201_/CLK _8201_/D vssd1 vssd1 vccd1 vccd1 _8201_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput123 _6059_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput112 _6037_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__buf_2
Xoutput134 _6026_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__buf_2
X_8132_ _8132_/CLK _8132_/D vssd1 vssd1 vccd1 vccd1 _8132_/Q sky130_fd_sc_hd__dfxtp_1
X_5344_ _5344_/A _5344_/B _5344_/C vssd1 vssd1 vccd1 vccd1 _5344_/X sky130_fd_sc_hd__or3_1
Xoutput145 _5977_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput156 _5999_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput167 _5957_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8063_ _8063_/CLK _8063_/D vssd1 vssd1 vccd1 vccd1 _8063_/Q sky130_fd_sc_hd__dfxtp_1
X_5275_ _8321_/Q _8337_/Q _5341_/S vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__mux2_1
Xoutput178 _6121_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput189 _6158_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_101_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4226_ _8574_/Q vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__buf_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7014_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7014_/X sky130_fd_sc_hd__buf_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4157_ _8258_/Q vssd1 vssd1 vccd1 vccd1 _4508_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4088_ _4088_/A vssd1 vssd1 vccd1 vccd1 _8508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7450__126 _7454__130/A vssd1 vssd1 vccd1 vccd1 _8465_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7916_ _7916_/CLK _7916_/D vssd1 vssd1 vccd1 vccd1 _7916_/Q sky130_fd_sc_hd__dfxtp_1
X_7094__493 _7094__493/A vssd1 vssd1 vccd1 vccd1 _8302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7847_ _7847_/CLK _7847_/D vssd1 vssd1 vccd1 vccd1 _7847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ _7778_/A vssd1 vssd1 vccd1 vccd1 _7778_/X sky130_fd_sc_hd__clkbuf_2
X_7742__41 _7743__42/A vssd1 vssd1 vccd1 vccd1 _8592_/CLK sky130_fd_sc_hd__inv_2
X_6729_ _6729_/A vssd1 vssd1 vccd1 vccd1 _8094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3657_ clkbuf_0__3657_/X vssd1 vssd1 vccd1 vccd1 _7529_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_4
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
Xinput36 wb_rst_i vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__clkbuf_4
Xinput58 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
Xinput69 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_4
Xinput47 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ _4460_/X _8223_/Q _5066_/S vssd1 vssd1 vccd1 vccd1 _5061_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4011_ _8539_/Q _3931_/X _4017_/S vssd1 vssd1 vccd1 vccd1 _4012_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5962_ _6008_/B vssd1 vssd1 vccd1 vccd1 _5971_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4913_ _8009_/Q _4716_/B _4821_/A vssd1 vssd1 vccd1 vccd1 _4913_/X sky130_fd_sc_hd__a21o_1
X_7701_ _8568_/Q _7687_/A _7700_/X _7684_/A vssd1 vssd1 vccd1 vccd1 _8567_/D sky130_fd_sc_hd__o211a_1
X_5893_ _5893_/A vssd1 vssd1 vccd1 vccd1 _7855_/D sky130_fd_sc_hd__clkbuf_1
X_4844_ _8011_/Q _4716_/B _4821_/X vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__a21o_1
X_7632_ _7630_/X _7649_/B vssd1 vssd1 vccd1 vccd1 _7633_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4775_ _4713_/X _4772_/X _4774_/X vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__a21o_1
X_7563_ _8629_/Q _7563_/B vssd1 vssd1 vccd1 vccd1 _7563_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6514_ _6514_/A vssd1 vssd1 vccd1 vccd1 _7962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6445_ _8145_/Q vssd1 vssd1 vccd1 vccd1 _6481_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6376_ _7962_/Q _6376_/B _7961_/Q vssd1 vssd1 vccd1 vccd1 _6381_/B sky130_fd_sc_hd__or3b_1
X_5327_ _8121_/Q _8148_/Q _5330_/S vssd1 vssd1 vccd1 vccd1 _5327_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8115_ _8115_/CLK _8115_/D vssd1 vssd1 vccd1 vccd1 _8115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8046_ _8046_/CLK _8046_/D vssd1 vssd1 vccd1 vccd1 _8046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5258_ _8123_/Q _8150_/Q _5258_/S vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__mux2_2
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5189_ _5189_/A _5189_/B vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__and2_1
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3442_ clkbuf_0__3442_/X vssd1 vssd1 vccd1 vccd1 _7051_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ _8189_/Q vssd1 vssd1 vccd1 vccd1 _4209_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8658__223 vssd1 vssd1 vccd1 vccd1 _8658__223/HI core1Index[3] sky130_fd_sc_hd__conb_1
XFILLER_73_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6966__397 _6968__399/A vssd1 vssd1 vccd1 vccd1 _8201_/CLK sky130_fd_sc_hd__inv_2
X_6782__338 _6782__338/A vssd1 vssd1 vccd1 vccd1 _8130_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _8317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4491_ _4491_/A vssd1 vssd1 vccd1 vccd1 _8340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6230_ _6222_/X _7893_/Q _6225_/X _6229_/X _7861_/Q vssd1 vssd1 vccd1 vccd1 _7861_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6195_/B vssd1 vssd1 vccd1 vccd1 _7794_/B sky130_fd_sc_hd__clkbuf_2
X_5112_ _5112_/A _5112_/B vssd1 vssd1 vccd1 vccd1 _5125_/B sky130_fd_sc_hd__nor2_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6149_/A vssd1 vssd1 vccd1 vccd1 _6107_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5043_ _8230_/Q _4516_/X _5047_/S vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _7000_/A vssd1 vssd1 vccd1 vccd1 _6994_/X sky130_fd_sc_hd__buf_1
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6991__413 _6991__413/A vssd1 vssd1 vccd1 vccd1 _8219_/CLK sky130_fd_sc_hd__inv_2
X_5945_ _7838_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__or2_1
Xclkbuf_0__3812_ _7747_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3812_/X sky130_fd_sc_hd__clkbuf_16
X_5876_ _7905_/Q _5613_/A _5878_/S vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4827_ _4845_/A vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__clkbuf_2
X_7615_ _8546_/Q vssd1 vssd1 vccd1 vccd1 _7615_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8595_ _8595_/CLK _8595_/D vssd1 vssd1 vccd1 vccd1 _8595_/Q sky130_fd_sc_hd__dfxtp_1
X_4758_ _4758_/A vssd1 vssd1 vccd1 vccd1 _4758_/X sky130_fd_sc_hd__clkbuf_4
X_7546_ _7588_/A _7546_/B vssd1 vssd1 vccd1 vccd1 _7546_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4689_ _4806_/B vssd1 vssd1 vccd1 vccd1 _4955_/S sky130_fd_sc_hd__buf_2
XFILLER_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6428_ _8053_/Q _6403_/A _6382_/X vssd1 vssd1 vccd1 vccd1 _6428_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _6430_/A vssd1 vssd1 vccd1 vccd1 _6359_/X sky130_fd_sc_hd__buf_2
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8029_ _8029_/CLK _8029_/D vssd1 vssd1 vccd1 vccd1 _8029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3425_ clkbuf_0__3425_/X vssd1 vssd1 vccd1 vccd1 _6968__399/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _3991_/A vssd1 vssd1 vccd1 vccd1 _8583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5730_ _8018_/Q _5636_/X _5734_/S vssd1 vssd1 vccd1 vccd1 _5731_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5661_ _5616_/X _8056_/Q _5661_/S vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__mux2_1
X_7400_ _7053_/A _7349_/B _7350_/A _7321_/Y _7399_/Y vssd1 vssd1 vccd1 vccd1 _7408_/B
+ sky130_fd_sc_hd__o221a_1
X_8380_ _8380_/CLK _8380_/D vssd1 vssd1 vccd1 vccd1 _8380_/Q sky130_fd_sc_hd__dfxtp_1
X_4612_ _4612_/A vssd1 vssd1 vccd1 vccd1 _8294_/D sky130_fd_sc_hd__clkbuf_1
X_5592_ _5592_/A vssd1 vssd1 vccd1 vccd1 _8104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4543_ _4543_/A vssd1 vssd1 vccd1 vccd1 _8323_/D sky130_fd_sc_hd__clkbuf_1
X_7331_ _7331_/A _7331_/B _7331_/C _7331_/D vssd1 vssd1 vccd1 vccd1 _7331_/X sky130_fd_sc_hd__and4_1
XFILLER_116_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7262_ _7324_/B _7324_/C vssd1 vssd1 vccd1 vccd1 _7263_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4474_ _4474_/A vssd1 vssd1 vccd1 vccd1 _8345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6144_ _7953_/Q input11/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6144_/X sky130_fd_sc_hd__mux2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_16 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6075_ _6147_/A vssd1 vssd1 vccd1 vccd1 _6188_/B sky130_fd_sc_hd__buf_4
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _8238_/D sky130_fd_sc_hd__clkbuf_1
X_6806__352 _6809__355/A vssd1 vssd1 vccd1 vccd1 _8147_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_27 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_38 _6178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_49 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6977_ _6977_/A vssd1 vssd1 vccd1 vccd1 _6977_/X sky130_fd_sc_hd__buf_1
X_5928_ _6281_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__and2_1
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5859_ _5859_/A vssd1 vssd1 vccd1 vccd1 _7913_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3657_ _7510_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3657_/X sky130_fd_sc_hd__clkbuf_16
X_8578_ _8578_/CLK _8578_/D vssd1 vssd1 vccd1 vccd1 _8578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7529_ _7529_/A vssd1 vssd1 vccd1 vccd1 _7529_/X sky130_fd_sc_hd__buf_1
XFILLER_119_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6998__419 _6999__420/A vssd1 vssd1 vccd1 vccd1 _8225_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4190_ _5645_/A _5682_/A vssd1 vssd1 vccd1 vccd1 _4213_/S sky130_fd_sc_hd__nor2_2
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7157__544 _7157__544/A vssd1 vssd1 vccd1 vccd1 _8353_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6900_ _8555_/Q _6900_/B vssd1 vssd1 vccd1 vccd1 _7549_/B sky130_fd_sc_hd__xnor2_4
X_7880_ _8091_/CLK _7880_/D vssd1 vssd1 vccd1 vccd1 _7880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6831_ _8555_/Q _6843_/A _6850_/A _6843_/C vssd1 vssd1 vccd1 vccd1 _6903_/D sky130_fd_sc_hd__and4_2
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7215__90 _7215__90/A vssd1 vssd1 vccd1 vccd1 _8399_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8501_ _8501_/CLK _8501_/D vssd1 vssd1 vccd1 vccd1 _8501_/Q sky130_fd_sc_hd__dfxtp_1
X_3974_ _8571_/Q vssd1 vssd1 vccd1 vccd1 _3974_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3474_ clkbuf_0__3474_/X vssd1 vssd1 vccd1 vccd1 _7222_/A sky130_fd_sc_hd__clkbuf_4
X_5713_ _5713_/A vssd1 vssd1 vccd1 vccd1 _8026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5644_ _5644_/A vssd1 vssd1 vccd1 vccd1 _8064_/D sky130_fd_sc_hd__clkbuf_1
X_8432_ _8440_/CLK _8432_/D vssd1 vssd1 vccd1 vccd1 _8432_/Q sky130_fd_sc_hd__dfxtp_1
X_8363_ _8363_/CLK _8363_/D vssd1 vssd1 vccd1 vccd1 _8363_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__3442_ _7038_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3442_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5575_ _5700_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5591_/S sky130_fd_sc_hd__or2_2
X_7314_ _7358_/B vssd1 vssd1 vccd1 vccd1 _7350_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8294_ _8294_/CLK _8294_/D vssd1 vssd1 vccd1 vccd1 _8294_/Q sky130_fd_sc_hd__dfxtp_1
X_4526_ _8329_/Q _4525_/X _4532_/S vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4457_ _4479_/S vssd1 vssd1 vccd1 vccd1 _4470_/S sky130_fd_sc_hd__clkbuf_4
X_7245_ _8440_/Q _7394_/A vssd1 vssd1 vccd1 vccd1 _7246_/B sky130_fd_sc_hd__xor2_1
XFILLER_112_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4388_ _4388_/A vssd1 vssd1 vccd1 vccd1 _8376_/D sky130_fd_sc_hd__clkbuf_1
X_6127_ _6117_/X _6125_/X _6126_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6127_/X sky130_fd_sc_hd__o211a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _8094_/Q _6058_/B vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__and2_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _8245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7749__47 _7752__50/A vssd1 vssd1 vccd1 vccd1 _8598_/CLK sky130_fd_sc_hd__inv_2
X_7058__464 _7058__464/A vssd1 vssd1 vccd1 vccd1 _8273_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6592__244 _6593__245/A vssd1 vssd1 vccd1 vccd1 _8004_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8638__254 vssd1 vssd1 vccd1 vccd1 partID[6] _8638__254/LO sky130_fd_sc_hd__conb_1
XFILLER_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7469__142 _7472__145/A vssd1 vssd1 vccd1 vccd1 _8481_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5360_ _8525_/Q _5276_/X _5274_/A _5358_/X _5359_/X vssd1 vssd1 vccd1 vccd1 _5360_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4311_ _4311_/A vssd1 vssd1 vccd1 vccd1 _8410_/D sky130_fd_sc_hd__clkbuf_1
X_5291_ _8495_/Q _5254_/X _5230_/B _8487_/Q _5239_/X vssd1 vssd1 vccd1 vccd1 _5291_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4242_ _4257_/S vssd1 vssd1 vccd1 vccd1 _4251_/S sky130_fd_sc_hd__buf_2
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _4454_/A _4666_/B _4666_/A _4172_/Y vssd1 vssd1 vccd1 vccd1 _4173_/X sky130_fd_sc_hd__a211o_1
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7932_ _7932_/CLK _7932_/D vssd1 vssd1 vccd1 vccd1 _7932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7863_ _8436_/CLK _7863_/D vssd1 vssd1 vccd1 vccd1 _7863_/Q sky130_fd_sc_hd__dfxtp_1
X_7794_ _8145_/Q _7794_/B _7820_/B vssd1 vssd1 vccd1 vccd1 _7818_/B sky130_fd_sc_hd__and3_1
XFILLER_51_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3957_ _3952_/X _8593_/Q _3969_/S vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__mux2_1
X_6745_ _6745_/A vssd1 vssd1 vccd1 vccd1 _8101_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3457_ clkbuf_0__3457_/X vssd1 vssd1 vccd1 vccd1 _7114__509/A sky130_fd_sc_hd__clkbuf_4
X_8415_ _8440_/CLK _8415_/D vssd1 vssd1 vccd1 vccd1 _8415_/Q sky130_fd_sc_hd__dfxtp_2
X_3888_ _3953_/A _5112_/A _3887_/Y vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__a21bo_1
X_5627_ _8193_/Q vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5558_ _5573_/S vssd1 vssd1 vccd1 vccd1 _5567_/S sky130_fd_sc_hd__clkbuf_4
X_8346_ _8346_/CLK _8346_/D vssd1 vssd1 vccd1 vccd1 _8346_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3811_ clkbuf_0__3811_/X vssd1 vssd1 vccd1 vccd1 _7746__45/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3425_ _6964_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3425_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8277_ _8277_/CLK _8277_/D vssd1 vssd1 vccd1 vccd1 _8277_/Q sky130_fd_sc_hd__dfxtp_1
X_4509_ _5862_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _4532_/S sky130_fd_sc_hd__nor2_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7228_ _7448_/A vssd1 vssd1 vccd1 vccd1 _7228_/X sky130_fd_sc_hd__buf_1
X_5489_ _8153_/Q _4486_/X _5495_/S vssd1 vssd1 vccd1 vccd1 _5490_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7159_ _7159_/A vssd1 vssd1 vccd1 vccd1 _7159_/X sky130_fd_sc_hd__buf_1
XFILLER_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_wb_clk_i _6197_/A vssd1 vssd1 vccd1 vccd1 _7972_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4860_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3311_ clkbuf_0__3311_/X vssd1 vssd1 vccd1 vccd1 _6776__333/A sky130_fd_sc_hd__clkbuf_4
X_4791_ _8176_/Q _8168_/Q _7996_/Q _8237_/Q _4710_/X _4702_/X vssd1 vssd1 vccd1 vccd1
+ _4791_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6530_ _6530_/A vssd1 vssd1 vccd1 vccd1 _7969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6461_ _8623_/Q vssd1 vssd1 vccd1 vccd1 _7811_/A sky130_fd_sc_hd__clkbuf_4
X_5412_ _5604_/A vssd1 vssd1 vccd1 vccd1 _5412_/X sky130_fd_sc_hd__buf_2
X_8200_ _8200_/CLK _8200_/D vssd1 vssd1 vccd1 vccd1 _8200_/Q sky130_fd_sc_hd__dfxtp_4
X_6392_ _7936_/Q _6359_/X _6389_/Y _6391_/X vssd1 vssd1 vccd1 vccd1 _7936_/D sky130_fd_sc_hd__a211o_1
Xoutput124 _6062_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput113 _6040_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8131_ _8131_/CLK _8131_/D vssd1 vssd1 vccd1 vccd1 _8131_/Q sky130_fd_sc_hd__dfxtp_1
X_5343_ _5274_/X _5341_/X _5342_/X _5142_/S vssd1 vssd1 vccd1 vccd1 _5344_/C sky130_fd_sc_hd__o211a_1
Xoutput135 _6029_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__buf_2
Xoutput157 _6001_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput168 _5959_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__buf_2
Xoutput146 _5979_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__buf_2
X_8062_ _8062_/CLK _8062_/D vssd1 vssd1 vccd1 vccd1 _8062_/Q sky130_fd_sc_hd__dfxtp_1
X_5274_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__clkbuf_2
Xoutput179 _6124_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__buf_2
X_4225_ _4225_/A vssd1 vssd1 vccd1 vccd1 _8474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4156_ _8195_/Q vssd1 vssd1 vccd1 vccd1 _4156_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _8508_/Q _3872_/X _4095_/S vssd1 vssd1 vccd1 vccd1 _4088_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7915_ _7915_/CLK _7915_/D vssd1 vssd1 vccd1 vccd1 _7915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7846_ _7846_/CLK _7846_/D vssd1 vssd1 vccd1 vccd1 _7846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7777_ _7777_/A vssd1 vssd1 vccd1 vccd1 _7777_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4989_ _4989_/A vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6728_ _5989_/A _8094_/Q _6730_/S vssd1 vssd1 vccd1 vccd1 _6729_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6659_ _8266_/Q _6663_/B vssd1 vssd1 vccd1 vccd1 _6660_/A sky130_fd_sc_hd__and2_1
X_8329_ _8329_/CLK _8329_/D vssd1 vssd1 vccd1 vccd1 _8329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3656_ clkbuf_0__3656_/X vssd1 vssd1 vccd1 vccd1 _7506__172/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _6186_/A sky130_fd_sc_hd__clkbuf_4
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_4
X_7194__73 _7194__73/A vssd1 vssd1 vccd1 vccd1 _8382_/CLK sky130_fd_sc_hd__inv_2
Xinput37 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _6010_/A sky130_fd_sc_hd__buf_4
XFILLER_116_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput59 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _6014_/A sky130_fd_sc_hd__buf_4
Xinput48 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _6012_/A sky130_fd_sc_hd__buf_4
XFILLER_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4010_ _4010_/A vssd1 vssd1 vccd1 vccd1 _8540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6978__406 _6982__410/A vssd1 vssd1 vccd1 vccd1 _8210_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5961_ _5961_/A vssd1 vssd1 vccd1 vccd1 _5961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7700_ _8567_/Q _7704_/B vssd1 vssd1 vccd1 vccd1 _7700_/X sky130_fd_sc_hd__or2_1
X_4912_ _4831_/X _8033_/Q _7846_/Q _4833_/X _4758_/A vssd1 vssd1 vccd1 vccd1 _4912_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5892_ _4206_/X _7855_/Q _5896_/S vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__mux2_1
X_7631_ _7683_/A vssd1 vssd1 vccd1 vccd1 _7649_/B sky130_fd_sc_hd__clkbuf_2
X_4843_ _4683_/X _4819_/X _4825_/X _4842_/X vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__o31a_1
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _4758_/X _4773_/X _4706_/X vssd1 vssd1 vccd1 vccd1 _4774_/X sky130_fd_sc_hd__a21o_1
X_7562_ _7562_/A _7562_/B _7562_/C _7562_/D vssd1 vssd1 vccd1 vccd1 _7562_/X sky130_fd_sc_hd__or4_1
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6513_ _6021_/A _7962_/Q _6515_/S vssd1 vssd1 vccd1 vccd1 _6514_/A sky130_fd_sc_hd__mux2_1
X_6444_ _6501_/A _6442_/X _6443_/X vssd1 vssd1 vccd1 vccd1 _7943_/D sky130_fd_sc_hd__a21o_1
X_6375_ _7967_/Q _6375_/B _7968_/Q _6371_/A vssd1 vssd1 vccd1 vccd1 _6377_/A sky130_fd_sc_hd__or4b_1
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8114_ _8114_/CLK _8114_/D vssd1 vssd1 vccd1 vccd1 _8114_/Q sky130_fd_sc_hd__dfxtp_1
X_5326_ _5393_/B _5324_/X _5325_/X vssd1 vssd1 vccd1 vccd1 _5326_/Y sky130_fd_sc_hd__o21ai_1
X_8045_ _8045_/CLK _8045_/D vssd1 vssd1 vccd1 vccd1 _8045_/Q sky130_fd_sc_hd__dfxtp_1
X_5257_ _5359_/B vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__clkbuf_2
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _8479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5188_ _8591_/Q _8340_/Q _8324_/Q _8364_/Q _5130_/X _5101_/A vssd1 vssd1 vccd1 vccd1
+ _5189_/B sky130_fd_sc_hd__mux4_2
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3441_ clkbuf_0__3441_/X vssd1 vssd1 vccd1 vccd1 _7034__447/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4139_ _4154_/S vssd1 vssd1 vccd1 vccd1 _4148_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7829_ _8627_/Q _7826_/X _7828_/X _6423_/X vssd1 vssd1 vccd1 vccd1 _8627_/D sky130_fd_sc_hd__a211o_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7151__539 _7152__540/A vssd1 vssd1 vccd1 vccd1 _8348_/CLK sky130_fd_sc_hd__inv_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4490_ _8340_/Q _4489_/X _4496_/S vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6160_/A _6188_/B vssd1 vssd1 vccd1 vccd1 _6160_/X sky130_fd_sc_hd__and2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5111_ _8601_/Q _8154_/Q _8127_/Q _8585_/Q _5345_/S _5110_/X vssd1 vssd1 vccd1 vccd1
+ _5111_/X sky130_fd_sc_hd__mux4_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _7939_/Q input28/X _6106_/S vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__mux2_1
X_5042_ _5042_/A vssd1 vssd1 vccd1 vccd1 _8231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3811_ _7741_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3811_/X sky130_fd_sc_hd__clkbuf_16
X_5944_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5875_ _5875_/A vssd1 vssd1 vccd1 vccd1 _7906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__clkbuf_2
X_8594_ _8594_/CLK _8594_/D vssd1 vssd1 vccd1 vccd1 _8594_/Q sky130_fd_sc_hd__dfxtp_1
X_7614_ _7614_/A vssd1 vssd1 vccd1 vccd1 _8545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7545_ _7793_/A _6846_/B _6905_/B vssd1 vssd1 vccd1 vccd1 _7573_/A sky130_fd_sc_hd__o21a_1
X_4757_ _4834_/A vssd1 vssd1 vccd1 vccd1 _4758_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4688_ _4723_/A vssd1 vssd1 vccd1 vccd1 _4994_/B sky130_fd_sc_hd__clkbuf_4
X_6427_ _8612_/Q vssd1 vssd1 vccd1 vccd1 _6427_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6358_ _6483_/A vssd1 vssd1 vccd1 vccd1 _6430_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ _5393_/B _5307_/X _5308_/X vssd1 vssd1 vccd1 vccd1 _5309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6289_ _7714_/A _7896_/Q _6291_/S vssd1 vssd1 vccd1 vccd1 _6290_/A sky130_fd_sc_hd__mux2_1
X_8028_ _8028_/CLK _8028_/D vssd1 vssd1 vccd1 vccd1 _8028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_wb_clk_i _6197_/A vssd1 vssd1 vccd1 vccd1 _8617_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7463__137 _7463__137/A vssd1 vssd1 vccd1 vccd1 _8476_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ _3962_/X _8583_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3991_/A sky130_fd_sc_hd__mux2_1
X_5660_ _5660_/A vssd1 vssd1 vccd1 vccd1 _8057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _8294_/Q _4481_/X _4619_/S vssd1 vssd1 vccd1 vccd1 _4612_/A sky130_fd_sc_hd__mux2_1
X_5591_ _5428_/X _8104_/Q _5591_/S vssd1 vssd1 vccd1 vccd1 _5592_/A sky130_fd_sc_hd__mux2_1
X_4542_ _4438_/X _8323_/Q _4544_/S vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__mux2_1
X_7330_ _7330_/A _7330_/B _7330_/C vssd1 vssd1 vccd1 vccd1 _7330_/X sky130_fd_sc_hd__and3_1
X_4473_ _4472_/X _8345_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__mux2_1
X_7261_ _8431_/Q _7274_/A _7282_/A _7282_/B _8432_/Q vssd1 vssd1 vccd1 vccd1 _7324_/C
+ sky130_fd_sc_hd__a41o_1
X_6212_ _6212_/A vssd1 vssd1 vccd1 vccd1 _6212_/X sky130_fd_sc_hd__buf_1
X_6143_ _6136_/X _6141_/X _6142_/X _6139_/X vssd1 vssd1 vccd1 vccd1 _6143_/X sky130_fd_sc_hd__o211a_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6195_/B _5918_/B _5919_/X _7844_/Q vssd1 vssd1 vccd1 vccd1 _6147_/A sky130_fd_sc_hd__a31oi_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_39 _6178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_28 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_17 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _8238_/Q _4516_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__mux2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5927_ _5927_/A vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7528__15 _7528__15/A vssd1 vssd1 vccd1 vccd1 _8529_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _4447_/X _7913_/Q _5860_/S vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__mux2_1
X_5789_ _5789_/A vssd1 vssd1 vccd1 vccd1 _7992_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3656_ _7504_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3656_/X sky130_fd_sc_hd__clkbuf_16
X_4809_ _4809_/A vssd1 vssd1 vccd1 vccd1 _4996_/B sky130_fd_sc_hd__buf_2
X_8577_ _8577_/CLK _8577_/D vssd1 vssd1 vccd1 vccd1 _8577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6830_ _8550_/Q _8549_/Q _8548_/Q _8547_/Q vssd1 vssd1 vccd1 vccd1 _6843_/C sky130_fd_sc_hd__and4_1
X_6795__349 _6796__350/A vssd1 vssd1 vccd1 vccd1 _8141_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8500_ _8500_/CLK _8500_/D vssd1 vssd1 vccd1 vccd1 _8500_/Q sky130_fd_sc_hd__dfxtp_1
X_5712_ _5610_/X _8026_/Q _5716_/S vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__mux2_1
X_3973_ _3973_/A vssd1 vssd1 vccd1 vccd1 _8588_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3473_ clkbuf_0__3473_/X vssd1 vssd1 vccd1 vccd1 _7194__73/A sky130_fd_sc_hd__clkbuf_4
X_5643_ _8064_/Q _5642_/X _5643_/S vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__mux2_1
X_8431_ _8440_/CLK _8431_/D vssd1 vssd1 vccd1 vccd1 _8431_/Q sky130_fd_sc_hd__dfxtp_1
X_5574_ _5574_/A vssd1 vssd1 vccd1 vccd1 _8112_/D sky130_fd_sc_hd__clkbuf_1
X_8362_ _8362_/CLK _8362_/D vssd1 vssd1 vccd1 vccd1 _8362_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3441_ _7032_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3441_/X sky130_fd_sc_hd__clkbuf_16
X_7313_ _7334_/B _7313_/B _7313_/C _7313_/D vssd1 vssd1 vccd1 vccd1 _7358_/B sky130_fd_sc_hd__and4_1
X_4525_ _8190_/Q vssd1 vssd1 vccd1 vccd1 _4525_/X sky130_fd_sc_hd__buf_2
X_8293_ _8293_/CLK _8293_/D vssd1 vssd1 vccd1 vccd1 _8293_/Q sky130_fd_sc_hd__dfxtp_1
X_4456_ _5645_/A _5880_/A vssd1 vssd1 vccd1 vccd1 _4479_/S sky130_fd_sc_hd__or2_2
X_7244_ _7244_/A vssd1 vssd1 vccd1 vccd1 _7394_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4387_ _8376_/Q _4235_/X _4389_/S vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6126_ _7873_/Q _6126_/B vssd1 vssd1 vccd1 vccd1 _6126_/X sky130_fd_sc_hd__or2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A vssd1 vssd1 vccd1 vccd1 _6057_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6626__271 _6626__271/A vssd1 vssd1 vccd1 vccd1 _8031_/CLK sky130_fd_sc_hd__inv_2
X_5008_ _8245_/Q _4519_/X _5010_/S vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__mux2_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0__3809_ clkbuf_0__3809_/X vssd1 vssd1 vccd1 vccd1 _7732__33/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6959_ _6959_/A vssd1 vssd1 vccd1 vccd1 _8195_/D sky130_fd_sc_hd__clkbuf_1
X_8629_ _8633_/CLK _8629_/D vssd1 vssd1 vccd1 vccd1 _8629_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4310_ _8410_/Q _4229_/X _4310_/S vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5290_ _8463_/Q _8471_/Q _5352_/S vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__mux2_1
X_4241_ _5539_/B _4241_/B vssd1 vssd1 vccd1 vccd1 _4257_/S sky130_fd_sc_hd__nor2_2
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4172_ _4172_/A vssd1 vssd1 vccd1 vccd1 _4172_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7931_ _7931_/CLK _7931_/D vssd1 vssd1 vccd1 vccd1 _7931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _8436_/CLK _7862_/D vssd1 vssd1 vccd1 vccd1 _7862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7793_ _7793_/A _7811_/B vssd1 vssd1 vccd1 vccd1 _7793_/Y sky130_fd_sc_hd__nand2_1
X_6209__183 _6209__183/A vssd1 vssd1 vccd1 vccd1 _7852_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6744_ _8101_/Q _6004_/A _6748_/S vssd1 vssd1 vccd1 vccd1 _6745_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _3978_/S vssd1 vssd1 vccd1 vccd1 _3969_/S sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3456_ clkbuf_0__3456_/X vssd1 vssd1 vccd1 vccd1 _7105__501/A sky130_fd_sc_hd__clkbuf_4
X_5626_ _5626_/A vssd1 vssd1 vccd1 vccd1 _8070_/D sky130_fd_sc_hd__clkbuf_1
X_8414_ _8414_/CLK _8414_/D vssd1 vssd1 vccd1 vccd1 _8414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ _8205_/Q _8200_/Q vssd1 vssd1 vccd1 vccd1 _3887_/Y sky130_fd_sc_hd__xnor2_1
X_8345_ _8345_/CLK _8345_/D vssd1 vssd1 vccd1 vccd1 _8345_/Q sky130_fd_sc_hd__dfxtp_1
X_5557_ _5700_/A _5718_/B vssd1 vssd1 vccd1 vccd1 _5573_/S sky130_fd_sc_hd__or2_2
Xclkbuf_1_0_0__3810_ clkbuf_0__3810_/X vssd1 vssd1 vccd1 vccd1 _7738__38/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5488_ _5488_/A vssd1 vssd1 vccd1 vccd1 _8154_/D sky130_fd_sc_hd__clkbuf_1
X_8276_ _8276_/CLK _8276_/D vssd1 vssd1 vccd1 vccd1 _8276_/Q sky130_fd_sc_hd__dfxtp_1
X_4508_ _5663_/A _4508_/B _5663_/B vssd1 vssd1 vccd1 vccd1 _5718_/B sky130_fd_sc_hd__or3_4
X_4439_ _4438_/X _8355_/Q _4442_/S vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6147_/A vssd1 vssd1 vccd1 vccd1 _6125_/S sky130_fd_sc_hd__buf_2
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6819__363 _6819__363/A vssd1 vssd1 vccd1 vccd1 _8158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4790_ _4713_/X _4787_/X _4789_/X vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6460_ _7945_/Q _6410_/X _6452_/X _6457_/X _6459_/X vssd1 vssd1 vccd1 vccd1 _7945_/D
+ sky130_fd_sc_hd__a221o_1
X_5411_ _8192_/Q vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__clkbuf_2
X_6391_ _7806_/A vssd1 vssd1 vccd1 vccd1 _6391_/X sky130_fd_sc_hd__clkbuf_4
Xoutput125 _6064_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput114 _6042_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__buf_2
X_8130_ _8130_/CLK _8130_/D vssd1 vssd1 vccd1 vccd1 _8130_/Q sky130_fd_sc_hd__dfxtp_1
X_5342_ _8359_/Q _5276_/X _5249_/A _8586_/Q vssd1 vssd1 vccd1 vccd1 _5342_/X sky130_fd_sc_hd__o22a_1
Xoutput158 _6003_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput136 _6031_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__buf_2
Xoutput147 _5981_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__buf_2
X_7009__426 _7009__426/A vssd1 vssd1 vccd1 vccd1 _8232_/CLK sky130_fd_sc_hd__inv_2
X_8061_ _8061_/CLK _8061_/D vssd1 vssd1 vccd1 vccd1 _8061_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput169 _5961_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_102_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5273_ _5269_/X _5270_/X _5272_/X vssd1 vssd1 vccd1 vccd1 _5279_/B sky130_fd_sc_hd__o21a_1
X_4224_ _8474_/Q _4223_/X _4230_/S vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4155_ _4155_/A vssd1 vssd1 vccd1 vccd1 _8485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4086_ _4101_/S vssd1 vssd1 vccd1 vccd1 _4095_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7914_ _7914_/CLK _7914_/D vssd1 vssd1 vccd1 vccd1 _7914_/Q sky130_fd_sc_hd__dfxtp_1
X_7845_ _7845_/CLK _7845_/D vssd1 vssd1 vccd1 vccd1 _7845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7776_ _7776_/A vssd1 vssd1 vccd1 vccd1 _7777_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4988_ _4988_/A vssd1 vssd1 vccd1 vccd1 _4988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3939_ _3939_/A vssd1 vssd1 vccd1 vccd1 _8598_/D sky130_fd_sc_hd__clkbuf_1
X_6727_ _6727_/A vssd1 vssd1 vccd1 vccd1 _8093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3439_ clkbuf_0__3439_/X vssd1 vssd1 vccd1 vccd1 _7025__440/A sky130_fd_sc_hd__clkbuf_4
X_6658_ _6658_/A vssd1 vssd1 vccd1 vccd1 _8052_/D sky130_fd_sc_hd__clkbuf_1
X_5609_ _5609_/A vssd1 vssd1 vccd1 vccd1 _8075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8328_ _8328_/CLK _8328_/D vssd1 vssd1 vccd1 vccd1 _8328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8259_ _8259_/CLK _8259_/D vssd1 vssd1 vccd1 vccd1 _8259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3655_ clkbuf_0__3655_/X vssd1 vssd1 vccd1 vccd1 _7503__170/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6752__314 _6753__315/A vssd1 vssd1 vccd1 vccd1 _8106_/CLK sky130_fd_sc_hd__inv_2
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__clkbuf_4
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _6160_/A sky130_fd_sc_hd__clkbuf_4
X_6639__281 _6641__283/A vssd1 vssd1 vccd1 vccd1 _8041_/CLK sky130_fd_sc_hd__inv_2
Xinput49 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _3902_/D sky130_fd_sc_hd__clkbuf_1
Xinput38 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _6032_/A sky130_fd_sc_hd__buf_4
XFILLER_115_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5960_ _7815_/A _5960_/B vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__or2_1
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5891_ _5891_/A vssd1 vssd1 vccd1 vccd1 _7856_/D sky130_fd_sc_hd__clkbuf_1
X_4911_ _4853_/X _7929_/Q _7854_/Q _4829_/X _4809_/A vssd1 vssd1 vccd1 vccd1 _4911_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7630_ _6861_/A _7620_/X _7625_/X _6864_/B vssd1 vssd1 vccd1 vccd1 _7630_/X sky130_fd_sc_hd__o22a_1
X_4842_ _4737_/X _4836_/X _4840_/X _4992_/B _4673_/A vssd1 vssd1 vccd1 vccd1 _4842_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4773_ _8222_/Q _8109_/Q _8005_/Q _7989_/Q _4691_/A _4725_/X vssd1 vssd1 vccd1 vccd1
+ _4773_/X sky130_fd_sc_hd__mux4_1
X_7561_ _7834_/A _7611_/A _7611_/B vssd1 vssd1 vccd1 vccd1 _7562_/D sky130_fd_sc_hd__and3b_1
X_7492_ _7498_/A vssd1 vssd1 vccd1 vccd1 _7492_/X sky130_fd_sc_hd__buf_1
X_6512_ _6512_/A vssd1 vssd1 vccd1 vccd1 _7961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6443_ _7943_/Q _6430_/A _7806_/A vssd1 vssd1 vccd1 vccd1 _6443_/X sky130_fd_sc_hd__a21o_1
X_6374_ _8633_/Q _6363_/X _6373_/X vssd1 vssd1 vccd1 vccd1 _6389_/B sky130_fd_sc_hd__a21oi_1
X_8113_ _8113_/CLK _8113_/D vssd1 vssd1 vccd1 vccd1 _8113_/Q sky130_fd_sc_hd__dfxtp_1
X_5325_ _8494_/Q _5236_/X _5249_/X _8486_/Q _5135_/X vssd1 vssd1 vccd1 vccd1 _5325_/X
+ sky130_fd_sc_hd__o221a_1
X_8044_ _8044_/CLK _8044_/D vssd1 vssd1 vccd1 vccd1 _8044_/Q sky130_fd_sc_hd__dfxtp_1
X_5256_ _5233_/X _5253_/X _5255_/X vssd1 vssd1 vccd1 vccd1 _5256_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3440_ clkbuf_0__3440_/X vssd1 vssd1 vccd1 vccd1 _7031__445/A sky130_fd_sc_hd__clkbuf_4
X_4207_ _8479_/Q _4206_/X _4213_/S vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5187_ _5185_/X _5186_/X _5246_/S vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4138_ _5826_/A _4241_/B vssd1 vssd1 vccd1 vccd1 _4154_/S sky130_fd_sc_hd__nor2_2
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4069_ _4069_/A vssd1 vssd1 vccd1 vccd1 _8516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7828_ _7828_/A _7842_/B _7840_/C vssd1 vssd1 vccd1 vccd1 _7828_/X sky130_fd_sc_hd__and3_1
X_7759_ _7759_/A vssd1 vssd1 vccd1 vccd1 _8606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5110_ _5123_/A vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6147_/A vssd1 vssd1 vccd1 vccd1 _6106_/S sky130_fd_sc_hd__buf_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5041_ _8231_/Q _4513_/X _5047_/S vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3810_ _7735_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3810_/X sky130_fd_sc_hd__clkbuf_16
X_5943_ _7840_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5944_/A sky130_fd_sc_hd__or2_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6620__266 _6621__267/A vssd1 vssd1 vccd1 vccd1 _8026_/CLK sky130_fd_sc_hd__inv_2
X_5874_ _7906_/Q _5610_/A _5878_/S vssd1 vssd1 vccd1 vccd1 _5875_/A sky130_fd_sc_hd__mux2_1
X_4825_ _8330_/Q _4817_/X _4994_/B _4824_/X vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__o211a_1
X_8593_ _8593_/CLK _8593_/D vssd1 vssd1 vccd1 vccd1 _8593_/Q sky130_fd_sc_hd__dfxtp_1
X_7613_ _7612_/X _7628_/B vssd1 vssd1 vccd1 vccd1 _7614_/A sky130_fd_sc_hd__and2b_1
X_6323__196 _6325__198/A vssd1 vssd1 vccd1 vccd1 _7908_/CLK sky130_fd_sc_hd__inv_2
X_7544_ _7581_/A vssd1 vssd1 vccd1 vccd1 _7664_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _4754_/X _4755_/X _4756_/S vssd1 vssd1 vccd1 vccd1 _4756_/X sky130_fd_sc_hd__mux2_1
X_4687_ _4687_/A vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6426_ _7564_/A _6403_/X _6387_/X vssd1 vssd1 vccd1 vccd1 _6430_/B sky130_fd_sc_hd__a21oi_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6357_ _6454_/A _6368_/A vssd1 vssd1 vccd1 vccd1 _6483_/A sky130_fd_sc_hd__nor2b_2
XFILLER_68_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5308_ _8304_/Q _5236_/X _5249_/X _8288_/Q _5095_/A vssd1 vssd1 vccd1 vccd1 _5308_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6288_ _6288_/A vssd1 vssd1 vccd1 vccd1 _7895_/D sky130_fd_sc_hd__clkbuf_1
X_8027_ _8027_/CLK _8027_/D vssd1 vssd1 vccd1 vccd1 _8027_/Q sky130_fd_sc_hd__dfxtp_1
X_5239_ _5239_/A vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4610_ _4625_/S vssd1 vssd1 vccd1 vccd1 _4619_/S sky130_fd_sc_hd__buf_2
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5590_ _5590_/A vssd1 vssd1 vccd1 vccd1 _8105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4541_ _4541_/A vssd1 vssd1 vccd1 vccd1 _8324_/D sky130_fd_sc_hd__clkbuf_1
X_8648__213 vssd1 vssd1 vccd1 vccd1 _8648__213/HI core0Index[0] sky130_fd_sc_hd__conb_1
X_6203__178 _6204__179/A vssd1 vssd1 vccd1 vccd1 _7847_/CLK sky130_fd_sc_hd__inv_2
X_7127__520 _7127__520/A vssd1 vssd1 vccd1 vccd1 _8329_/CLK sky130_fd_sc_hd__inv_2
X_7260_ _7260_/A vssd1 vssd1 vccd1 vccd1 _7282_/B sky130_fd_sc_hd__clkbuf_2
X_4472_ _8190_/Q vssd1 vssd1 vccd1 vccd1 _4472_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7191_ _7191_/A vssd1 vssd1 vccd1 vccd1 _7191_/X sky130_fd_sc_hd__buf_1
X_6142_ _7877_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6142_/X sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6073_ _6136_/A vssd1 vssd1 vccd1 vccd1 _6073_/X sky130_fd_sc_hd__clkbuf_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_29 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5024_ _5024_/A vssd1 vssd1 vccd1 vccd1 _8239_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_18 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7232__103 _7234__105/A vssd1 vssd1 vccd1 vccd1 _8412_/CLK sky130_fd_sc_hd__inv_2
X_5926_ _6303_/C _5930_/B vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__and2_1
XFILLER_110_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5857_ _5857_/A vssd1 vssd1 vccd1 vccd1 _7914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3655_ _7498_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3655_/X sky130_fd_sc_hd__clkbuf_16
X_5788_ _7992_/Q _5616_/A _5788_/S vssd1 vssd1 vccd1 vccd1 _5789_/A sky130_fd_sc_hd__mux2_1
X_4808_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__clkbuf_2
X_8576_ _8612_/CLK _8576_/D vssd1 vssd1 vccd1 vccd1 _8576_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6813__358 _6813__358/A vssd1 vssd1 vccd1 vccd1 _8153_/CLK sky130_fd_sc_hd__inv_2
X_4739_ _4683_/X _4708_/X _4720_/X _4738_/X vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__a31o_2
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6409_ _7938_/Q _6359_/X _6408_/Y _6391_/X vssd1 vssd1 vccd1 vccd1 _7938_/D sky130_fd_sc_hd__a211o_1
X_7389_ _7398_/A _7389_/B vssd1 vssd1 vccd1 vccd1 _8436_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7515__4 _7516__5/A vssd1 vssd1 vccd1 vccd1 _8518_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ _6760_/A vssd1 vssd1 vccd1 vccd1 _6760_/X sky130_fd_sc_hd__buf_1
XFILLER_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3472_ clkbuf_0__3472_/X vssd1 vssd1 vccd1 vccd1 _7190__70/A sky130_fd_sc_hd__clkbuf_4
X_5711_ _5711_/A vssd1 vssd1 vccd1 vccd1 _8027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3972_ _3971_/X _8588_/Q _3978_/S vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__mux2_1
X_5642_ _8188_/Q vssd1 vssd1 vccd1 vccd1 _5642_/X sky130_fd_sc_hd__clkbuf_2
X_8430_ _8452_/CLK _8430_/D vssd1 vssd1 vccd1 vccd1 _8430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5573_ _5428_/X _8112_/Q _5573_/S vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3440_ _7026_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3440_/X sky130_fd_sc_hd__clkbuf_16
X_8361_ _8361_/CLK _8361_/D vssd1 vssd1 vccd1 vccd1 _8361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4524_ _4524_/A vssd1 vssd1 vccd1 vccd1 _8330_/D sky130_fd_sc_hd__clkbuf_1
X_7312_ _7299_/Y _7300_/X _7304_/Y _7307_/Y _7327_/B vssd1 vssd1 vccd1 vccd1 _7313_/D
+ sky130_fd_sc_hd__o2111a_1
X_8292_ _8292_/CLK _8292_/D vssd1 vssd1 vccd1 vccd1 _8292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7243_ _8439_/Q _8438_/Q _7306_/B vssd1 vssd1 vccd1 vccd1 _7244_/A sky130_fd_sc_hd__nand3_1
X_4455_ _4979_/A _4985_/A _4970_/C vssd1 vssd1 vccd1 vccd1 _5880_/A sky130_fd_sc_hd__or3_4
X_4386_ _4386_/A vssd1 vssd1 vccd1 vccd1 _8377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6125_ _7948_/Q input6/X _6125_/S vssd1 vssd1 vccd1 vccd1 _6125_/X sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _8093_/Q _6058_/B vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__and2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _8246_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6958_ _8569_/Q _6958_/B vssd1 vssd1 vccd1 vccd1 _6959_/A sky130_fd_sc_hd__and2_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5909_ _5909_/A vssd1 vssd1 vccd1 vccd1 _7848_/D sky130_fd_sc_hd__clkbuf_1
X_6889_ _8551_/Q vssd1 vssd1 vccd1 vccd1 _6891_/A sky130_fd_sc_hd__inv_2
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7221__95 _7221__95/A vssd1 vssd1 vccd1 vccd1 _8404_/CLK sky130_fd_sc_hd__inv_2
X_8628_ _8633_/CLK _8628_/D vssd1 vssd1 vccd1 vccd1 _8628_/Q sky130_fd_sc_hd__dfxtp_1
X_8559_ _8561_/CLK _8559_/D vssd1 vssd1 vccd1 vccd1 _8559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6633__276 _6636__279/A vssd1 vssd1 vccd1 vccd1 _8036_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4240_ _4240_/A vssd1 vssd1 vccd1 vccd1 _8469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7476__148 _7477__149/A vssd1 vssd1 vccd1 vccd1 _8487_/CLK sky130_fd_sc_hd__inv_2
X_4171_ _4259_/A _4171_/B vssd1 vssd1 vccd1 vccd1 _4666_/A sky130_fd_sc_hd__nand2_1
X_7930_ _7930_/CLK _7930_/D vssd1 vssd1 vccd1 vccd1 _7930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _8436_/CLK _7861_/D vssd1 vssd1 vccd1 vccd1 _7861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7792_ _7817_/B vssd1 vssd1 vccd1 vccd1 _7811_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6743_ _6743_/A vssd1 vssd1 vccd1 vccd1 _8100_/D sky130_fd_sc_hd__clkbuf_1
X_3955_ _4355_/A _4534_/A vssd1 vssd1 vccd1 vccd1 _3978_/S sky130_fd_sc_hd__or2_2
X_6674_ _6674_/A vssd1 vssd1 vccd1 vccd1 _6674_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3455_ clkbuf_0__3455_/X vssd1 vssd1 vccd1 vccd1 _7128_/A sky130_fd_sc_hd__clkbuf_4
X_5625_ _8070_/Q _5624_/X _5634_/S vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__mux2_1
X_8413_ _8413_/CLK _8413_/D vssd1 vssd1 vccd1 vccd1 _8413_/Q sky130_fd_sc_hd__dfxtp_1
X_3886_ _8199_/Q vssd1 vssd1 vccd1 vccd1 _5112_/A sky130_fd_sc_hd__clkbuf_2
X_5556_ _5556_/A vssd1 vssd1 vccd1 vccd1 _8120_/D sky130_fd_sc_hd__clkbuf_1
X_8344_ _8344_/CLK _8344_/D vssd1 vssd1 vccd1 vccd1 _8344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5487_ _8154_/Q _4481_/X _5495_/S vssd1 vssd1 vccd1 vccd1 _5488_/A sky130_fd_sc_hd__mux2_1
X_4507_ _8195_/Q vssd1 vssd1 vccd1 vccd1 _4507_/X sky130_fd_sc_hd__buf_2
X_8275_ _8275_/CLK _8275_/D vssd1 vssd1 vccd1 vccd1 _8275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4438_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4369_ _4131_/X _8384_/Q _4371_/S vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6098_/X _6106_/X _6107_/X _6101_/X vssd1 vssd1 vccd1 vccd1 _6108_/X sky130_fd_sc_hd__o211a_1
X_6039_ _6039_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6040_/A sky130_fd_sc_hd__and2_1
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6575__230 _6575__230/A vssd1 vssd1 vccd1 vccd1 _7990_/CLK sky130_fd_sc_hd__inv_2
X_7482__152 _7483__153/A vssd1 vssd1 vccd1 vccd1 _8491_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5410_ _5410_/A vssd1 vssd1 vccd1 vccd1 _8185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6390_ _6390_/A vssd1 vssd1 vccd1 vccd1 _7806_/A sky130_fd_sc_hd__clkbuf_2
Xoutput115 _6044_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__buf_2
X_5341_ _8319_/Q _8335_/Q _5341_/S vssd1 vssd1 vccd1 vccd1 _5341_/X sky130_fd_sc_hd__mux2_1
Xoutput126 _6066_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput148 _5983_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput137 _5930_/B vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__buf_2
Xoutput159 _6005_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__buf_2
X_8060_ _8060_/CLK _8060_/D vssd1 vssd1 vccd1 vccd1 _8060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5272_ _8305_/Q _5271_/X _5257_/X _8289_/Q _5135_/A vssd1 vssd1 vccd1 vccd1 _5272_/X
+ sky130_fd_sc_hd__o221a_1
X_4223_ _8575_/Q vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__buf_2
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4154_ _8485_/Q _3949_/X _4154_/S vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4085_ _5826_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _4101_/S sky130_fd_sc_hd__nor2_2
XFILLER_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7913_ _7913_/CLK _7913_/D vssd1 vssd1 vccd1 vccd1 _7913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7844_ _8617_/CLK _7844_/D vssd1 vssd1 vccd1 vccd1 _7844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7775_ _8146_/Q _7820_/B vssd1 vssd1 vccd1 vccd1 _7776_/A sky130_fd_sc_hd__and2_1
XFILLER_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6726_ _5987_/A _8093_/Q _6730_/S vssd1 vssd1 vccd1 vccd1 _6727_/A sky130_fd_sc_hd__mux2_1
X_4987_ _4987_/A vssd1 vssd1 vccd1 vccd1 _8255_/D sky130_fd_sc_hd__clkbuf_1
X_3938_ _8598_/Q _3937_/X _3941_/S vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3438_ clkbuf_0__3438_/X vssd1 vssd1 vccd1 vccd1 _7017__433/A sky130_fd_sc_hd__clkbuf_4
X_6657_ _8265_/Q _6663_/B vssd1 vssd1 vccd1 vccd1 _6658_/A sky130_fd_sc_hd__and2_1
X_6588_ _6594_/A vssd1 vssd1 vccd1 vccd1 _6588_/X sky130_fd_sc_hd__buf_1
X_5608_ _5607_/X _8075_/Q _5608_/S vssd1 vssd1 vccd1 vccd1 _5609_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5539_ _5539_/A _5539_/B vssd1 vssd1 vccd1 vccd1 _5555_/S sky130_fd_sc_hd__nor2_2
X_8327_ _8327_/CLK _8327_/D vssd1 vssd1 vccd1 vccd1 _8327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8258_ _8258_/CLK _8258_/D vssd1 vssd1 vccd1 vccd1 _8258_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3654_ clkbuf_0__3654_/X vssd1 vssd1 vccd1 vccd1 _7496__164/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8553_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_8189_ _8568_/CLK _8189_/D vssd1 vssd1 vccd1 vccd1 _8189_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3019_ clkbuf_0__3019_/X vssd1 vssd1 vccd1 vccd1 _6217__190/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput39 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _6034_/A sky130_fd_sc_hd__buf_4
X_8681__246 vssd1 vssd1 vccd1 vccd1 _8681__246/HI versionID[0] sky130_fd_sc_hd__conb_1
XFILLER_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7121__515 _7121__515/A vssd1 vssd1 vccd1 vccd1 _8324_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _4203_/X _7856_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__mux2_1
X_4910_ _8328_/Q _4817_/X _4723_/A _4909_/X vssd1 vssd1 vccd1 vccd1 _4910_/X sky130_fd_sc_hd__o211a_1
X_4841_ _4841_/A vssd1 vssd1 vccd1 vccd1 _4992_/B sky130_fd_sc_hd__buf_2
X_7015__431 _7017__433/A vssd1 vssd1 vccd1 vccd1 _8237_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4772_ _8177_/Q _8169_/Q _7997_/Q _8238_/Q _4710_/X _4702_/X vssd1 vssd1 vccd1 vccd1
+ _4772_/X sky130_fd_sc_hd__mux4_1
X_7560_ _8631_/Q _7608_/B vssd1 vssd1 vccd1 vccd1 _7562_/C sky130_fd_sc_hd__xor2_1
XFILLER_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6511_ _6019_/A _7961_/Q _6515_/S vssd1 vssd1 vccd1 vccd1 _6512_/A sky130_fd_sc_hd__mux2_1
X_6442_ _7821_/A _6363_/X _6452_/A _6436_/Y _6441_/X vssd1 vssd1 vccd1 vccd1 _6442_/X
+ sky130_fd_sc_hd__a32o_1
X_8112_ _8112_/CLK _8112_/D vssd1 vssd1 vccd1 vccd1 _8112_/Q sky130_fd_sc_hd__dfxtp_1
X_6373_ _6387_/A vssd1 vssd1 vccd1 vccd1 _6373_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5324_ _8462_/Q _8470_/Q _5324_/S vssd1 vssd1 vccd1 vccd1 _5324_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8043_ _8043_/CLK _8043_/D vssd1 vssd1 vccd1 vccd1 _8043_/Q sky130_fd_sc_hd__dfxtp_1
X_5255_ _8496_/Q _5254_/X _5230_/B _8488_/Q _5239_/X vssd1 vssd1 vccd1 vccd1 _5255_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4206_ _8190_/Q vssd1 vssd1 vccd1 vccd1 _4206_/X sky130_fd_sc_hd__clkbuf_4
X_5186_ _8388_/Q _8380_/Q _8372_/Q _8396_/Q _5138_/X _5131_/X vssd1 vssd1 vccd1 vccd1
+ _5186_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4137_ _4137_/A vssd1 vssd1 vccd1 vccd1 _8493_/D sky130_fd_sc_hd__clkbuf_1
X_4068_ _8516_/Q _3872_/X _4076_/S vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7489__158 _7491__160/A vssd1 vssd1 vccd1 vccd1 _8497_/CLK sky130_fd_sc_hd__inv_2
X_7827_ _7842_/C vssd1 vssd1 vccd1 vccd1 _7840_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7758_ _8206_/Q _7836_/A vssd1 vssd1 vccd1 vccd1 _7759_/A sky130_fd_sc_hd__and2_1
X_6709_ _6709_/A vssd1 vssd1 vccd1 vccd1 _8085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7689_ _7704_/B vssd1 vssd1 vccd1 vccd1 _7698_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5040_ _5040_/A vssd1 vssd1 vccd1 vccd1 _8232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5942_ _5942_/A vssd1 vssd1 vccd1 vccd1 _7840_/A sky130_fd_sc_hd__buf_6
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5873_ _5873_/A vssd1 vssd1 vccd1 vccd1 _7907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824_ _8019_/Q _4821_/X _4823_/X _4996_/B vssd1 vssd1 vccd1 vccd1 _4824_/X sky130_fd_sc_hd__o22a_1
X_8592_ _8592_/CLK _8592_/D vssd1 vssd1 vccd1 vccd1 _8592_/Q sky130_fd_sc_hd__dfxtp_1
X_7612_ _7610_/Y _7667_/B _7604_/X _7611_/Y vssd1 vssd1 vccd1 vccd1 _7612_/X sky130_fd_sc_hd__o22a_1
X_4755_ _8231_/Q _8186_/Q _8078_/Q _8423_/Q _4710_/A _4729_/X vssd1 vssd1 vccd1 vccd1
+ _4755_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4686_ _4733_/A vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__clkbuf_2
X_6425_ _8628_/Q vssd1 vssd1 vccd1 vccd1 _7564_/A sky130_fd_sc_hd__buf_4
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5307_ _8534_/Q _8272_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__mux2_1
X_8026_ _8026_/CLK _8026_/D vssd1 vssd1 vccd1 vccd1 _8026_/Q sky130_fd_sc_hd__dfxtp_1
X_6287_ _7838_/A _7895_/Q _6291_/S vssd1 vssd1 vccd1 vccd1 _6288_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5238_ _5238_/A vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__buf_2
X_5169_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__buf_2
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8441_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4540_ _4435_/X _8324_/Q _4544_/S vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4471_ _4471_/A vssd1 vssd1 vccd1 vccd1 _8346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6141_ _7952_/Q input10/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6141_/X sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6765__325 _6765__325/A vssd1 vssd1 vccd1 vccd1 _8117_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6136_/A sky130_fd_sc_hd__clkbuf_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _8239_/Q _4513_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _5024_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_19 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5856_ _4444_/X _7914_/Q _5860_/S vssd1 vssd1 vccd1 vccd1 _5857_/A sky130_fd_sc_hd__mux2_1
X_4807_ _4807_/A _4856_/A vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__nand2_2
Xclkbuf_0__3654_ _7492_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3654_/X sky130_fd_sc_hd__clkbuf_16
X_5787_ _5787_/A vssd1 vssd1 vccd1 vccd1 _7993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8575_ _8612_/CLK _8575_/D vssd1 vssd1 vccd1 vccd1 _8575_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4738_ _4723_/X _4728_/X _4734_/X _4735_/X _4737_/X vssd1 vssd1 vccd1 vccd1 _4738_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4669_ _4669_/A vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6408_ _6416_/A _6408_/B _6408_/C vssd1 vssd1 vccd1 vccd1 _6408_/Y sky130_fd_sc_hd__nor3_2
X_7388_ _8436_/Q _7384_/X _7376_/X _7311_/B vssd1 vssd1 vccd1 vccd1 _7389_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6666__289 _6667__290/A vssd1 vssd1 vccd1 vccd1 _8057_/CLK sky130_fd_sc_hd__inv_2
X_8009_ _8009_/CLK _8009_/D vssd1 vssd1 vccd1 vccd1 _8009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3019_ _6212_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3019_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ _8572_/Q vssd1 vssd1 vccd1 vccd1 _3971_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3471_ clkbuf_0__3471_/X vssd1 vssd1 vccd1 vccd1 _7183__64/A sky130_fd_sc_hd__clkbuf_4
X_5710_ _5607_/X _8027_/Q _5710_/S vssd1 vssd1 vccd1 vccd1 _5711_/A sky130_fd_sc_hd__mux2_1
X_5641_ _5641_/A vssd1 vssd1 vccd1 vccd1 _8065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5572_ _5572_/A vssd1 vssd1 vccd1 vccd1 _8113_/D sky130_fd_sc_hd__clkbuf_1
X_8360_ _8360_/CLK _8360_/D vssd1 vssd1 vccd1 vccd1 _8360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8291_ _8291_/CLK _8291_/D vssd1 vssd1 vccd1 vccd1 _8291_/Q sky130_fd_sc_hd__dfxtp_1
X_4523_ _8330_/Q _4522_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__mux2_1
X_7311_ _7808_/A _7311_/B vssd1 vssd1 vccd1 vccd1 _7327_/B sky130_fd_sc_hd__xor2_1
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7242_ _8437_/Q _7260_/A _7280_/C _7308_/C vssd1 vssd1 vccd1 vccd1 _7306_/B sky130_fd_sc_hd__and4_2
X_4454_ _4454_/A vssd1 vssd1 vccd1 vccd1 _4979_/A sky130_fd_sc_hd__inv_2
X_4385_ _8377_/Q _4232_/X _4389_/S vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__mux2_1
X_7173_ _7173_/A vssd1 vssd1 vccd1 vccd1 _7173_/X sky130_fd_sc_hd__buf_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6124_ _6117_/X _6122_/X _6123_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6124_/X sky130_fd_sc_hd__o211a_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _8246_/Q _4516_/X _5010_/S vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__mux2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7206__82 _7208__84/A vssd1 vssd1 vccd1 vccd1 _8391_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6957_ _6957_/A vssd1 vssd1 vccd1 vccd1 _8194_/D sky130_fd_sc_hd__clkbuf_1
X_5908_ _4203_/X _7848_/Q _5908_/S vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__mux2_1
X_6888_ _7554_/B _7554_/C vssd1 vssd1 vccd1 vccd1 _7590_/B sky130_fd_sc_hd__nand2_2
XFILLER_22_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5839_ _5839_/A vssd1 vssd1 vccd1 vccd1 _7922_/D sky130_fd_sc_hd__clkbuf_1
X_8627_ _8633_/CLK _8627_/D vssd1 vssd1 vccd1 vccd1 _8627_/Q sky130_fd_sc_hd__dfxtp_2
X_8558_ _8561_/CLK _8558_/D vssd1 vssd1 vccd1 vccd1 _8558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8489_ _8489_/CLK _8489_/D vssd1 vssd1 vccd1 vccd1 _8489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7002__422 _7002__422/A vssd1 vssd1 vccd1 vccd1 _8228_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _8257_/Q _8252_/Q vssd1 vssd1 vccd1 vccd1 _4666_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _7860_/CLK _7860_/D vssd1 vssd1 vccd1 vccd1 _7860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7791_ _7791_/A _7791_/B vssd1 vssd1 vccd1 vccd1 _7817_/B sky130_fd_sc_hd__or2_1
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6742_ _8100_/Q _6002_/A _6742_/S vssd1 vssd1 vccd1 vccd1 _6743_/A sky130_fd_sc_hd__mux2_1
X_3954_ _4336_/A _5373_/A _4027_/B vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__or3_2
Xclkbuf_1_1_0__3454_ clkbuf_0__3454_/X vssd1 vssd1 vccd1 vccd1 _7102__500/A sky130_fd_sc_hd__clkbuf_4
X_3885_ _8204_/Q vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__inv_2
X_8412_ _8412_/CLK _8412_/D vssd1 vssd1 vccd1 vccd1 _8412_/Q sky130_fd_sc_hd__dfxtp_1
X_5624_ _8194_/Q vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__buf_2
X_8343_ _8343_/CLK _8343_/D vssd1 vssd1 vccd1 vccd1 _8343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5555_ _8120_/Q _4450_/A _5555_/S vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5486_ _5501_/S vssd1 vssd1 vccd1 vccd1 _5495_/S sky130_fd_sc_hd__clkbuf_2
X_4506_ _4506_/A vssd1 vssd1 vccd1 vccd1 _8335_/D sky130_fd_sc_hd__clkbuf_1
X_8274_ _8274_/CLK _8274_/D vssd1 vssd1 vccd1 vccd1 _8274_/Q sky130_fd_sc_hd__dfxtp_1
X_4437_ _4437_/A vssd1 vssd1 vccd1 vccd1 _8356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6216__189 _6216__189/A vssd1 vssd1 vccd1 vccd1 _7858_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4368_ _4368_/A vssd1 vssd1 vccd1 vccd1 _8385_/D sky130_fd_sc_hd__clkbuf_1
X_6107_ _7868_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6107_/X sky130_fd_sc_hd__or2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4299_/A _4336_/B _5376_/A vssd1 vssd1 vccd1 vccd1 _5826_/B sky130_fd_sc_hd__nand3_4
X_6038_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6778__335 _6778__335/A vssd1 vssd1 vccd1 vccd1 _8127_/CLK sky130_fd_sc_hd__inv_2
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7989_ _7989_/CLK _7989_/D vssd1 vssd1 vccd1 vccd1 _7989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7071__475 _7071__475/A vssd1 vssd1 vccd1 vccd1 _8284_/CLK sky130_fd_sc_hd__inv_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7200__77 _7200__77/A vssd1 vssd1 vccd1 vccd1 _8386_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput116 _6046_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__buf_2
X_5340_ _5269_/X _5338_/X _5339_/X vssd1 vssd1 vccd1 vccd1 _5344_/B sky130_fd_sc_hd__o21a_1
Xoutput127 _6068_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput149 _5944_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput138 _5941_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__buf_2
X_5271_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__buf_2
X_4222_ _4222_/A vssd1 vssd1 vccd1 vccd1 _8475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4153_ _4153_/A vssd1 vssd1 vccd1 vccd1 _8486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4084_ _4299_/A _4336_/B _5376_/A vssd1 vssd1 vccd1 vccd1 _5503_/B sky130_fd_sc_hd__or3_4
X_7912_ _7912_/CLK _7912_/D vssd1 vssd1 vccd1 vccd1 _7912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7843_ _8633_/Q _7826_/X _7842_/X _6269_/X vssd1 vssd1 vccd1 vccd1 _8633_/D sky130_fd_sc_hd__a211o_1
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7774_ _7790_/B _7774_/B _7774_/C vssd1 vssd1 vccd1 vccd1 _7820_/B sky130_fd_sc_hd__nor3_2
X_4986_ _7053_/C _4986_/B _4986_/C vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__and3_1
X_3937_ _8574_/Q vssd1 vssd1 vccd1 vccd1 _3937_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6725_ _6725_/A vssd1 vssd1 vccd1 vccd1 _8092_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3437_ clkbuf_0__3437_/X vssd1 vssd1 vccd1 vccd1 _7009__426/A sky130_fd_sc_hd__clkbuf_4
X_6656_ _6656_/A vssd1 vssd1 vccd1 vccd1 _8051_/D sky130_fd_sc_hd__clkbuf_1
X_5607_ _5607_/A vssd1 vssd1 vccd1 vccd1 _5607_/X sky130_fd_sc_hd__clkbuf_2
X_5538_ _5538_/A vssd1 vssd1 vccd1 vccd1 _8128_/D sky130_fd_sc_hd__clkbuf_1
X_8326_ _8326_/CLK _8326_/D vssd1 vssd1 vccd1 vccd1 _8326_/Q sky130_fd_sc_hd__dfxtp_1
X_8257_ _8257_/CLK _8257_/D vssd1 vssd1 vccd1 vccd1 _8257_/Q sky130_fd_sc_hd__dfxtp_1
X_5469_ _4427_/X _8162_/Q _5477_/S vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3653_ clkbuf_0__3653_/X vssd1 vssd1 vccd1 vccd1 _7488__157/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8188_ _8568_/CLK _8188_/D vssd1 vssd1 vccd1 vccd1 _8188_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0_0__3584_ clkbuf_0__3584_/X vssd1 vssd1 vccd1 vccd1 _7435__115/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6936__386 _6937__387/A vssd1 vssd1 vccd1 vccd1 _8182_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _6168_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3018_ clkbuf_0__3018_/X vssd1 vssd1 vccd1 vccd1 _6211__185/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7733__34 _7734__35/A vssd1 vssd1 vccd1 vccd1 _8585_/CLK sky130_fd_sc_hd__inv_2
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6646__287 _6646__287/A vssd1 vssd1 vccd1 vccd1 _8047_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4840_ _4996_/B _4837_/X _4839_/X vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4771_ _4994_/B _4768_/X _4770_/X vssd1 vssd1 vccd1 vccd1 _4771_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6510_ _6510_/A vssd1 vssd1 vccd1 vccd1 _7960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6441_ _8055_/Q _6395_/X _7055_/B vssd1 vssd1 vccd1 vccd1 _6441_/X sky130_fd_sc_hd__a21o_1
X_6372_ _6433_/A _6433_/B vssd1 vssd1 vccd1 vccd1 _6387_/A sky130_fd_sc_hd__or2_1
X_8111_ _8111_/CLK _8111_/D vssd1 vssd1 vccd1 vccd1 _8111_/Q sky130_fd_sc_hd__dfxtp_1
X_5323_ _5393_/B _5321_/X _5322_/X vssd1 vssd1 vccd1 vccd1 _5323_/Y sky130_fd_sc_hd__o21ai_1
X_8042_ _8042_/CLK _8042_/D vssd1 vssd1 vccd1 vccd1 _8042_/Q sky130_fd_sc_hd__dfxtp_1
X_5254_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5254_/X sky130_fd_sc_hd__clkbuf_2
X_5185_ _8506_/Q _8404_/Q _8141_/Q _8356_/Q _5169_/A _5140_/X vssd1 vssd1 vccd1 vccd1
+ _5185_/X sky130_fd_sc_hd__mux4_2
X_4205_ _4205_/A vssd1 vssd1 vccd1 vccd1 _8480_/D sky130_fd_sc_hd__clkbuf_1
X_4136_ _4135_/X _8493_/Q _4136_/S vssd1 vssd1 vccd1 vccd1 _4137_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4082_/S vssd1 vssd1 vccd1 vccd1 _4076_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _7826_/A vssd1 vssd1 vccd1 vccd1 _7826_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ _5055_/B _4969_/B _4985_/B vssd1 vssd1 vccd1 vccd1 _4976_/B sky130_fd_sc_hd__nand3_1
X_7757_ _7757_/A _7757_/B vssd1 vssd1 vccd1 vccd1 _8605_/D sky130_fd_sc_hd__nor2_1
X_6708_ _7803_/A _8085_/Q _6712_/S vssd1 vssd1 vccd1 vccd1 _6709_/A sky130_fd_sc_hd__mux2_1
X_7688_ _7688_/A _7688_/B vssd1 vssd1 vccd1 vccd1 _7704_/B sky130_fd_sc_hd__and2_1
XFILLER_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8309_ _8309_/CLK _8309_/D vssd1 vssd1 vccd1 vccd1 _8309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7084__485 _7084__485/A vssd1 vssd1 vccd1 vccd1 _8294_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5941_ _5941_/A vssd1 vssd1 vccd1 vccd1 _5941_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5872_ _7907_/Q _5607_/A _5872_/S vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8440_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4823_ _4812_/X _8115_/Q _8067_/Q _4822_/X vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__a22o_1
X_7611_ _7611_/A _7611_/B vssd1 vssd1 vccd1 vccd1 _7611_/Y sky130_fd_sc_hd__nand2_1
X_8591_ _8591_/CLK _8591_/D vssd1 vssd1 vccd1 vccd1 _8591_/Q sky130_fd_sc_hd__dfxtp_1
X_4754_ _8333_/Q _8118_/Q _8070_/Q _8022_/Q _4710_/A _4729_/X vssd1 vssd1 vccd1 vccd1
+ _4754_/X sky130_fd_sc_hd__mux4_1
X_7542_ _7735_/A vssd1 vssd1 vccd1 vccd1 _7542_/X sky130_fd_sc_hd__buf_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7473_ _7473_/A vssd1 vssd1 vccd1 vccd1 _7473_/X sky130_fd_sc_hd__buf_1
X_4685_ _4820_/A _4704_/A vssd1 vssd1 vccd1 vccd1 _4733_/A sky130_fd_sc_hd__or2_1
X_6424_ _7940_/Q _6410_/X _6422_/Y _6423_/X vssd1 vssd1 vccd1 vccd1 _7940_/D sky130_fd_sc_hd__a211o_1
X_5306_ _5355_/S vssd1 vssd1 vccd1 vccd1 _5321_/S sky130_fd_sc_hd__buf_2
X_6286_ _6286_/A vssd1 vssd1 vccd1 vccd1 _7894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8025_ _8025_/CLK _8025_/D vssd1 vssd1 vccd1 vccd1 _8025_/Q sky130_fd_sc_hd__dfxtp_1
X_7495__163 _7496__164/A vssd1 vssd1 vccd1 vccd1 _8502_/CLK sky130_fd_sc_hd__inv_2
X_5237_ _5237_/A vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _5283_/S vssd1 vssd1 vccd1 vccd1 _5341_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4119_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4119_/X sky130_fd_sc_hd__clkbuf_2
X_5099_ _5221_/A vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _7809_/A _7812_/B vssd1 vssd1 vccd1 vccd1 _7809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _4469_/X _8346_/Q _4470_/S vssd1 vssd1 vccd1 vccd1 _4471_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6140_ _6136_/X _6137_/X _6138_/X _6139_/X vssd1 vssd1 vccd1 vccd1 _6140_/X sky130_fd_sc_hd__o211a_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6071_ _6077_/A vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__inv_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5022_ _5022_/A vssd1 vssd1 vccd1 vccd1 _8240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5924_ _6505_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__and2_1
X_5855_ _5855_/A vssd1 vssd1 vccd1 vccd1 _7915_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3653_ _7486_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3653_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _8251_/Q _4806_/B vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__or2_2
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5786_ _7993_/Q _5613_/A _5788_/S vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__mux2_1
X_8574_ _8612_/CLK _8574_/D vssd1 vssd1 vccd1 vccd1 _8574_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_119_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3584_ _7344_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3584_/X sky130_fd_sc_hd__clkbuf_16
X_4737_ _4763_/A vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__clkbuf_4
X_4668_ _8269_/Q _6647_/B vssd1 vssd1 vccd1 vccd1 _4669_/A sky130_fd_sc_hd__nand2_1
X_6407_ _6405_/Y _6385_/X _6406_/Y _6398_/X _6387_/X vssd1 vssd1 vccd1 vccd1 _6408_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7028__442 _7028__442/A vssd1 vssd1 vccd1 vccd1 _8248_/CLK sky130_fd_sc_hd__inv_2
X_7503__170 _7503__170/A vssd1 vssd1 vccd1 vccd1 _8509_/CLK sky130_fd_sc_hd__inv_2
X_4599_ _4466_/X _8299_/Q _4601_/S vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__mux2_1
X_7387_ _7387_/A vssd1 vssd1 vccd1 vccd1 _7398_/A sky130_fd_sc_hd__buf_2
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6269_ _6390_/A vssd1 vssd1 vccd1 vccd1 _6269_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8008_ _8008_/CLK _8008_/D vssd1 vssd1 vccd1 vccd1 _8008_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3018_ _6206_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3018_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6603__252 _6603__252/A vssd1 vssd1 vccd1 vccd1 _8012_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6684__302 _6685__303/A vssd1 vssd1 vccd1 vccd1 _8070_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6348__216 _6351__219/A vssd1 vssd1 vccd1 vccd1 _7928_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3970_ _3970_/A vssd1 vssd1 vccd1 vccd1 _8589_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3470_ clkbuf_0__3470_/X vssd1 vssd1 vccd1 vccd1 _7178__60/A sky130_fd_sc_hd__clkbuf_4
X_7446__124 _7447__125/A vssd1 vssd1 vccd1 vccd1 _8463_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5640_ _8065_/Q _5639_/X _5643_/S vssd1 vssd1 vccd1 vccd1 _5641_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5571_ _5424_/X _8113_/Q _5573_/S vssd1 vssd1 vccd1 vccd1 _5572_/A sky130_fd_sc_hd__mux2_1
X_8290_ _8290_/CLK _8290_/D vssd1 vssd1 vccd1 vccd1 _8290_/Q sky130_fd_sc_hd__dfxtp_1
X_4522_ _8191_/Q vssd1 vssd1 vccd1 vccd1 _4522_/X sky130_fd_sc_hd__buf_2
X_7310_ _7310_/A _7310_/B vssd1 vssd1 vccd1 vccd1 _7311_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7241_ _8436_/Q _8435_/Q _8434_/Q _8433_/Q vssd1 vssd1 vccd1 vccd1 _7308_/C sky130_fd_sc_hd__and4_1
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4453_ _8195_/Q vssd1 vssd1 vccd1 vccd1 _4453_/X sky130_fd_sc_hd__clkbuf_4
X_4384_ _4384_/A vssd1 vssd1 vccd1 vccd1 _8378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7140__530 _7140__530/A vssd1 vssd1 vccd1 vccd1 _8339_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6123_ _7872_/Q _6126_/B vssd1 vssd1 vccd1 vccd1 _6123_/X sky130_fd_sc_hd__or2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _8092_/Q _6058_/B vssd1 vssd1 vccd1 vccd1 _6055_/A sky130_fd_sc_hd__and2_1
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A vssd1 vssd1 vccd1 vccd1 _8247_/D sky130_fd_sc_hd__clkbuf_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6956_ _8568_/Q _6958_/B vssd1 vssd1 vccd1 vccd1 _6957_/A sky130_fd_sc_hd__and2_1
X_5907_ _5907_/A vssd1 vssd1 vccd1 vccd1 _7849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6887_ _8551_/Q _6842_/C _6843_/C _8552_/Q vssd1 vssd1 vccd1 vccd1 _7554_/C sky130_fd_sc_hd__a31o_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _7922_/Q _4444_/A _5842_/S vssd1 vssd1 vccd1 vccd1 _5839_/A sky130_fd_sc_hd__mux2_1
X_8626_ _8631_/CLK _8626_/D vssd1 vssd1 vccd1 vccd1 _8626_/Q sky130_fd_sc_hd__dfxtp_2
X_5769_ _5769_/A vssd1 vssd1 vccd1 vccd1 _8001_/D sky130_fd_sc_hd__clkbuf_1
X_8557_ _8561_/CLK _8557_/D vssd1 vssd1 vccd1 vccd1 _8557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6672__294 _6672__294/A vssd1 vssd1 vccd1 vccd1 _8062_/CLK sky130_fd_sc_hd__inv_2
X_8488_ _8488_/CLK _8488_/D vssd1 vssd1 vccd1 vccd1 _8488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3249_ clkbuf_0__3249_/X vssd1 vssd1 vccd1 vccd1 _6591__243/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6810_ _6822_/A vssd1 vssd1 vccd1 vccd1 _6810_/X sky130_fd_sc_hd__buf_1
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7790_ _7790_/A _7790_/B _7790_/C _7790_/D vssd1 vssd1 vccd1 vccd1 _7791_/B sky130_fd_sc_hd__or4_1
X_6741_ _6741_/A vssd1 vssd1 vccd1 vccd1 _8099_/D sky130_fd_sc_hd__clkbuf_1
X_3953_ _3953_/A vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0__3453_ clkbuf_0__3453_/X vssd1 vssd1 vccd1 vccd1 _7094__493/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3884_ _5074_/C _5074_/D _5074_/B vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__mux2_1
X_5623_ _5623_/A vssd1 vssd1 vccd1 vccd1 _8071_/D sky130_fd_sc_hd__clkbuf_1
X_8411_ _8411_/CLK _8411_/D vssd1 vssd1 vccd1 vccd1 _8411_/Q sky130_fd_sc_hd__dfxtp_1
X_8342_ _8342_/CLK _8342_/D vssd1 vssd1 vccd1 vccd1 _8342_/Q sky130_fd_sc_hd__dfxtp_1
X_5554_ _5554_/A vssd1 vssd1 vccd1 vccd1 _8121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5485_ _5539_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _5501_/S sky130_fd_sc_hd__nor2_2
X_4505_ _8335_/Q _4504_/X _4505_/S vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__mux2_1
X_8273_ _8273_/CLK _8273_/D vssd1 vssd1 vccd1 vccd1 _8273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4436_ _4435_/X _8356_/Q _4442_/S vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4367_ _4127_/X _8385_/Q _4371_/S vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _7943_/Q input32/X _6106_/S vssd1 vssd1 vccd1 vccd1 _6106_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4298_ _4298_/A vssd1 vssd1 vccd1 vccd1 _8417_/D sky130_fd_sc_hd__clkbuf_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ _6037_/A vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ _7988_/CLK _7988_/D vssd1 vssd1 vccd1 vccd1 _7988_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8609_ _8612_/CLK _8609_/D vssd1 vssd1 vccd1 vccd1 _8609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput128 _6070_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput117 _6048_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__buf_2
Xoutput139 _5964_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__buf_2
X_5270_ _8535_/Q _8273_/Q _5355_/S vssd1 vssd1 vccd1 vccd1 _5270_/X sky130_fd_sc_hd__mux2_1
X_4221_ _8475_/Q _4220_/X _4230_/S vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4152_ _8486_/Q _3946_/X _4154_/S vssd1 vssd1 vccd1 vccd1 _4153_/A sky130_fd_sc_hd__mux2_1
X_4083_ _4083_/A vssd1 vssd1 vccd1 vccd1 _8509_/D sky130_fd_sc_hd__clkbuf_1
X_7911_ _7911_/CLK _7911_/D vssd1 vssd1 vccd1 vccd1 _7911_/Q sky130_fd_sc_hd__dfxtp_1
X_7842_ _7842_/A _7842_/B _7842_/C vssd1 vssd1 vccd1 vccd1 _7842_/X sky130_fd_sc_hd__and3_1
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7773_ _7790_/A _7790_/D _6448_/C vssd1 vssd1 vccd1 vccd1 _7774_/C sky130_fd_sc_hd__o21a_1
X_4985_ _4985_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4986_/C sky130_fd_sc_hd__or2_1
X_3936_ _3936_/A vssd1 vssd1 vccd1 vccd1 _8599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6724_ _5985_/A _8092_/Q _6724_/S vssd1 vssd1 vccd1 vccd1 _6725_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3436_ clkbuf_0__3436_/X vssd1 vssd1 vccd1 vccd1 _7020_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6655_ _8264_/Q _8249_/D vssd1 vssd1 vccd1 vccd1 _6656_/A sky130_fd_sc_hd__and2_1
X_5606_ _5606_/A vssd1 vssd1 vccd1 vccd1 _8076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5537_ _8128_/Q _4450_/A _5537_/S vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__mux2_1
X_8325_ _8325_/CLK _8325_/D vssd1 vssd1 vccd1 vccd1 _8325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8256_ _8256_/CLK _8256_/D vssd1 vssd1 vccd1 vccd1 _8256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459__134 _7460__135/A vssd1 vssd1 vccd1 vccd1 _8473_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5468_ _5483_/S vssd1 vssd1 vccd1 vccd1 _5477_/S sky130_fd_sc_hd__clkbuf_4
X_8187_ _8187_/CLK _8187_/D vssd1 vssd1 vccd1 vccd1 _8187_/Q sky130_fd_sc_hd__dfxtp_1
X_6784__340 _6784__340/A vssd1 vssd1 vccd1 vccd1 _8132_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3652_ clkbuf_0__3652_/X vssd1 vssd1 vccd1 vccd1 _7485__155/A sky130_fd_sc_hd__clkbuf_4
X_4419_ _4123_/X _8362_/Q _4419_/S vssd1 vssd1 vccd1 vccd1 _4420_/A sky130_fd_sc_hd__mux2_1
X_5399_ _5594_/A _5880_/A vssd1 vssd1 vccd1 vccd1 _5429_/S sky130_fd_sc_hd__or2_2
XFILLER_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3583_ clkbuf_0__3583_/X vssd1 vssd1 vccd1 vccd1 _7342__109/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8633_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3017_ clkbuf_0__3017_/X vssd1 vssd1 vccd1 vccd1 _6204__179/A sky130_fd_sc_hd__clkbuf_4
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _4758_/X _4769_/X _4946_/A vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6440_ _8626_/Q vssd1 vssd1 vccd1 vccd1 _7821_/A sky130_fd_sc_hd__clkbuf_4
X_6371_ _6371_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6433_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8110_ _8110_/CLK _8110_/D vssd1 vssd1 vccd1 vccd1 _8110_/Q sky130_fd_sc_hd__dfxtp_1
X_5322_ _8526_/Q _5220_/X _5249_/X _8518_/Q _5209_/A vssd1 vssd1 vccd1 vccd1 _5322_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5253_ _8464_/Q _8472_/Q _5352_/S vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__mux2_1
X_8041_ _8041_/CLK _8041_/D vssd1 vssd1 vccd1 vccd1 _8041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5184_ _5095_/A _5181_/X _5183_/X vssd1 vssd1 vccd1 vccd1 _5184_/X sky130_fd_sc_hd__a21o_1
X_4204_ _8480_/Q _4203_/X _4204_/S vssd1 vssd1 vccd1 vccd1 _4205_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4135_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4135_/X sky130_fd_sc_hd__buf_2
X_7022__437 _7023__438/A vssd1 vssd1 vccd1 vccd1 _8243_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4066_ _5844_/B _5485_/B vssd1 vssd1 vccd1 vccd1 _4082_/S sky130_fd_sc_hd__nor2_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7825_ _7825_/A vssd1 vssd1 vccd1 vccd1 _8626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8634__250 vssd1 vssd1 vccd1 vccd1 core1Index[0] _8634__250/LO sky130_fd_sc_hd__conb_1
X_4968_ _8258_/Q vssd1 vssd1 vccd1 vccd1 _5055_/B sky130_fd_sc_hd__clkbuf_4
X_7756_ _7757_/A _7756_/B vssd1 vssd1 vccd1 vccd1 _8604_/D sky130_fd_sc_hd__nor2_1
X_4899_ _4894_/X _4895_/X _4727_/X _4898_/X vssd1 vssd1 vccd1 vccd1 _4899_/X sky130_fd_sc_hd__a211o_1
X_6707_ _6707_/A vssd1 vssd1 vccd1 vccd1 _8084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7687_ _7687_/A vssd1 vssd1 vccd1 vccd1 _7687_/X sky130_fd_sc_hd__clkbuf_2
X_3919_ _7973_/Q _7974_/Q _7975_/Q _7976_/Q vssd1 vssd1 vccd1 vccd1 _6366_/B sky130_fd_sc_hd__or4_2
X_6638_ _6674_/A vssd1 vssd1 vccd1 vccd1 _6638_/X sky130_fd_sc_hd__buf_1
XFILLER_22_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8308_ _8308_/CLK _8308_/D vssd1 vssd1 vccd1 vccd1 _8308_/Q sky130_fd_sc_hd__dfxtp_1
X_6569_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6569_/X sky130_fd_sc_hd__buf_1
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8239_ _8239_/CLK _8239_/D vssd1 vssd1 vccd1 vccd1 _8239_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3249_ _6588_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3249_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6942__391 _6942__391/A vssd1 vssd1 vccd1 vccd1 _8187_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7518__6 _7519__7/A vssd1 vssd1 vccd1 vccd1 _8520_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7440__119 _7441__120/A vssd1 vssd1 vccd1 vccd1 _8458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _7842_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__or2_1
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5871_ _5871_/A vssd1 vssd1 vccd1 vccd1 _7908_/D sky130_fd_sc_hd__clkbuf_1
X_7610_ _7610_/A vssd1 vssd1 vccd1 vccd1 _7610_/Y sky130_fd_sc_hd__inv_2
X_4822_ _4822_/A vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8590_ _8590_/CLK _8590_/D vssd1 vssd1 vccd1 vccd1 _8590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _4699_/X _4750_/X _4752_/X vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__a21o_1
X_7541_ _7541_/A vssd1 vssd1 vccd1 vccd1 _7541_/X sky130_fd_sc_hd__buf_1
X_4684_ _4684_/A _4684_/B vssd1 vssd1 vccd1 vccd1 _4820_/A sky130_fd_sc_hd__and2_1
X_6423_ _6423_/A vssd1 vssd1 vccd1 vccd1 _6423_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5305_ _5305_/A vssd1 vssd1 vccd1 vccd1 _5393_/B sky130_fd_sc_hd__clkbuf_2
X_6285_ _7840_/A _7894_/Q _6291_/S vssd1 vssd1 vccd1 vccd1 _6286_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8024_ _8024_/CLK _8024_/D vssd1 vssd1 vccd1 vccd1 _8024_/Q sky130_fd_sc_hd__dfxtp_1
X_5236_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__buf_2
X_5167_ _5189_/A _5167_/B vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__and2_1
XFILLER_110_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4118_ _8574_/Q vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__buf_2
X_5098_ _5330_/S vssd1 vssd1 vccd1 vccd1 _5324_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4049_ _4049_/A vssd1 vssd1 vccd1 vccd1 _8524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8671__236 vssd1 vssd1 vccd1 vccd1 _8671__236/HI manufacturerID[8] sky130_fd_sc_hd__conb_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7808_ _7808_/A _7811_/B vssd1 vssd1 vccd1 vccd1 _7808_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6595__246 _6596__247/A vssd1 vssd1 vccd1 vccd1 _8006_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7090__490 _7090__490/A vssd1 vssd1 vccd1 vccd1 _8299_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5021_ _8240_/Q _4507_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _5022_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7218__92 _7219__93/A vssd1 vssd1 vccd1 vccd1 _8401_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5923_ _6060_/A vssd1 vssd1 vccd1 vccd1 _5930_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5854_ _4441_/X _7915_/Q _5854_/S vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3652_ _7480_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3652_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8573_ _8612_/CLK _8573_/D vssd1 vssd1 vccd1 vccd1 _8573_/Q sky130_fd_sc_hd__dfxtp_2
X_4805_ _4466_/X _4669_/X _4804_/X _4744_/X vssd1 vssd1 vccd1 vccd1 _8265_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5785_ _5785_/A vssd1 vssd1 vccd1 vccd1 _7994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3583_ _7338_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3583_/X sky130_fd_sc_hd__clkbuf_16
X_4736_ _8254_/Q _4736_/B vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7455_ _7473_/A vssd1 vssd1 vccd1 vccd1 _7455_/X sky130_fd_sc_hd__buf_1
X_4667_ _4985_/A _4665_/X _4172_/Y _4666_/X vssd1 vssd1 vccd1 vccd1 _6647_/B sky130_fd_sc_hd__o211a_2
X_7386_ _7386_/A _7386_/B vssd1 vssd1 vccd1 vccd1 _8435_/D sky130_fd_sc_hd__nor2_1
X_6406_ _8050_/Q _6395_/X _6382_/X vssd1 vssd1 vccd1 vccd1 _6406_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4598_ _4598_/A vssd1 vssd1 vccd1 vccd1 _8300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6268_ _6265_/X _8095_/Q _6261_/X _6263_/X _7884_/Q vssd1 vssd1 vccd1 vccd1 _7884_/D
+ sky130_fd_sc_hd__o32a_1
X_8007_ _8007_/CLK _8007_/D vssd1 vssd1 vccd1 vccd1 _8007_/Q sky130_fd_sc_hd__dfxtp_1
X_6199_ _6631_/A vssd1 vssd1 vccd1 vccd1 _6199_/X sky130_fd_sc_hd__buf_1
X_5219_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5276_/A sky130_fd_sc_hd__inv_2
Xclkbuf_0__3017_ _6200_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3017_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5570_ _5570_/A vssd1 vssd1 vccd1 vccd1 _8114_/D sky130_fd_sc_hd__clkbuf_1
X_4521_ _4521_/A vssd1 vssd1 vccd1 vccd1 _8331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4452_ _4452_/A vssd1 vssd1 vccd1 vccd1 _8351_/D sky130_fd_sc_hd__clkbuf_1
X_7240_ _8432_/Q _8431_/Q _8430_/Q _8429_/Q vssd1 vssd1 vccd1 vccd1 _7280_/C sky130_fd_sc_hd__and4_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4383_ _8378_/Q _4229_/X _4383_/S vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6122_ _7947_/Q input5/X _6125_/S vssd1 vssd1 vccd1 vccd1 _6122_/X sky130_fd_sc_hd__mux2_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7453__129 _7453__129/A vssd1 vssd1 vccd1 vccd1 _8468_/CLK sky130_fd_sc_hd__inv_2
X_5004_ _8247_/Q _4513_/X _5010_/S vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__mux2_1
X_6962__394 _6963__395/A vssd1 vssd1 vccd1 vccd1 _8198_/CLK sky130_fd_sc_hd__inv_2
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6955_ _6955_/A vssd1 vssd1 vccd1 vccd1 _8193_/D sky130_fd_sc_hd__clkbuf_1
X_5906_ _4200_/X _7849_/Q _5908_/S vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__mux2_1
X_8625_ _8625_/CLK _8625_/D vssd1 vssd1 vccd1 vccd1 _8625_/Q sky130_fd_sc_hd__dfxtp_2
X_6886_ _6886_/A _6886_/B _6886_/C vssd1 vssd1 vccd1 vccd1 _7554_/B sky130_fd_sc_hd__nand3_1
XFILLER_14_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5837_ _5837_/A vssd1 vssd1 vccd1 vccd1 _7923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5768_ _8001_/Q _5639_/X _5770_/S vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__mux2_1
X_7524__11 _7526__13/A vssd1 vssd1 vccd1 vccd1 _8525_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8556_ _8556_/CLK _8556_/D vssd1 vssd1 vccd1 vccd1 _8556_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4719_ _4713_/X _4715_/X _4946_/A vssd1 vssd1 vccd1 vccd1 _4719_/X sky130_fd_sc_hd__a21o_1
X_8487_ _8487_/CLK _8487_/D vssd1 vssd1 vccd1 vccd1 _8487_/Q sky130_fd_sc_hd__dfxtp_1
X_5699_ _5699_/A vssd1 vssd1 vccd1 vccd1 _8032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7369_ _7369_/A _7369_/B vssd1 vssd1 vccd1 vccd1 _7369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8677__242 vssd1 vssd1 vccd1 vccd1 _8677__242/HI partID[7] sky130_fd_sc_hd__conb_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7117__511 _7119__513/A vssd1 vssd1 vccd1 vccd1 _8320_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3248_ clkbuf_0__3248_/X vssd1 vssd1 vccd1 vccd1 _6587__240/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7212__87 _7214__89/A vssd1 vssd1 vccd1 vccd1 _8396_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6354__221 _6356__223/A vssd1 vssd1 vccd1 vccd1 _7933_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6740_ _8099_/Q _6000_/A _6742_/S vssd1 vssd1 vccd1 vccd1 _6741_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3952_ _8577_/Q vssd1 vssd1 vccd1 vccd1 _3952_/X sky130_fd_sc_hd__buf_2
XFILLER_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3452_ clkbuf_0__3452_/X vssd1 vssd1 vccd1 vccd1 _7090__490/A sky130_fd_sc_hd__clkbuf_4
X_3883_ _8202_/Q _8197_/Q vssd1 vssd1 vccd1 vccd1 _5074_/B sky130_fd_sc_hd__xnor2_1
X_5622_ _8071_/Q _5619_/X _5634_/S vssd1 vssd1 vccd1 vccd1 _5623_/A sky130_fd_sc_hd__mux2_1
X_8410_ _8410_/CLK _8410_/D vssd1 vssd1 vccd1 vccd1 _8410_/Q sky130_fd_sc_hd__dfxtp_1
X_5553_ _8121_/Q _4447_/A _5555_/S vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__mux2_1
X_8341_ _8341_/CLK _8341_/D vssd1 vssd1 vccd1 vccd1 _8341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4504_ _8570_/Q vssd1 vssd1 vccd1 vccd1 _4504_/X sky130_fd_sc_hd__clkbuf_4
X_5484_ _5484_/A vssd1 vssd1 vccd1 vccd1 _8155_/D sky130_fd_sc_hd__clkbuf_1
X_8272_ _8272_/CLK _8272_/D vssd1 vssd1 vccd1 vccd1 _8272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4435_ _4435_/A vssd1 vssd1 vccd1 vccd1 _4435_/X sky130_fd_sc_hd__buf_2
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _4366_/A vssd1 vssd1 vccd1 vccd1 _8386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6098_/X _6103_/X _6104_/X _6101_/X vssd1 vssd1 vccd1 vccd1 _6105_/X sky130_fd_sc_hd__o211a_1
X_7085_ _7097_/A vssd1 vssd1 vccd1 vccd1 _7085_/X sky130_fd_sc_hd__buf_1
X_4297_ _8417_/Q _4212_/X _4297_/S vssd1 vssd1 vccd1 vccd1 _4298_/A sky130_fd_sc_hd__mux2_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6037_/A sky130_fd_sc_hd__and2_1
XFILLER_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7987_ _7987_/CLK _7987_/D vssd1 vssd1 vccd1 vccd1 _7987_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7745__44 _7746__45/A vssd1 vssd1 vccd1 vccd1 _8595_/CLK sky130_fd_sc_hd__inv_2
X_6869_ _7821_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6869_/X sky130_fd_sc_hd__and2_1
X_8608_ _8608_/CLK _8608_/D vssd1 vssd1 vccd1 vccd1 _8608_/Q sky130_fd_sc_hd__dfxtp_1
X_8539_ _8539_/CLK _8539_/D vssd1 vssd1 vccd1 vccd1 _8539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6616__263 _6616__263/A vssd1 vssd1 vccd1 vccd1 _8023_/CLK sky130_fd_sc_hd__inv_2
Xoutput129 _6015_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput118 _6051_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__buf_2
XFILLER_5_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4220_ _8576_/Q vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__buf_2
X_6319__193 _6321__195/A vssd1 vssd1 vccd1 vccd1 _7905_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4151_ _4151_/A vssd1 vssd1 vccd1 vccd1 _8487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4082_ _8509_/Q _3949_/X _4082_/S vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__mux2_1
X_7910_ _7910_/CLK _7910_/D vssd1 vssd1 vccd1 vccd1 _7910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7841_ _8632_/Q _7826_/X _7840_/X _6423_/X vssd1 vssd1 vccd1 vccd1 _8632_/D sky130_fd_sc_hd__a211o_1
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4984_ _4984_/A _4984_/B vssd1 vssd1 vccd1 vccd1 _8256_/D sky130_fd_sc_hd__nor2_1
X_7772_ _7772_/A vssd1 vssd1 vccd1 vccd1 _8612_/D sky130_fd_sc_hd__clkbuf_1
X_3935_ _8599_/Q _3934_/X _3941_/S vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__mux2_1
X_6723_ _6723_/A vssd1 vssd1 vccd1 vccd1 _8091_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3435_ clkbuf_0__3435_/X vssd1 vssd1 vccd1 vccd1 _7134_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6654_ _6654_/A vssd1 vssd1 vccd1 vccd1 _8050_/D sky130_fd_sc_hd__clkbuf_1
X_5605_ _5604_/X _8076_/Q _5608_/S vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5536_ _5536_/A vssd1 vssd1 vccd1 vccd1 _8129_/D sky130_fd_sc_hd__clkbuf_1
X_8324_ _8324_/CLK _8324_/D vssd1 vssd1 vccd1 vccd1 _8324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5467_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5483_/S sky130_fd_sc_hd__or2_2
X_8255_ _8255_/CLK _8255_/D vssd1 vssd1 vccd1 vccd1 _8255_/Q sky130_fd_sc_hd__dfxtp_1
X_4418_ _4418_/A vssd1 vssd1 vccd1 vccd1 _8363_/D sky130_fd_sc_hd__clkbuf_1
X_8186_ _8186_/CLK _8186_/D vssd1 vssd1 vccd1 vccd1 _8186_/Q sky130_fd_sc_hd__dfxtp_1
X_5398_ _5593_/A vssd1 vssd1 vccd1 vccd1 _5398_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0__3651_ clkbuf_0__3651_/X vssd1 vssd1 vccd1 vccd1 _7504_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4349_ _4127_/X _8393_/Q _4353_/S vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6019_ _6019_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__and2_1
XFILLER_100_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3016_ clkbuf_0__3016_/X vssd1 vssd1 vccd1 vccd1 _6322_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6370_ _6501_/B _7790_/D vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0__3082_ clkbuf_0__3082_/X vssd1 vssd1 vccd1 vccd1 _6356__223/A sky130_fd_sc_hd__clkbuf_4
X_5321_ _7913_/Q _8510_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8040_ _8040_/CLK _8040_/D vssd1 vssd1 vccd1 vccd1 _8040_/Q sky130_fd_sc_hd__dfxtp_1
X_5252_ _8520_/Q _5249_/X _5209_/A _5251_/X vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__o211a_1
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6809__355 _6809__355/A vssd1 vssd1 vccd1 vccd1 _8150_/CLK sky130_fd_sc_hd__inv_2
X_5183_ _5121_/X _5182_/X _5344_/A vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__a21o_1
X_4203_ _8191_/Q vssd1 vssd1 vccd1 vccd1 _4203_/X sky130_fd_sc_hd__clkbuf_4
X_7339__106 _7342__109/A vssd1 vssd1 vccd1 vccd1 _8417_/CLK sky130_fd_sc_hd__inv_2
X_4134_ _8570_/Q vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4065_ _5521_/A vssd1 vssd1 vccd1 vccd1 _5485_/B sky130_fd_sc_hd__buf_4
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7824_ _7836_/A _7824_/B _7824_/C vssd1 vssd1 vccd1 vccd1 _7825_/A sky130_fd_sc_hd__and3_1
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _8260_/Q _8269_/Q _4964_/X _4966_/Y vssd1 vssd1 vccd1 vccd1 _8260_/D sky130_fd_sc_hd__o211a_1
X_7755_ _7755_/A vssd1 vssd1 vccd1 vccd1 _8603_/D sky130_fd_sc_hd__clkbuf_1
X_4898_ _8174_/Q _4865_/X _4713_/A _4897_/X vssd1 vssd1 vccd1 vccd1 _4898_/X sky130_fd_sc_hd__o211a_1
X_6706_ _5967_/A _8084_/Q _6706_/S vssd1 vssd1 vccd1 vccd1 _6707_/A sky130_fd_sc_hd__mux2_1
X_7686_ _7688_/A _7688_/B vssd1 vssd1 vccd1 vccd1 _7687_/A sky130_fd_sc_hd__nand2_1
X_3918_ _7982_/Q _7981_/Q vssd1 vssd1 vccd1 vccd1 _6505_/B sky130_fd_sc_hd__nor2_2
XFILLER_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5519_ _8136_/Q _4504_/X _5519_/S vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__mux2_1
X_8307_ _8307_/CLK _8307_/D vssd1 vssd1 vccd1 vccd1 _8307_/Q sky130_fd_sc_hd__dfxtp_1
X_6499_ _6499_/A _6499_/B vssd1 vssd1 vccd1 vccd1 _6983_/B sky130_fd_sc_hd__nor2_1
X_8238_ _8238_/CLK _8238_/D vssd1 vssd1 vccd1 vccd1 _8238_/Q sky130_fd_sc_hd__dfxtp_1
X_8169_ _8169_/CLK _8169_/D vssd1 vssd1 vccd1 vccd1 _8169_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3248_ _6582_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3248_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7190__70 _7190__70/A vssd1 vssd1 vccd1 vccd1 _8379_/CLK sky130_fd_sc_hd__inv_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _7908_/Q _5604_/A _5872_/S vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4821_ _4821_/A vssd1 vssd1 vccd1 vccd1 _4821_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _4713_/X _4751_/X _4946_/A vssd1 vssd1 vccd1 vccd1 _4752_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4683_ _4683_/A vssd1 vssd1 vccd1 vccd1 _4683_/X sky130_fd_sc_hd__buf_2
XFILLER_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6422_ _6430_/A _6422_/B _6422_/C vssd1 vssd1 vccd1 vccd1 _6422_/Y sky130_fd_sc_hd__nor3_1
XFILLER_115_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6353_ _6353_/A vssd1 vssd1 vccd1 vccd1 _6353_/X sky130_fd_sc_hd__buf_1
XFILLER_103_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6284_ _6284_/A vssd1 vssd1 vccd1 vccd1 _7893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5304_ _3971_/X _5078_/A _5302_/X _5303_/X vssd1 vssd1 vccd1 vccd1 _8209_/D sky130_fd_sc_hd__o211a_1
X_8023_ _8023_/CLK _8023_/D vssd1 vssd1 vccd1 vccd1 _8023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5235_ _8536_/Q _8274_/Q _5352_/S vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5166_ _8592_/Q _8341_/Q _8325_/Q _8365_/Q _5130_/X _5101_/A vssd1 vssd1 vccd1 vccd1
+ _5167_/B sky130_fd_sc_hd__mux4_1
X_4117_ _4117_/A vssd1 vssd1 vccd1 vccd1 _8498_/D sky130_fd_sc_hd__clkbuf_1
X_5097_ _5283_/S vssd1 vssd1 vccd1 vccd1 _5330_/S sky130_fd_sc_hd__buf_2
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4048_ _3952_/X _8524_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4049_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _5999_/A vssd1 vssd1 vccd1 vccd1 _5999_/X sky130_fd_sc_hd__clkbuf_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7807_ _7807_/A vssd1 vssd1 vccd1 vccd1 _8621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7111__506 _7114__509/A vssd1 vssd1 vccd1 vccd1 _8315_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7669_ _8559_/Q vssd1 vssd1 vccd1 vccd1 _7672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7520__8 _7521__9/A vssd1 vssd1 vccd1 vccd1 _8522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3479_ clkbuf_0__3479_/X vssd1 vssd1 vccd1 vccd1 _7226__99/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5035_/S vssd1 vssd1 vccd1 vccd1 _5029_/S sky130_fd_sc_hd__clkbuf_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6971_ _6977_/A vssd1 vssd1 vccd1 vccd1 _6971_/X sky130_fd_sc_hd__buf_1
X_5922_ _5995_/A vssd1 vssd1 vccd1 vccd1 _6060_/A sky130_fd_sc_hd__inv_6
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5853_ _5853_/A vssd1 vssd1 vccd1 vccd1 _7916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3651_ _7479_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3651_/X sky130_fd_sc_hd__clkbuf_16
X_5784_ _7994_/Q _5610_/A _5788_/S vssd1 vssd1 vccd1 vccd1 _5785_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8572_ _8612_/CLK _8572_/D vssd1 vssd1 vccd1 vccd1 _8572_/Q sky130_fd_sc_hd__dfxtp_2
X_4804_ _4672_/A _8265_/Q _4988_/A _4803_/X _4741_/A vssd1 vssd1 vccd1 vccd1 _4804_/X
+ sky130_fd_sc_hd__a221o_1
X_7523_ _7529_/A vssd1 vssd1 vccd1 vccd1 _7523_/X sky130_fd_sc_hd__buf_1
X_4735_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__buf_2
XFILLER_119_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4666_ _4666_/A _4666_/B _4666_/C _4666_/D vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__and4_1
X_4597_ _4463_/X _8300_/Q _4601_/S vssd1 vssd1 vccd1 vccd1 _4598_/A sky130_fd_sc_hd__mux2_1
X_7067__471 _7069__473/A vssd1 vssd1 vccd1 vccd1 _8280_/CLK sky130_fd_sc_hd__inv_2
X_7385_ _8435_/Q _7384_/X _7376_/X _7268_/B vssd1 vssd1 vccd1 vccd1 _7386_/B sky130_fd_sc_hd__o2bb2a_1
X_6405_ _8609_/Q vssd1 vssd1 vccd1 vccd1 _6405_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6267_ _6265_/X _8094_/Q _6261_/X _6263_/X _7883_/Q vssd1 vssd1 vccd1 vccd1 _7883_/D
+ sky130_fd_sc_hd__o32a_1
X_8006_ _8006_/CLK _8006_/D vssd1 vssd1 vccd1 vccd1 _8006_/Q sky130_fd_sc_hd__dfxtp_1
X_6198_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6198_/X sky130_fd_sc_hd__buf_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5218_ _8198_/Q vssd1 vssd1 vccd1 vccd1 _5271_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3016_ _6199_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3016_/X sky130_fd_sc_hd__clkbuf_16
X_5149_ _8214_/Q _5080_/X _5385_/A _5146_/X _5148_/X vssd1 vssd1 vccd1 vccd1 _5149_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6974__403 _6976__405/A vssd1 vssd1 vccd1 vccd1 _8207_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7035__448 _7037__450/A vssd1 vssd1 vccd1 vccd1 _8255_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6610__258 _6611__259/A vssd1 vssd1 vccd1 vccd1 _8018_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6691__308 _6693__310/A vssd1 vssd1 vccd1 vccd1 _8076_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4520_ _8331_/Q _4519_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451_ _4450_/X _8351_/Q _4451_/S vssd1 vssd1 vccd1 vccd1 _4452_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _8379_/D sky130_fd_sc_hd__clkbuf_1
X_6121_ _6117_/X _6118_/X _6119_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6121_/X sky130_fd_sc_hd__o211a_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _8091_/Q _6058_/B vssd1 vssd1 vccd1 vccd1 _6053_/A sky130_fd_sc_hd__and2_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5003_ _5003_/A vssd1 vssd1 vccd1 vccd1 _8248_/D sky130_fd_sc_hd__clkbuf_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6954_ _8567_/Q _6958_/B vssd1 vssd1 vccd1 vccd1 _6955_/A sky130_fd_sc_hd__and2_1
X_5905_ _5905_/A vssd1 vssd1 vccd1 vccd1 _7850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6885_ _7811_/A _7589_/B _6865_/X _6869_/X _6884_/Y vssd1 vssd1 vccd1 vccd1 _6885_/X
+ sky130_fd_sc_hd__a2111o_1
X_8624_ _8631_/CLK _8624_/D vssd1 vssd1 vccd1 vccd1 _8624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5836_ _7923_/Q _4441_/A _5836_/S vssd1 vssd1 vccd1 vccd1 _5837_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5767_ _5767_/A vssd1 vssd1 vccd1 vccd1 _8002_/D sky130_fd_sc_hd__clkbuf_1
X_8555_ _8561_/CLK _8555_/D vssd1 vssd1 vccd1 vccd1 _8555_/Q sky130_fd_sc_hd__dfxtp_2
X_8486_ _8486_/CLK _8486_/D vssd1 vssd1 vccd1 vccd1 _8486_/Q sky130_fd_sc_hd__dfxtp_1
X_4718_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__buf_2
X_5698_ _8032_/Q _5642_/X _5698_/S vssd1 vssd1 vccd1 vccd1 _5699_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4649_ _4649_/A vssd1 vssd1 vccd1 vccd1 _8278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7368_ _7384_/A vssd1 vssd1 vccd1 vccd1 _7368_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7299_ _7379_/A _7379_/B _7817_/A vssd1 vssd1 vccd1 vccd1 _7299_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_wb_clk_i _6197_/A vssd1 vssd1 vccd1 vccd1 _8630_/CLK sky130_fd_sc_hd__clkbuf_16
X_7041__452 _7041__452/A vssd1 vssd1 vccd1 vccd1 _8259_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3316_ clkbuf_0__3316_/X vssd1 vssd1 vccd1 vccd1 _6809__355/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3247_ clkbuf_0__3247_/X vssd1 vssd1 vccd1 vccd1 _6581__235/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6755__316 _6758__319/A vssd1 vssd1 vccd1 vccd1 _8108_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _3951_/A vssd1 vssd1 vccd1 vccd1 _8594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3451_ clkbuf_0__3451_/X vssd1 vssd1 vccd1 vccd1 _7083__484/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3882_ _8201_/Q _8196_/Q vssd1 vssd1 vccd1 vccd1 _5074_/D sky130_fd_sc_hd__or2b_1
X_5621_ _5643_/S vssd1 vssd1 vccd1 vccd1 _5634_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5552_ _5552_/A vssd1 vssd1 vccd1 vccd1 _8122_/D sky130_fd_sc_hd__clkbuf_1
X_8340_ _8340_/CLK _8340_/D vssd1 vssd1 vccd1 vccd1 _8340_/Q sky130_fd_sc_hd__dfxtp_1
X_4503_ _4503_/A vssd1 vssd1 vccd1 vccd1 _8336_/D sky130_fd_sc_hd__clkbuf_1
X_8271_ _8271_/CLK _8271_/D vssd1 vssd1 vccd1 vccd1 _8271_/Q sky130_fd_sc_hd__dfxtp_1
X_5483_ _4450_/X _8155_/Q _5483_/S vssd1 vssd1 vccd1 vccd1 _5484_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4434_ _4434_/A vssd1 vssd1 vccd1 vccd1 _8357_/D sky130_fd_sc_hd__clkbuf_1
X_7222_ _7222_/A vssd1 vssd1 vccd1 vccd1 _7222_/X sky130_fd_sc_hd__buf_1
XFILLER_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4365_ _4123_/X _8386_/Q _4365_/S vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__mux2_1
X_7153_ _7159_/A vssd1 vssd1 vccd1 vccd1 _7153_/X sky130_fd_sc_hd__buf_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _7867_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__or2_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6035_/A vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4296_/A vssd1 vssd1 vccd1 vccd1 _8418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7986_ _7986_/CLK _7986_/D vssd1 vssd1 vccd1 vccd1 _7986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3649_ clkbuf_0__3649_/X vssd1 vssd1 vccd1 vccd1 _7472__145/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6868_ _7552_/B _7552_/C vssd1 vssd1 vccd1 vccd1 _6869_/B sky130_fd_sc_hd__nand2_2
X_5819_ _5819_/A vssd1 vssd1 vccd1 vccd1 _7931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8607_ _8608_/CLK _8607_/D vssd1 vssd1 vccd1 vccd1 _8607_/Q sky130_fd_sc_hd__dfxtp_1
X_8538_ _8538_/CLK _8538_/D vssd1 vssd1 vccd1 vccd1 _8538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8469_ _8469_/CLK _8469_/D vssd1 vssd1 vccd1 vccd1 _8469_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3479_ _7222_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3479_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput119 _6053_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput108 _7903_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__buf_2
X_7048__458 _7049__459/A vssd1 vssd1 vccd1 vccd1 _8265_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4150_ _8487_/Q _3943_/X _4154_/S vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__mux2_1
X_4081_ _4081_/A vssd1 vssd1 vccd1 vccd1 _8510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7840_ _7840_/A _7842_/B _7840_/C vssd1 vssd1 vccd1 vccd1 _7840_/X sky130_fd_sc_hd__and3_1
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _4979_/A _4986_/B _7055_/A vssd1 vssd1 vccd1 vccd1 _4984_/B sky130_fd_sc_hd__a21o_1
X_7771_ _7771_/A _8606_/Q vssd1 vssd1 vccd1 vccd1 _7772_/A sky130_fd_sc_hd__and2_1
X_3934_ _8575_/Q vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6722_ _5982_/A _8091_/Q _6724_/S vssd1 vssd1 vccd1 vccd1 _6723_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3434_ clkbuf_0__3434_/X vssd1 vssd1 vccd1 vccd1 _7005__425/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6653_ _8263_/Q _8249_/D vssd1 vssd1 vccd1 vccd1 _6654_/A sky130_fd_sc_hd__and2_1
X_5604_ _5604_/A vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__buf_2
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5535_ _8129_/Q _4447_/A _5537_/S vssd1 vssd1 vccd1 vccd1 _5536_/A sky130_fd_sc_hd__mux2_1
X_8323_ _8323_/CLK _8323_/D vssd1 vssd1 vccd1 vccd1 _8323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5466_ _5466_/A vssd1 vssd1 vccd1 vccd1 _8164_/D sky130_fd_sc_hd__clkbuf_1
X_8254_ _8254_/CLK _8254_/D vssd1 vssd1 vccd1 vccd1 _8254_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4417_ _4119_/X _8363_/Q _4419_/S vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3650_ clkbuf_0__3650_/X vssd1 vssd1 vccd1 vccd1 _7477__149/A sky130_fd_sc_hd__clkbuf_4
X_8185_ _8185_/CLK _8185_/D vssd1 vssd1 vccd1 vccd1 _8185_/Q sky130_fd_sc_hd__dfxtp_1
X_5397_ _8195_/Q vssd1 vssd1 vccd1 vccd1 _5593_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4348_ _4348_/A vssd1 vssd1 vccd1 vccd1 _8394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4279_ _4279_/A vssd1 vssd1 vccd1 vccd1 _8453_/D sky130_fd_sc_hd__clkbuf_1
X_6018_ _6018_/A vssd1 vssd1 vccd1 vccd1 _6018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _8577_/CLK _7969_/D vssd1 vssd1 vccd1 vccd1 _7969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3015_ clkbuf_0__3015_/X vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7160__546 _7162__548/A vssd1 vssd1 vccd1 vccd1 _8355_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3081_ clkbuf_0__3081_/X vssd1 vssd1 vccd1 vccd1 _6352__220/A sky130_fd_sc_hd__clkbuf_4
X_5320_ _5247_/A _5309_/Y _5312_/Y _5319_/X vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__a31o_1
XFILLER_114_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6768__326 _6769__327/A vssd1 vssd1 vccd1 vccd1 _8118_/CLK sky130_fd_sc_hd__inv_2
X_5251_ _8528_/Q _5103_/B _5250_/X _5294_/A vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4202_ _4202_/A vssd1 vssd1 vccd1 vccd1 _8481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5182_ _8599_/Q _8152_/Q _8125_/Q _8583_/Q _5330_/S _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5182_/X sky130_fd_sc_hd__mux4_2
X_7061__466 _7063__468/A vssd1 vssd1 vccd1 vccd1 _8275_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4133_ _4133_/A vssd1 vssd1 vccd1 vccd1 _8494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4064_ _5382_/A _4064_/B _5150_/A _4004_/A vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__or4bb_4
XFILLER_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7823_ _7723_/A _7778_/A _7826_/A vssd1 vssd1 vccd1 vccd1 _7824_/C sky130_fd_sc_hd__a21o_1
XFILLER_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7754_ _8260_/Q _7836_/A vssd1 vssd1 vccd1 vccd1 _7755_/A sky130_fd_sc_hd__and2_1
XFILLER_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6705_ _6705_/A vssd1 vssd1 vccd1 vccd1 _8083_/D sky130_fd_sc_hd__clkbuf_1
X_4966_ _4985_/B vssd1 vssd1 vccd1 vccd1 _4966_/Y sky130_fd_sc_hd__inv_2
X_4897_ _8235_/Q _4821_/A _4896_/X _4861_/A vssd1 vssd1 vccd1 vccd1 _4897_/X sky130_fd_sc_hd__o22a_1
X_7685_ _8561_/Q _7679_/Y _7682_/X _7684_/X vssd1 vssd1 vccd1 vccd1 _8561_/D sky130_fd_sc_hd__o211a_1
X_3917_ _7960_/Q _7967_/Q _7968_/Q _6375_/B vssd1 vssd1 vccd1 vccd1 _3923_/C sky130_fd_sc_hd__or4_1
XFILLER_32_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5518_ _5518_/A vssd1 vssd1 vccd1 vccd1 _8137_/D sky130_fd_sc_hd__clkbuf_1
X_8306_ _8306_/CLK _8306_/D vssd1 vssd1 vccd1 vccd1 _8306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3316_ _6798_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3316_/X sky130_fd_sc_hd__clkbuf_16
X_6498_ _8616_/Q vssd1 vssd1 vccd1 vccd1 _7575_/A sky130_fd_sc_hd__inv_2
X_8237_ _8237_/CLK _8237_/D vssd1 vssd1 vccd1 vccd1 _8237_/Q sky130_fd_sc_hd__dfxtp_1
X_5449_ _5700_/A _5772_/B vssd1 vssd1 vccd1 vccd1 _5465_/S sky130_fd_sc_hd__or2_2
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8168_ _8168_/CLK _8168_/D vssd1 vssd1 vccd1 vccd1 _8168_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3247_ _6576_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3247_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8099_ _8569_/CLK _8099_/D vssd1 vssd1 vccd1 vccd1 _8099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6205__180 _6205__180/A vssd1 vssd1 vccd1 vccd1 _7849_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4820_ _4820_/A vssd1 vssd1 vccd1 vccd1 _4821_/A sky130_fd_sc_hd__clkbuf_2
X_6919__373 _6920__374/A vssd1 vssd1 vccd1 vccd1 _8169_/CLK sky130_fd_sc_hd__inv_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _8459_/Q _8349_/Q _8062_/Q _8483_/Q _4691_/A _4714_/X vssd1 vssd1 vccd1 vccd1
+ _4751_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4682_ _8254_/Q _4736_/B vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__xor2_4
X_7345__111 _7347__113/A vssd1 vssd1 vccd1 vccd1 _8422_/CLK sky130_fd_sc_hd__inv_2
X_6815__360 _6815__360/A vssd1 vssd1 vccd1 vccd1 _8155_/CLK sky130_fd_sc_hd__inv_2
X_6421_ _6419_/Y _6385_/X _6420_/Y _6398_/X _6387_/A vssd1 vssd1 vccd1 vccd1 _6422_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6283_ _7842_/A _7893_/Q _6291_/S vssd1 vssd1 vccd1 vccd1 _6284_/A sky130_fd_sc_hd__mux2_1
X_5303_ _5377_/A vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__clkbuf_2
X_8022_ _8022_/CLK _8022_/D vssd1 vssd1 vccd1 vccd1 _8022_/Q sky130_fd_sc_hd__dfxtp_1
X_5234_ _5361_/S vssd1 vssd1 vccd1 vccd1 _5352_/S sky130_fd_sc_hd__buf_4
X_5165_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5189_/A sky130_fd_sc_hd__clkbuf_2
X_4116_ _4115_/X _8498_/Q _4124_/S vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6629__274 _6630__275/A vssd1 vssd1 vccd1 vccd1 _8034_/CLK sky130_fd_sc_hd__inv_2
X_5096_ _5222_/B vssd1 vssd1 vccd1 vccd1 _5283_/S sky130_fd_sc_hd__buf_2
XFILLER_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4047_ _4062_/S vssd1 vssd1 vccd1 vccd1 _4056_/S sky130_fd_sc_hd__buf_2
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7806_ _7806_/A _7806_/B vssd1 vssd1 vccd1 vccd1 _7807_/A sky130_fd_sc_hd__or2_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _5999_/A sky130_fd_sc_hd__or2_1
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4949_ _4845_/X _4947_/X _4948_/X vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__o21a_1
X_7668_ _7664_/X _7667_/X _7601_/X vssd1 vssd1 vccd1 vccd1 _8558_/D sky130_fd_sc_hd__o21a_1
X_6619_ _6619_/A vssd1 vssd1 vccd1 vccd1 _6619_/X sky130_fd_sc_hd__buf_1
X_7599_ _7667_/B _7575_/X vssd1 vssd1 vccd1 vccd1 _7599_/X sky130_fd_sc_hd__or2b_1
XFILLER_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3478_ clkbuf_0__3478_/X vssd1 vssd1 vccd1 vccd1 _7219__93/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6970_ _6970_/A vssd1 vssd1 vccd1 vccd1 _6970_/X sky130_fd_sc_hd__buf_1
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5921_ _5921_/A _6195_/C vssd1 vssd1 vccd1 vccd1 _5995_/A sky130_fd_sc_hd__or2_4
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5852_ _4438_/X _7916_/Q _5854_/S vssd1 vssd1 vccd1 vccd1 _5853_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4803_ _4683_/X _4790_/X _4794_/X _4802_/X vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__a31o_2
X_5783_ _5783_/A vssd1 vssd1 vccd1 vccd1 _7995_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3650_ _7473_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3650_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7536__21 _7537__22/A vssd1 vssd1 vccd1 vccd1 _8535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8571_ _8612_/CLK _8571_/D vssd1 vssd1 vccd1 vccd1 _8571_/Q sky130_fd_sc_hd__dfxtp_2
X_4734_ _4730_/X _4732_/X _4796_/A vssd1 vssd1 vccd1 vccd1 _4734_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ _4822_/A vssd1 vssd1 vccd1 vccd1 _4665_/X sky130_fd_sc_hd__clkbuf_4
X_4596_ _4596_/A vssd1 vssd1 vccd1 vccd1 _8301_/D sky130_fd_sc_hd__clkbuf_1
X_7384_ _7384_/A vssd1 vssd1 vccd1 vccd1 _7384_/X sky130_fd_sc_hd__clkbuf_2
X_6404_ _6872_/A _6403_/X _6373_/X vssd1 vssd1 vccd1 vccd1 _6408_/B sky130_fd_sc_hd__a21oi_1
X_6335_ _6341_/A vssd1 vssd1 vccd1 vccd1 _6335_/X sky130_fd_sc_hd__buf_1
X_8005_ _8005_/CLK _8005_/D vssd1 vssd1 vccd1 vccd1 _8005_/Q sky130_fd_sc_hd__dfxtp_1
X_6266_ _6265_/X _8093_/Q _6261_/X _6263_/X _7882_/Q vssd1 vssd1 vccd1 vccd1 _7882_/D
+ sky130_fd_sc_hd__o32a_1
X_6197_ _6197_/A vssd1 vssd1 vccd1 vccd1 _6197_/X sky130_fd_sc_hd__buf_1
X_5217_ _5217_/A vssd1 vssd1 vccd1 vccd1 _5387_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3015_ _6198_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3015_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5148_ _5148_/A vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _8216_/Q vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__inv_2
XFILLER_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7224__97 _7224__97/A vssd1 vssd1 vccd1 vccd1 _8406_/CLK sky130_fd_sc_hd__inv_2
X_7074__476 _7075__477/A vssd1 vssd1 vccd1 vccd1 _8285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7478__150 _7478__150/A vssd1 vssd1 vccd1 vccd1 _8489_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6578__232 _6578__232/A vssd1 vssd1 vccd1 vccd1 _7992_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4450_/A vssd1 vssd1 vccd1 vccd1 _4450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4381_ _8379_/Q _4226_/X _4383_/S vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__mux2_1
X_6120_ _6173_/A vssd1 vssd1 vccd1 vccd1 _6120_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8661__226 vssd1 vssd1 vccd1 vccd1 _8661__226/HI core1Index[6] sky130_fd_sc_hd__conb_1
X_6051_ _6051_/A vssd1 vssd1 vccd1 vccd1 _6051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5002_ _8248_/Q _4507_/X _5010_/S vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__mux2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6953_ _6953_/A vssd1 vssd1 vccd1 vccd1 _8192_/D sky130_fd_sc_hd__clkbuf_1
X_5904_ _4197_/X _7850_/Q _5908_/S vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6884_ _7821_/A _6869_/B _7582_/A _6881_/X _7582_/B vssd1 vssd1 vccd1 vccd1 _6884_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5835_ _5835_/A vssd1 vssd1 vccd1 vccd1 _7924_/D sky130_fd_sc_hd__clkbuf_1
X_8623_ _8623_/CLK _8623_/D vssd1 vssd1 vccd1 vccd1 _8623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5766_ _8002_/Q _5636_/X _5770_/S vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8554_ _8554_/CLK _8554_/D vssd1 vssd1 vccd1 vccd1 _8554_/Q sky130_fd_sc_hd__dfxtp_1
X_8485_ _8485_/CLK _8485_/D vssd1 vssd1 vccd1 vccd1 _8485_/Q sky130_fd_sc_hd__dfxtp_1
X_4717_ _4736_/B _4717_/B vssd1 vssd1 vccd1 vccd1 _4869_/A sky130_fd_sc_hd__nor2_1
X_5697_ _5697_/A vssd1 vssd1 vccd1 vccd1 _8033_/D sky130_fd_sc_hd__clkbuf_1
X_7436_ _7436_/A vssd1 vssd1 vccd1 vccd1 _7436_/X sky130_fd_sc_hd__buf_1
X_4648_ _8278_/Q _4481_/X _4656_/S vssd1 vssd1 vccd1 vccd1 _4649_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4579_ _4435_/X _8308_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__mux2_1
X_7367_ _7371_/A _7367_/B vssd1 vssd1 vccd1 vccd1 _8429_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7298_ _7308_/A _7308_/B _8433_/Q vssd1 vssd1 vccd1 vccd1 _7379_/B sky130_fd_sc_hd__a21o_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6249_ _6423_/A vssd1 vssd1 vccd1 vccd1 _6249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3315_ clkbuf_0__3315_/X vssd1 vssd1 vccd1 vccd1 _6822_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3246_ clkbuf_0__3246_/X vssd1 vssd1 vccd1 vccd1 _6572__227/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7530__16 _7532__18/A vssd1 vssd1 vccd1 vccd1 _8530_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7124__517 _7124__517/A vssd1 vssd1 vccd1 vccd1 _8326_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3950_ _8594_/Q _3949_/X _3950_/S vssd1 vssd1 vccd1 vccd1 _3951_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3450_ clkbuf_0__3450_/X vssd1 vssd1 vccd1 vccd1 _7075__477/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3881_ _8196_/Q _3983_/B vssd1 vssd1 vccd1 vccd1 _5074_/C sky130_fd_sc_hd__or2b_1
X_5620_ _5718_/B _5772_/A vssd1 vssd1 vccd1 vccd1 _5643_/S sky130_fd_sc_hd__nor2_2
X_5551_ _8122_/Q _4444_/A _5555_/S vssd1 vssd1 vccd1 vccd1 _5552_/A sky130_fd_sc_hd__mux2_1
X_4502_ _8336_/Q _4501_/X _4505_/S vssd1 vssd1 vccd1 vccd1 _4503_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8270_ _8270_/CLK _8270_/D vssd1 vssd1 vccd1 vccd1 _8270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5482_ _5482_/A vssd1 vssd1 vccd1 vccd1 _8156_/D sky130_fd_sc_hd__clkbuf_1
X_4433_ _4432_/X _8357_/Q _4442_/S vssd1 vssd1 vccd1 vccd1 _4434_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4364_ _4364_/A vssd1 vssd1 vccd1 vccd1 _8387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _7942_/Q input31/X _6106_/S vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__mux2_1
X_4295_ _8418_/Q _4209_/X _4297_/S vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__mux2_1
X_6034_ _6034_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6035_/A sky130_fd_sc_hd__and2_1
XFILLER_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7985_ _7985_/CLK _7985_/D vssd1 vssd1 vccd1 vccd1 _7985_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3648_ clkbuf_0__3648_/X vssd1 vssd1 vccd1 vccd1 _7463__137/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6867_ _8549_/Q _6850_/A _6852_/B _8550_/Q vssd1 vssd1 vccd1 vccd1 _7552_/C sky130_fd_sc_hd__a31o_1
X_6798_ _6822_/A vssd1 vssd1 vccd1 vccd1 _6798_/X sky130_fd_sc_hd__buf_1
X_5818_ _5607_/X _7931_/Q _5818_/S vssd1 vssd1 vccd1 vccd1 _5819_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8606_ _8612_/CLK _8606_/D vssd1 vssd1 vccd1 vccd1 _8606_/Q sky130_fd_sc_hd__dfxtp_1
X_8537_ _8537_/CLK _8537_/D vssd1 vssd1 vccd1 vccd1 _8537_/Q sky130_fd_sc_hd__dfxtp_1
X_5749_ _5749_/A vssd1 vssd1 vccd1 vccd1 _8010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8468_ _8468_/CLK _8468_/D vssd1 vssd1 vccd1 vccd1 _8468_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3478_ _7216_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3478_/X sky130_fd_sc_hd__clkbuf_16
X_8399_ _8399_/CLK _8399_/D vssd1 vssd1 vccd1 vccd1 _8399_/Q sky130_fd_sc_hd__dfxtp_1
X_7419_ _8446_/Q _7424_/B vssd1 vssd1 vccd1 vccd1 _7419_/X sky130_fd_sc_hd__or2_1
XFILLER_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6761__321 _6763__323/A vssd1 vssd1 vccd1 vccd1 _8113_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7751__49 _7751__49/A vssd1 vssd1 vccd1 vccd1 _8600_/CLK sky130_fd_sc_hd__inv_2
X_6913__368 _6915__370/A vssd1 vssd1 vccd1 vccd1 _8164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput109 _6011_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4080_ _8510_/Q _3946_/X _4082_/S vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6623__269 _6624__270/A vssd1 vssd1 vccd1 vccd1 _8029_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4982_ _4969_/B _4985_/B _4980_/Y _7055_/A vssd1 vssd1 vccd1 vccd1 _8257_/D sky130_fd_sc_hd__a211oi_1
X_7770_ _7770_/A vssd1 vssd1 vccd1 vccd1 _8611_/D sky130_fd_sc_hd__clkbuf_1
X_6326__199 _6327__200/A vssd1 vssd1 vccd1 vccd1 _7911_/CLK sky130_fd_sc_hd__inv_2
X_3933_ _3933_/A vssd1 vssd1 vccd1 vccd1 _8600_/D sky130_fd_sc_hd__clkbuf_1
X_6721_ _6721_/A vssd1 vssd1 vccd1 vccd1 _8090_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8570_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1_0__3433_ clkbuf_0__3433_/X vssd1 vssd1 vccd1 vccd1 _6997__418/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6652_ _6652_/A vssd1 vssd1 vccd1 vccd1 _8049_/D sky130_fd_sc_hd__clkbuf_1
X_5603_ _5603_/A vssd1 vssd1 vccd1 vccd1 _8077_/D sky130_fd_sc_hd__clkbuf_1
X_8322_ _8322_/CLK _8322_/D vssd1 vssd1 vccd1 vccd1 _8322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5534_ _5534_/A vssd1 vssd1 vccd1 vccd1 _8130_/D sky130_fd_sc_hd__clkbuf_1
X_8667__232 vssd1 vssd1 vccd1 vccd1 _8667__232/HI manufacturerID[4] sky130_fd_sc_hd__conb_1
X_5465_ _5428_/X _8164_/Q _5465_/S vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__mux2_1
X_8253_ _8253_/CLK _8253_/D vssd1 vssd1 vccd1 vccd1 _8253_/Q sky130_fd_sc_hd__dfxtp_1
X_8184_ _8184_/CLK _8184_/D vssd1 vssd1 vccd1 vccd1 _8184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7204_ _7210_/A vssd1 vssd1 vccd1 vccd1 _7204_/X sky130_fd_sc_hd__buf_1
X_4416_ _4416_/A vssd1 vssd1 vccd1 vccd1 _8364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7135_ _7159_/A vssd1 vssd1 vccd1 vccd1 _7135_/X sky130_fd_sc_hd__buf_1
X_5396_ _5321_/S _5385_/X _5395_/Y vssd1 vssd1 vccd1 vccd1 _8196_/D sky130_fd_sc_hd__a21oi_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4347_ _4123_/X _8394_/Q _4347_/S vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__mux2_1
X_7066_ _7066_/A vssd1 vssd1 vccd1 vccd1 _7066_/X sky130_fd_sc_hd__buf_1
X_4278_ _8453_/Q _4212_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__mux2_1
X_6017_ _6017_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__and2_1
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _8570_/CLK _7968_/D vssd1 vssd1 vccd1 vccd1 _7968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7899_ _8631_/CLK _7899_/D vssd1 vssd1 vccd1 vccd1 _7899_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3014_ clkbuf_0__3014_/X vssd1 vssd1 vccd1 vccd1 _7541_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3080_ clkbuf_0__3080_/X vssd1 vssd1 vccd1 vccd1 _6346__215/A sky130_fd_sc_hd__clkbuf_4
X_5250_ _7915_/Q _8512_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4201_ _8481_/Q _4200_/X _4204_/S vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5181_ _7925_/Q _8133_/Q _8412_/Q _8160_/Q _5313_/S _5110_/X vssd1 vssd1 vccd1 vccd1
+ _5181_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _4131_/X _8494_/Q _4136_/S vssd1 vssd1 vccd1 vccd1 _4133_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4063_ _4063_/A vssd1 vssd1 vccd1 vccd1 _8517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7137__527 _7139__529/A vssd1 vssd1 vccd1 vccd1 _8336_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7822_ _7842_/C vssd1 vssd1 vccd1 vccd1 _7826_/A sky130_fd_sc_hd__inv_2
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7753_ _7757_/A _7753_/B vssd1 vssd1 vccd1 vccd1 _8602_/D sky130_fd_sc_hd__nor2_1
X_4965_ _4965_/A vssd1 vssd1 vccd1 vccd1 _4985_/B sky130_fd_sc_hd__clkbuf_2
X_6704_ _7809_/A _8083_/Q _6706_/S vssd1 vssd1 vccd1 vccd1 _6705_/A sky130_fd_sc_hd__mux2_1
X_3916_ _6454_/A _6368_/A _7959_/Q vssd1 vssd1 vccd1 vccd1 _6375_/B sky130_fd_sc_hd__o21ai_1
X_4896_ _4849_/A _8166_/Q _7994_/Q _4847_/A vssd1 vssd1 vccd1 vccd1 _4896_/X sky130_fd_sc_hd__a22o_1
X_7176__58 _7177__59/A vssd1 vssd1 vccd1 vccd1 _8367_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7684_ _7684_/A vssd1 vssd1 vccd1 vccd1 _7684_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6566_ _6225_/X _6306_/B _7757_/A vssd1 vssd1 vccd1 vccd1 _7983_/D sky130_fd_sc_hd__a21oi_1
X_5517_ _8137_/Q _4501_/X _5519_/S vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__mux2_1
X_8305_ _8305_/CLK _8305_/D vssd1 vssd1 vccd1 vccd1 _8305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3315_ _6797_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3315_/X sky130_fd_sc_hd__clkbuf_16
X_8236_ _8236_/CLK _8236_/D vssd1 vssd1 vccd1 vccd1 _8236_/Q sky130_fd_sc_hd__dfxtp_1
X_6497_ _8617_/Q vssd1 vssd1 vccd1 vccd1 _6500_/A sky130_fd_sc_hd__inv_2
X_5448_ _5448_/A vssd1 vssd1 vccd1 vccd1 _8172_/D sky130_fd_sc_hd__clkbuf_1
X_8167_ _8167_/CLK _8167_/D vssd1 vssd1 vccd1 vccd1 _8167_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3246_ _6570_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3246_/X sky130_fd_sc_hd__clkbuf_16
X_5379_ _5147_/A _5382_/A _7757_/B _4004_/A vssd1 vssd1 vccd1 vccd1 _5380_/B sky130_fd_sc_hd__a31o_1
X_8641__257 vssd1 vssd1 vccd1 vccd1 partID[11] _8641__257/LO sky130_fd_sc_hd__conb_1
X_8098_ _8569_/CLK _8098_/D vssd1 vssd1 vccd1 vccd1 _8098_/Q sky130_fd_sc_hd__dfxtp_1
X_7472__145 _7472__145/A vssd1 vssd1 vccd1 vccd1 _8484_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6572__227 _6572__227/A vssd1 vssd1 vccd1 vccd1 _7987_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6774__331 _6778__335/A vssd1 vssd1 vccd1 vccd1 _8123_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _8301_/Q _8285_/Q _8247_/Q _8317_/Q _4710_/X _4702_/X vssd1 vssd1 vccd1 vccd1
+ _4750_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4681_ _4716_/A _4704_/A vssd1 vssd1 vccd1 vccd1 _4736_/B sky130_fd_sc_hd__and2_2
X_6420_ _8052_/Q _6395_/X _6382_/X vssd1 vssd1 vccd1 vccd1 _6420_/Y sky130_fd_sc_hd__a21oi_1
X_5302_ _8209_/Q _5081_/A _5386_/A _5301_/X _5148_/A vssd1 vssd1 vccd1 vccd1 _5302_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6282_ _6297_/S vssd1 vssd1 vccd1 vccd1 _6291_/S sky130_fd_sc_hd__buf_2
X_8021_ _8021_/CLK _8021_/D vssd1 vssd1 vccd1 vccd1 _8021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5233_ _5294_/A vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__clkbuf_2
X_5164_ _5162_/X _5163_/X _5246_/S vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__mux2_1
X_6926__378 _6927__379/A vssd1 vssd1 vccd1 vccd1 _8174_/CLK sky130_fd_sc_hd__inv_2
X_4115_ _4435_/A vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5095_ _5095_/A vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4046_ _4355_/A _5844_/B vssd1 vssd1 vccd1 vccd1 _4062_/S sky130_fd_sc_hd__or2_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7805_ _7548_/A _7817_/B _7818_/B _5967_/A vssd1 vssd1 vccd1 vccd1 _7806_/B sky130_fd_sc_hd__a22o_1
X_5997_ _5997_/A vssd1 vssd1 vccd1 vccd1 _5997_/X sky130_fd_sc_hd__clkbuf_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4948_ _8477_/Q _4680_/A _4817_/A _8453_/Q _4687_/A vssd1 vssd1 vccd1 vccd1 _4948_/X
+ sky130_fd_sc_hd__o221a_1
X_4879_ _8018_/Q _4821_/X _4878_/X _4861_/X vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__o22a_1
X_7667_ _6905_/B _7667_/B _7682_/A vssd1 vssd1 vccd1 vccd1 _7667_/X sky130_fd_sc_hd__and3b_1
XFILLER_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6636__279 _6636__279/A vssd1 vssd1 vccd1 vccd1 _8039_/CLK sky130_fd_sc_hd__inv_2
X_7598_ _7642_/A vssd1 vssd1 vccd1 vccd1 _7667_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6549_ _6549_/A vssd1 vssd1 vccd1 vccd1 _7978_/D sky130_fd_sc_hd__clkbuf_1
X_8219_ _8219_/CLK _8219_/D vssd1 vssd1 vccd1 vccd1 _8219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3477_ clkbuf_0__3477_/X vssd1 vssd1 vccd1 vccd1 _7214__89/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5920_ _6195_/B _5918_/B _5919_/X _7844_/Q vssd1 vssd1 vccd1 vccd1 _6195_/C sky130_fd_sc_hd__a31o_4
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5851_ _5851_/A vssd1 vssd1 vccd1 vccd1 _7917_/D sky130_fd_sc_hd__clkbuf_1
X_4802_ _4796_/X _4798_/X _4801_/X _4735_/X _4737_/X vssd1 vssd1 vccd1 vccd1 _4802_/X
+ sky130_fd_sc_hd__o221a_1
X_5782_ _7995_/Q _5607_/A _5782_/S vssd1 vssd1 vccd1 vccd1 _5783_/A sky130_fd_sc_hd__mux2_1
X_8570_ _8570_/CLK _8570_/D vssd1 vssd1 vccd1 vccd1 _8570_/Q sky130_fd_sc_hd__dfxtp_2
X_4733_ _4733_/A vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__buf_2
XFILLER_119_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664_ _4852_/A vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__clkbuf_2
X_6403_ _6403_/A vssd1 vssd1 vccd1 vccd1 _6403_/X sky130_fd_sc_hd__clkbuf_2
X_4595_ _4460_/X _8301_/Q _4601_/S vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__mux2_1
X_7383_ _7386_/A _7383_/B vssd1 vssd1 vccd1 vccd1 _8434_/D sky130_fd_sc_hd__nor2_1
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _6390_/A vssd1 vssd1 vccd1 vccd1 _6265_/X sky130_fd_sc_hd__buf_2
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8004_ _8004_/CLK _8004_/D vssd1 vssd1 vccd1 vccd1 _8004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5216_ _5216_/A vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__clkbuf_2
X_6196_ _6196_/A vssd1 vssd1 vccd1 vccd1 _7844_/D sky130_fd_sc_hd__buf_2
XFILLER_111_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3014_ _6197_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3014_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5147_ _5147_/A _7410_/A vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__and2_1
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5078_ _5078_/A vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4029_ _4044_/S vssd1 vssd1 vccd1 vccd1 _4038_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_71_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7719_ _7719_/A _7723_/B _7723_/C vssd1 vssd1 vccd1 vccd1 _7720_/A sky130_fd_sc_hd__and3_1
XFILLER_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6981__409 _6982__410/A vssd1 vssd1 vccd1 vccd1 _8213_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7485__155 _7485__155/A vssd1 vssd1 vccd1 vccd1 _8494_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4380_ _4380_/A vssd1 vssd1 vccd1 vccd1 _8380_/D sky130_fd_sc_hd__clkbuf_1
X_6331__202 _6331__202/A vssd1 vssd1 vccd1 vccd1 _7914_/CLK sky130_fd_sc_hd__inv_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _8090_/Q _6058_/B vssd1 vssd1 vccd1 vccd1 _6051_/A sky130_fd_sc_hd__and2_1
XFILLER_86_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5001_ _5016_/S vssd1 vssd1 vccd1 vccd1 _5010_/S sky130_fd_sc_hd__buf_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952_ _8566_/Q _6958_/B vssd1 vssd1 vccd1 vccd1 _6953_/A sky130_fd_sc_hd__and2_1
X_5903_ _5903_/A vssd1 vssd1 vccd1 vccd1 _7851_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3664_ clkbuf_0__3664_/X vssd1 vssd1 vccd1 vccd1 _7543__26/A sky130_fd_sc_hd__clkbuf_4
X_6883_ _8629_/Q _7564_/B vssd1 vssd1 vccd1 vccd1 _7582_/B sky130_fd_sc_hd__xor2_1
X_5834_ _7924_/Q _4438_/A _5836_/S vssd1 vssd1 vccd1 vccd1 _5835_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8622_ _8622_/CLK _8622_/D vssd1 vssd1 vccd1 vccd1 _8622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5765_ _5765_/A vssd1 vssd1 vccd1 vccd1 _8003_/D sky130_fd_sc_hd__clkbuf_1
X_8553_ _8553_/CLK _8553_/D vssd1 vssd1 vccd1 vccd1 _8553_/Q sky130_fd_sc_hd__dfxtp_2
X_8484_ _8484_/CLK _8484_/D vssd1 vssd1 vccd1 vccd1 _8484_/Q sky130_fd_sc_hd__dfxtp_1
X_7504_ _7504_/A vssd1 vssd1 vccd1 vccd1 _7504_/X sky130_fd_sc_hd__buf_1
X_4716_ _4716_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4717_/B sky130_fd_sc_hd__nor2_1
X_5696_ _8033_/Q _5639_/X _5698_/S vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__mux2_1
X_4647_ _4662_/S vssd1 vssd1 vccd1 vccd1 _4656_/S sky130_fd_sc_hd__buf_2
X_7366_ _7282_/A _7352_/X _7360_/X _7283_/B vssd1 vssd1 vccd1 vccd1 _7367_/B sky130_fd_sc_hd__o2bb2a_1
X_4578_ _4578_/A vssd1 vssd1 vccd1 vccd1 _8309_/D sky130_fd_sc_hd__clkbuf_1
X_6317_ _7407_/D _6314_/X _7358_/A _7387_/A vssd1 vssd1 vccd1 vccd1 _7903_/D sky130_fd_sc_hd__a211o_4
X_7297_ _7297_/A _7297_/B _7297_/C _7297_/D vssd1 vssd1 vccd1 vccd1 _7313_/C sky130_fd_sc_hd__and4_1
X_7080__481 _7084__485/A vssd1 vssd1 vccd1 vccd1 _8290_/CLK sky130_fd_sc_hd__inv_2
X_6248_ _6240_/X _8082_/Q _6245_/X _6247_/X _7871_/Q vssd1 vssd1 vccd1 vccd1 _7871_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6179_ _7887_/Q _6175_/X _6176_/X _6178_/X _6173_/X vssd1 vssd1 vccd1 vccd1 _6179_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3314_ clkbuf_0__3314_/X vssd1 vssd1 vccd1 vccd1 _6794__348/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3245_ clkbuf_0__3245_/X vssd1 vssd1 vccd1 vccd1 _6576_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8631_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8684__249 vssd1 vssd1 vccd1 vccd1 _8684__249/HI versionID[3] sky130_fd_sc_hd__conb_1
XFILLER_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7018__434 _7019__435/A vssd1 vssd1 vccd1 vccd1 _8240_/CLK sky130_fd_sc_hd__inv_2
X_3880_ _3983_/B vssd1 vssd1 vccd1 vccd1 _5382_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5550_ _5550_/A vssd1 vssd1 vccd1 vccd1 _8123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5481_ _4447_/X _8156_/Q _5483_/S vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__mux2_1
X_4501_ _8571_/Q vssd1 vssd1 vccd1 vccd1 _4501_/X sky130_fd_sc_hd__clkbuf_4
X_4432_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4432_/X sky130_fd_sc_hd__clkbuf_4
X_4363_ _4119_/X _8387_/Q _4365_/S vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4294_ _4294_/A vssd1 vssd1 vccd1 vccd1 _8419_/D sky130_fd_sc_hd__clkbuf_1
X_6102_ _6098_/X _6099_/X _6100_/X _6101_/X vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__o211a_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6033_/A vssd1 vssd1 vccd1 vccd1 _6033_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7984_ _7984_/CLK _7984_/D vssd1 vssd1 vccd1 vccd1 _7984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6935_ _6935_/A vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__buf_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3647_ clkbuf_0__3647_/X vssd1 vssd1 vccd1 vccd1 _7460__135/A sky130_fd_sc_hd__clkbuf_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6866_ _6886_/B _6886_/C vssd1 vssd1 vccd1 vccd1 _7552_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5817_ _5817_/A vssd1 vssd1 vccd1 vccd1 _7932_/D sky130_fd_sc_hd__clkbuf_1
X_6797_ _6797_/A vssd1 vssd1 vccd1 vccd1 _6797_/X sky130_fd_sc_hd__buf_1
XFILLER_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8605_ _8612_/CLK _8605_/D vssd1 vssd1 vccd1 vccd1 _8605_/Q sky130_fd_sc_hd__dfxtp_1
X_8536_ _8536_/CLK _8536_/D vssd1 vssd1 vccd1 vccd1 _8536_/Q sky130_fd_sc_hd__dfxtp_1
X_5748_ _8010_/Q _5636_/X _5752_/S vssd1 vssd1 vccd1 vccd1 _5749_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6338__208 _6338__208/A vssd1 vssd1 vccd1 vccd1 _7920_/CLK sky130_fd_sc_hd__inv_2
X_8467_ _8467_/CLK _8467_/D vssd1 vssd1 vccd1 vccd1 _8467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5679_ _5679_/A vssd1 vssd1 vccd1 vccd1 _8041_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3477_ _7210_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3477_/X sky130_fd_sc_hd__clkbuf_16
X_8398_ _8398_/CLK _8398_/D vssd1 vssd1 vccd1 vccd1 _8398_/Q sky130_fd_sc_hd__dfxtp_1
X_7418_ _8208_/Q _7756_/B _7413_/X _7417_/X _7336_/X vssd1 vssd1 vccd1 vccd1 _8445_/D
+ sky130_fd_sc_hd__o311a_1
X_7349_ _8616_/Q _7349_/B vssd1 vssd1 vccd1 vccd1 _7350_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7736__36 _7738__38/A vssd1 vssd1 vccd1 vccd1 _8587_/CLK sky130_fd_sc_hd__inv_2
X_7130__522 _7132__524/A vssd1 vssd1 vccd1 vccd1 _8331_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7087__487 _7089__489/A vssd1 vssd1 vccd1 vccd1 _8296_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4981_ _4981_/A vssd1 vssd1 vccd1 vccd1 _7055_/A sky130_fd_sc_hd__inv_2
X_3932_ _8600_/Q _3931_/X _3941_/S vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6720_ _5980_/A _8090_/Q _6724_/S vssd1 vssd1 vccd1 vccd1 _6721_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6651_ _8262_/Q _8249_/D vssd1 vssd1 vccd1 vccd1 _6652_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3432_ clkbuf_0__3432_/X vssd1 vssd1 vccd1 vccd1 _6991__413/A sky130_fd_sc_hd__clkbuf_4
X_5602_ _5601_/X _8077_/Q _5608_/S vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__mux2_1
X_6582_ _6594_/A vssd1 vssd1 vccd1 vccd1 _6582_/X sky130_fd_sc_hd__buf_1
X_5533_ _8130_/Q _4444_/A _5537_/S vssd1 vssd1 vccd1 vccd1 _5534_/A sky130_fd_sc_hd__mux2_1
X_8321_ _8321_/CLK _8321_/D vssd1 vssd1 vccd1 vccd1 _8321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5464_ _5464_/A vssd1 vssd1 vccd1 vccd1 _8165_/D sky130_fd_sc_hd__clkbuf_1
X_8252_ _8252_/CLK _8252_/D vssd1 vssd1 vccd1 vccd1 _8252_/Q sky130_fd_sc_hd__dfxtp_1
X_4415_ _4115_/X _8364_/Q _4419_/S vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__mux2_1
X_8183_ _8183_/CLK _8183_/D vssd1 vssd1 vccd1 vccd1 _8183_/Q sky130_fd_sc_hd__dfxtp_1
X_5395_ _5321_/S _5393_/A _5377_/A vssd1 vssd1 vccd1 vccd1 _5395_/Y sky130_fd_sc_hd__o21ai_1
X_4346_ _4346_/A vssd1 vssd1 vccd1 vccd1 _8395_/D sky130_fd_sc_hd__clkbuf_1
X_7134_ _7134_/A vssd1 vssd1 vccd1 vccd1 _7134_/X sky130_fd_sc_hd__buf_1
XFILLER_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4277_ _4277_/A vssd1 vssd1 vccd1 vccd1 _8454_/D sky130_fd_sc_hd__clkbuf_1
X_6016_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ _8570_/CLK _7967_/D vssd1 vssd1 vccd1 vccd1 _7967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7898_ _8439_/CLK _7898_/D vssd1 vssd1 vccd1 vccd1 _7898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6849_ _7555_/B _7555_/C vssd1 vssd1 vccd1 vccd1 _7589_/B sky130_fd_sc_hd__nand2_2
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8519_ _8519_/CLK _8519_/D vssd1 vssd1 vccd1 vccd1 _8519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4200_ _8192_/Q vssd1 vssd1 vccd1 vccd1 _4200_/X sky130_fd_sc_hd__clkbuf_4
X_5180_ _5095_/X _5177_/X _5179_/X vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4131_ _4447_/A vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4062_ _3977_/X _8517_/Q _4062_/S vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ _7821_/A _7842_/C vssd1 vssd1 vccd1 vccd1 _7824_/B sky130_fd_sc_hd__or2_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4964_ _7053_/C vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6703_ _6703_/A vssd1 vssd1 vccd1 vccd1 _8082_/D sky130_fd_sc_hd__clkbuf_1
X_3915_ _8144_/Q _6361_/A vssd1 vssd1 vccd1 vccd1 _6384_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0__3415_ clkbuf_0__3415_/X vssd1 vssd1 vccd1 vccd1 _6942__391/A sky130_fd_sc_hd__clkbuf_4
X_4895_ _4831_/X _7986_/Q _4838_/X _8219_/Q _4758_/A vssd1 vssd1 vccd1 vccd1 _4895_/X
+ sky130_fd_sc_hd__o221a_1
X_7683_ _7683_/A vssd1 vssd1 vccd1 vccd1 _7684_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6565_ _7806_/A vssd1 vssd1 vccd1 vccd1 _7757_/A sky130_fd_sc_hd__buf_6
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5516_ _5516_/A vssd1 vssd1 vccd1 vccd1 _8138_/D sky130_fd_sc_hd__clkbuf_1
X_8304_ _8304_/CLK _8304_/D vssd1 vssd1 vccd1 vccd1 _8304_/Q sky130_fd_sc_hd__dfxtp_1
X_7506__172 _7506__172/A vssd1 vssd1 vccd1 vccd1 _8511_/CLK sky130_fd_sc_hd__inv_2
X_6496_ _7957_/Q _6359_/X _6459_/X vssd1 vssd1 vccd1 vccd1 _7957_/D sky130_fd_sc_hd__a21o_1
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3314_ _6791_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3314_/X sky130_fd_sc_hd__clkbuf_16
X_5447_ _5428_/X _8172_/Q _5447_/S vssd1 vssd1 vccd1 vccd1 _5448_/A sky130_fd_sc_hd__mux2_1
X_8235_ _8235_/CLK _8235_/D vssd1 vssd1 vccd1 vccd1 _8235_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3245_ _6569_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3245_/X sky130_fd_sc_hd__clkbuf_16
X_8166_ _8166_/CLK _8166_/D vssd1 vssd1 vccd1 vccd1 _8166_/Q sky130_fd_sc_hd__dfxtp_1
X_5378_ _5378_/A vssd1 vssd1 vccd1 vccd1 _8203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4329_ _4329_/A vssd1 vssd1 vccd1 vccd1 _8402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8097_ _8569_/CLK _8097_/D vssd1 vssd1 vccd1 vccd1 _8097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _4680_/A _4807_/A vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7181__62 _7184__65/A vssd1 vssd1 vccd1 vccd1 _8371_/CLK sky130_fd_sc_hd__inv_2
X_5301_ _5387_/B _5279_/X _5286_/X _5300_/X vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__a31o_1
X_7143__532 _7144__533/A vssd1 vssd1 vccd1 vccd1 _8341_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6281_ _6281_/A _6732_/B vssd1 vssd1 vccd1 vccd1 _6297_/S sky130_fd_sc_hd__nand2_2
X_8020_ _8020_/CLK _8020_/D vssd1 vssd1 vccd1 vccd1 _8020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5232_ _5232_/A vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__clkbuf_2
X_5163_ _8389_/Q _8381_/Q _8373_/Q _8397_/Q _5138_/X _5131_/X vssd1 vssd1 vccd1 vccd1
+ _5163_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _8575_/Q vssd1 vssd1 vccd1 vccd1 _4435_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5094_ _5246_/S vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4045_ _4045_/A vssd1 vssd1 vccd1 vccd1 _8525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7804_ _7802_/Y _7803_/Y _7800_/X vssd1 vssd1 vccd1 vccd1 _8620_/D sky130_fd_sc_hd__a21oi_1
X_5996_ _5996_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _5997_/A sky130_fd_sc_hd__or2_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4947_ _8343_/Q _4849_/X _4847_/X _8056_/Q vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7735_ _7735_/A vssd1 vssd1 vccd1 vccd1 _7735_/X sky130_fd_sc_hd__buf_1
X_4878_ _4812_/A _8114_/Q _8066_/Q _4853_/A vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__a22o_1
X_7666_ _7677_/A vssd1 vssd1 vccd1 vccd1 _7682_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6675__296 _6678__299/A vssd1 vssd1 vccd1 vccd1 _8064_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7597_ _7597_/A vssd1 vssd1 vccd1 vccd1 _8541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6548_ _8093_/Q _7978_/Q _6548_/S vssd1 vssd1 vccd1 vccd1 _6549_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6479_ _7950_/Q _6464_/X _6474_/X _6478_/X _6472_/X vssd1 vssd1 vccd1 vccd1 _7950_/D
+ sky130_fd_sc_hd__a221o_1
X_8218_ _8218_/CLK _8218_/D vssd1 vssd1 vccd1 vccd1 _8218_/Q sky130_fd_sc_hd__dfxtp_1
X_7005__425 _7005__425/A vssd1 vssd1 vccd1 vccd1 _8231_/CLK sky130_fd_sc_hd__inv_2
X_8149_ _8149_/CLK _8149_/D vssd1 vssd1 vccd1 vccd1 _8149_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_0 _7903_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3476_ clkbuf_0__3476_/X vssd1 vssd1 vccd1 vccd1 _7208__84/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7012__429 _7013__430/A vssd1 vssd1 vccd1 vccd1 _8235_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5850_ _4435_/X _7917_/Q _5854_/S vssd1 vssd1 vccd1 vccd1 _5851_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4801_ _4799_/X _4800_/X _4801_/S vssd1 vssd1 vccd1 vccd1 _4801_/X sky130_fd_sc_hd__mux2_1
X_5781_ _5781_/A vssd1 vssd1 vccd1 vccd1 _7996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4732_ _8334_/Q _8119_/Q _8071_/Q _8023_/Q _4731_/X _4702_/A vssd1 vssd1 vccd1 vccd1
+ _4732_/X sky130_fd_sc_hd__mux4_1
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _8271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6932__383 _6932__383/A vssd1 vssd1 vccd1 vccd1 _8179_/CLK sky130_fd_sc_hd__inv_2
X_6402_ _8631_/Q vssd1 vssd1 vccd1 vccd1 _6872_/A sky130_fd_sc_hd__buf_4
X_4594_ _4594_/A vssd1 vssd1 vccd1 vccd1 _8302_/D sky130_fd_sc_hd__clkbuf_1
X_7382_ _8434_/Q _7368_/X _7376_/X _7281_/X vssd1 vssd1 vccd1 vccd1 _7383_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6264_ _6257_/X _8092_/Q _6261_/X _6263_/X _7881_/Q vssd1 vssd1 vccd1 vccd1 _7881_/D
+ sky130_fd_sc_hd__o32a_1
X_8003_ _8003_/CLK _8003_/D vssd1 vssd1 vccd1 vccd1 _8003_/Q sky130_fd_sc_hd__dfxtp_1
X_5215_ _3965_/X _5078_/X _5214_/X _5152_/X vssd1 vssd1 vccd1 vccd1 _8211_/D sky130_fd_sc_hd__o211a_1
X_6195_ _6300_/A _6195_/B _6195_/C vssd1 vssd1 vccd1 vccd1 _6196_/A sky130_fd_sc_hd__and3_1
X_5146_ _5087_/X _5116_/X _5128_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5146_/X sky130_fd_sc_hd__a31o_2
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5077_ _5147_/A _7410_/A vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__nand2_1
X_7209__85 _7209__85/A vssd1 vssd1 vccd1 vccd1 _8394_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4028_ _4573_/A _5844_/B vssd1 vssd1 vccd1 vccd1 _4044_/S sky130_fd_sc_hd__or2_2
X_6642__284 _6643__285/A vssd1 vssd1 vccd1 vccd1 _8044_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ _5979_/A vssd1 vssd1 vccd1 vccd1 _5979_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7718_ _7778_/A vssd1 vssd1 vccd1 vccd1 _7723_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7649_ _7648_/X _7649_/B vssd1 vssd1 vccd1 vccd1 _7650_/A sky130_fd_sc_hd__and2b_1
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3459_ clkbuf_0__3459_/X vssd1 vssd1 vccd1 vccd1 _7124__517/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6585__238 _6585__238/A vssd1 vssd1 vccd1 vccd1 _7998_/CLK sky130_fd_sc_hd__inv_2
X_5000_ _5000_/A _5772_/A vssd1 vssd1 vccd1 vccd1 _5016_/S sky130_fd_sc_hd__nor2_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6951_ _6951_/A vssd1 vssd1 vccd1 vccd1 _8191_/D sky130_fd_sc_hd__clkbuf_1
X_5902_ _4194_/X _7851_/Q _5908_/S vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3663_ clkbuf_0__3663_/X vssd1 vssd1 vccd1 vccd1 _7747_/A sky130_fd_sc_hd__clkbuf_4
X_6882_ _8547_/Q _6886_/B vssd1 vssd1 vccd1 vccd1 _7564_/B sky130_fd_sc_hd__xnor2_4
X_5833_ _5833_/A vssd1 vssd1 vccd1 vccd1 _7925_/D sky130_fd_sc_hd__clkbuf_1
X_8621_ _8623_/CLK _8621_/D vssd1 vssd1 vccd1 vccd1 _8621_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8552_ _8553_/CLK _8552_/D vssd1 vssd1 vccd1 vccd1 _8552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5764_ _8003_/Q _5633_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__mux2_1
X_4715_ _8460_/Q _8350_/Q _8063_/Q _8484_/Q _4700_/X _4714_/X vssd1 vssd1 vccd1 vccd1
+ _4715_/X sky130_fd_sc_hd__mux4_1
X_8483_ _8483_/CLK _8483_/D vssd1 vssd1 vccd1 vccd1 _8483_/Q sky130_fd_sc_hd__dfxtp_1
X_5695_ _5695_/A vssd1 vssd1 vccd1 vccd1 _8034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4646_ _4646_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _4662_/S sky130_fd_sc_hd__nor2_2
X_4577_ _4432_/X _8309_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4578_/A sky130_fd_sc_hd__mux2_1
X_7365_ _7371_/A _7365_/B vssd1 vssd1 vccd1 vccd1 _8428_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6787__342 _6788__343/A vssd1 vssd1 vccd1 vccd1 _8134_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _7840_/A _4164_/X _6390_/A vssd1 vssd1 vccd1 vccd1 _7387_/A sky130_fd_sc_hd__a21o_1
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7296_ _8624_/Q _7281_/X _7331_/C _7330_/C _7331_/D vssd1 vssd1 vccd1 vccd1 _7297_/D
+ sky130_fd_sc_hd__o2111a_1
X_6247_ _6247_/A vssd1 vssd1 vccd1 vccd1 _6247_/X sky130_fd_sc_hd__clkbuf_2
X_6178_ _6178_/A _6186_/B vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__and2_1
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5209_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3313_ clkbuf_0__3313_/X vssd1 vssd1 vccd1 vccd1 _6790__345/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6939__389 _6940__390/A vssd1 vssd1 vccd1 vccd1 _8185_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7491__160 _7491__160/A vssd1 vssd1 vccd1 vccd1 _8499_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5480_ _5480_/A vssd1 vssd1 vccd1 vccd1 _8157_/D sky130_fd_sc_hd__clkbuf_1
X_4500_ _4500_/A vssd1 vssd1 vccd1 vccd1 _8337_/D sky130_fd_sc_hd__clkbuf_1
X_4431_ _4431_/A vssd1 vssd1 vccd1 vccd1 _8358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4362_ _4362_/A vssd1 vssd1 vccd1 vccd1 _8388_/D sky130_fd_sc_hd__clkbuf_1
X_7500__167 _7502__169/A vssd1 vssd1 vccd1 vccd1 _8506_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4293_ _8419_/Q _4206_/X _4297_/S vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__mux2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6101_/A vssd1 vssd1 vccd1 vccd1 _6101_/X sky130_fd_sc_hd__clkbuf_2
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6032_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6033_/A sky130_fd_sc_hd__and2_1
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7983_ _8441_/CLK _7983_/D vssd1 vssd1 vccd1 vccd1 _7983_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3646_ clkbuf_0__3646_/X vssd1 vssd1 vccd1 vccd1 _7453__129/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _7584_/A _7584_/B _6864_/Y vssd1 vssd1 vccd1 vccd1 _6865_/X sky130_fd_sc_hd__a21o_1
X_8604_ _8604_/CLK _8604_/D vssd1 vssd1 vccd1 vccd1 _8604_/Q sky130_fd_sc_hd__dfxtp_1
X_5816_ _5604_/X _7932_/Q _5818_/S vssd1 vssd1 vccd1 vccd1 _5817_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5747_ _5747_/A vssd1 vssd1 vccd1 vccd1 _8011_/D sky130_fd_sc_hd__clkbuf_1
X_8535_ _8535_/CLK _8535_/D vssd1 vssd1 vccd1 vccd1 _8535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8466_ _8466_/CLK _8466_/D vssd1 vssd1 vccd1 vccd1 _8466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _5613_/X _8041_/Q _5680_/S vssd1 vssd1 vccd1 vccd1 _5679_/A sky130_fd_sc_hd__mux2_1
X_7417_ _8445_/Q _7424_/B vssd1 vssd1 vccd1 vccd1 _7417_/X sky130_fd_sc_hd__or2_1
X_8397_ _8397_/CLK _8397_/D vssd1 vssd1 vccd1 vccd1 _8397_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3476_ _7204_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3476_/X sky130_fd_sc_hd__clkbuf_16
X_4629_ _4644_/S vssd1 vssd1 vccd1 vccd1 _4638_/S sky130_fd_sc_hd__buf_2
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7348_ _8416_/Q _8415_/Q vssd1 vssd1 vccd1 vccd1 _7349_/B sky130_fd_sc_hd__or2_1
XFILLER_104_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7279_ _8434_/Q vssd1 vssd1 vccd1 vccd1 _7279_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8651__216 vssd1 vssd1 vccd1 vccd1 _8651__216/HI core0Index[3] sky130_fd_sc_hd__conb_1
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4980_ _5055_/C _4984_/A vssd1 vssd1 vccd1 vccd1 _4980_/Y sky130_fd_sc_hd__nor2_1
X_3931_ _8576_/Q vssd1 vssd1 vccd1 vccd1 _3931_/X sky130_fd_sc_hd__buf_4
XFILLER_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7188__68 _7188__68/A vssd1 vssd1 vccd1 vccd1 _8377_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6650_ _6650_/A vssd1 vssd1 vccd1 vccd1 _8048_/D sky130_fd_sc_hd__clkbuf_1
X_5601_ _5601_/A vssd1 vssd1 vccd1 vccd1 _5601_/X sky130_fd_sc_hd__buf_2
X_5532_ _5532_/A vssd1 vssd1 vccd1 vccd1 _8131_/D sky130_fd_sc_hd__clkbuf_1
X_8320_ _8320_/CLK _8320_/D vssd1 vssd1 vccd1 vccd1 _8320_/Q sky130_fd_sc_hd__dfxtp_1
X_5463_ _5424_/X _8165_/Q _5465_/S vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8251_ _8251_/CLK _8251_/D vssd1 vssd1 vccd1 vccd1 _8251_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4414_ _4414_/A vssd1 vssd1 vccd1 vccd1 _8365_/D sky130_fd_sc_hd__clkbuf_1
X_8182_ _8182_/CLK _8182_/D vssd1 vssd1 vccd1 vccd1 _8182_/Q sky130_fd_sc_hd__dfxtp_1
X_5394_ _5101_/X _5385_/X _5393_/Y _5374_/X vssd1 vssd1 vccd1 vccd1 _8197_/D sky130_fd_sc_hd__o211a_1
X_7107__503 _7109__505/A vssd1 vssd1 vccd1 vccd1 _8312_/CLK sky130_fd_sc_hd__inv_2
X_4345_ _4119_/X _8395_/Q _4347_/S vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4276_ _8454_/Q _4209_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__mux2_1
X_6015_ _6015_/A vssd1 vssd1 vccd1 vccd1 _6015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6344__213 _6346__215/A vssd1 vssd1 vccd1 vccd1 _7925_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _8570_/CLK _7966_/D vssd1 vssd1 vccd1 vccd1 _7966_/Q sky130_fd_sc_hd__dfxtp_1
X_7897_ _8436_/CLK _7897_/D vssd1 vssd1 vccd1 vccd1 _7897_/Q sky130_fd_sc_hd__dfxtp_1
X_6848_ _6886_/A _6842_/C _6886_/C _8553_/Q vssd1 vssd1 vccd1 vccd1 _7555_/C sky130_fd_sc_hd__a31o_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6779_ _6785_/A vssd1 vssd1 vccd1 vccd1 _6779_/X sky130_fd_sc_hd__buf_1
X_8518_ _8518_/CLK _8518_/D vssd1 vssd1 vccd1 vccd1 _8518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8449_ _8604_/CLK _8449_/D vssd1 vssd1 vccd1 vccd1 _8449_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3459_ _7122_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3459_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7093__492 _7094__493/A vssd1 vssd1 vccd1 vccd1 _8301_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8568_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4130_ _8571_/Q vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ _4061_/A vssd1 vssd1 vccd1 vccd1 _8518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7820_ _8144_/Q _7820_/B vssd1 vssd1 vccd1 vccd1 _7842_/C sky130_fd_sc_hd__and2_1
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _4981_/A vssd1 vssd1 vccd1 vccd1 _7053_/C sky130_fd_sc_hd__clkbuf_2
X_6702_ _7812_/A _8082_/Q _6706_/S vssd1 vssd1 vccd1 vccd1 _6703_/A sky130_fd_sc_hd__mux2_1
X_7682_ _7682_/A _7682_/B _7681_/X vssd1 vssd1 vccd1 vccd1 _7682_/X sky130_fd_sc_hd__or3b_1
X_3914_ _6454_/A _6368_/A vssd1 vssd1 vccd1 vccd1 _6361_/A sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__3414_ clkbuf_0__3414_/X vssd1 vssd1 vccd1 vccd1 _6940__390/A sky130_fd_sc_hd__clkbuf_4
X_4894_ _4874_/X _8106_/Q _8002_/Q _4847_/X _4809_/A vssd1 vssd1 vccd1 vccd1 _4894_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6564_ _6564_/A vssd1 vssd1 vccd1 vccd1 _7982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5515_ _8138_/Q _4498_/X _5519_/S vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3276_ clkbuf_0__3276_/X vssd1 vssd1 vccd1 vccd1 _6695__311/A sky130_fd_sc_hd__clkbuf_4
X_8303_ _8303_/CLK _8303_/D vssd1 vssd1 vccd1 vccd1 _8303_/Q sky130_fd_sc_hd__dfxtp_1
X_6495_ _7956_/Q _6483_/X _6452_/A _6494_/X _6472_/A vssd1 vssd1 vccd1 vccd1 _7956_/D
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_0__3313_ _6785_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3313_/X sky130_fd_sc_hd__clkbuf_16
X_5446_ _5446_/A vssd1 vssd1 vccd1 vccd1 _8173_/D sky130_fd_sc_hd__clkbuf_1
X_8234_ _8234_/CLK _8234_/D vssd1 vssd1 vccd1 vccd1 _8234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8165_ _8165_/CLK _8165_/D vssd1 vssd1 vccd1 vccd1 _8165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5377_ _5377_/A _5377_/B _5377_/C vssd1 vssd1 vccd1 vccd1 _5378_/A sky130_fd_sc_hd__and3_1
X_4328_ _8402_/Q _4229_/X _4328_/S vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7116_ _7122_/A vssd1 vssd1 vccd1 vccd1 _7116_/X sky130_fd_sc_hd__buf_1
X_8096_ _8569_/CLK _8096_/D vssd1 vssd1 vccd1 vccd1 _8096_/Q sky130_fd_sc_hd__dfxtp_1
X_4259_ _4259_/A vssd1 vssd1 vccd1 vccd1 _4970_/B sky130_fd_sc_hd__inv_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6606__255 _6606__255/A vssd1 vssd1 vccd1 vccd1 _8015_/CLK sky130_fd_sc_hd__inv_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _8622_/CLK _7949_/D vssd1 vssd1 vccd1 vccd1 _7949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6687__305 _6687__305/A vssd1 vssd1 vccd1 vccd1 _8073_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8657__222 vssd1 vssd1 vccd1 vccd1 _8657__222/HI core1Index[2] sky130_fd_sc_hd__conb_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _5351_/A _5289_/X _5292_/X _5299_/X _5087_/A vssd1 vssd1 vccd1 vccd1 _5300_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6280_ _6280_/A _6306_/B vssd1 vssd1 vccd1 vccd1 _6732_/B sky130_fd_sc_hd__nor2_4
X_5231_ _8362_/Q _5220_/X _5305_/A _5227_/X _5230_/X vssd1 vssd1 vccd1 vccd1 _5231_/X
+ sky130_fd_sc_hd__o221a_1
X_5162_ _8507_/Q _8405_/Q _8142_/Q _8357_/Q _5169_/A _5140_/X vssd1 vssd1 vccd1 vccd1
+ _5162_/X sky130_fd_sc_hd__mux4_2
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6965__396 _6969__400/A vssd1 vssd1 vccd1 vccd1 _8200_/CLK sky130_fd_sc_hd__inv_2
X_4113_ _4113_/A vssd1 vssd1 vccd1 vccd1 _8499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6781__337 _6782__338/A vssd1 vssd1 vccd1 vccd1 _8129_/CLK sky130_fd_sc_hd__inv_2
X_5093_ _5239_/A vssd1 vssd1 vccd1 vccd1 _5246_/S sky130_fd_sc_hd__buf_2
XFILLER_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _3977_/X _8525_/Q _4044_/S vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7803_ _7803_/A _7812_/B vssd1 vssd1 vccd1 vccd1 _7803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5995_ _5995_/A vssd1 vssd1 vccd1 vccd1 _6004_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _4946_/A _4946_/B _4946_/C vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__or3_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _4827_/X _4875_/X _4876_/X vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__o21a_1
X_7665_ _7681_/A _7688_/B _7664_/C vssd1 vssd1 vccd1 vccd1 _7677_/A sky130_fd_sc_hd__o21bai_1
X_7596_ _7580_/X _7683_/A _7596_/C vssd1 vssd1 vccd1 vccd1 _7597_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6547_ _6547_/A vssd1 vssd1 vccd1 vccd1 _7977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3259_ clkbuf_0__3259_/X vssd1 vssd1 vccd1 vccd1 _6643__285/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6478_ _7798_/A _6490_/B _6481_/C vssd1 vssd1 vccd1 vccd1 _6478_/X sky130_fd_sc_hd__and3_1
X_5429_ _5428_/X _8180_/Q _5429_/S vssd1 vssd1 vccd1 vccd1 _5430_/A sky130_fd_sc_hd__mux2_1
X_8217_ _8217_/CLK _8217_/D vssd1 vssd1 vccd1 vccd1 _8217_/Q sky130_fd_sc_hd__dfxtp_1
X_8148_ _8148_/CLK _8148_/D vssd1 vssd1 vccd1 vccd1 _8148_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_1 _7903_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8079_ _8079_/CLK _8079_/D vssd1 vssd1 vccd1 vccd1 _8079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3475_ clkbuf_0__3475_/X vssd1 vssd1 vccd1 vccd1 _7200__77/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990__412 _6991__413/A vssd1 vssd1 vccd1 vccd1 _8218_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4800_ _8229_/Q _8184_/Q _8076_/Q _8421_/Q _4731_/X _4702_/A vssd1 vssd1 vccd1 vccd1
+ _4800_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5780_ _7996_/Q _5604_/A _5782_/S vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4731_ _4806_/B vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__buf_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4662_ _8271_/Q _4504_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6401_ _7937_/Q _6359_/X _6400_/Y _6391_/X vssd1 vssd1 vccd1 vccd1 _7937_/D sky130_fd_sc_hd__a211o_1
X_4593_ _4453_/X _8302_/Q _4601_/S vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__mux2_1
X_7381_ _7386_/A _7381_/B vssd1 vssd1 vccd1 vccd1 _8433_/D sky130_fd_sc_hd__nor2_1
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6263_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8002_ _8002_/CLK _8002_/D vssd1 vssd1 vccd1 vccd1 _8002_/Q sky130_fd_sc_hd__dfxtp_1
X_5214_ _8211_/Q _5080_/X _5385_/A _5213_/X _5148_/X vssd1 vssd1 vccd1 vccd1 _5214_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6194_ _6280_/A vssd1 vssd1 vccd1 vccd1 _6300_/A sky130_fd_sc_hd__inv_2
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5145_ _5133_/X _5137_/X _5142_/X _5247_/A _5217_/A vssd1 vssd1 vccd1 vccd1 _5145_/X
+ sky130_fd_sc_hd__o221a_1
X_5076_ _6986_/C vssd1 vssd1 vccd1 vccd1 _7410_/A sky130_fd_sc_hd__clkinv_2
Xclkbuf_1_0_0__3260_ clkbuf_0__3260_/X vssd1 vssd1 vccd1 vccd1 _6667__290/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _4336_/B _4027_/B _4336_/A vssd1 vssd1 vccd1 vccd1 _5844_/B sky130_fd_sc_hd__or3b_2
XFILLER_71_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5978_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__or2_1
XFILLER_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4924_/X _4925_/X _4928_/X _4992_/B vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__a211o_1
X_7717_ _7717_/A vssd1 vssd1 vccd1 vccd1 _8574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7648_ _7646_/Y _7642_/X _7647_/X _7589_/B vssd1 vssd1 vccd1 vccd1 _7648_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7579_ _7579_/A vssd1 vssd1 vccd1 vccd1 _7664_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3458_ clkbuf_0__3458_/X vssd1 vssd1 vccd1 vccd1 _7119__513/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6997__418 _6997__418/A vssd1 vssd1 vccd1 vccd1 _8224_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6950_ _8565_/Q _6958_/B vssd1 vssd1 vccd1 vccd1 _6951_/A sky130_fd_sc_hd__and2_1
X_5901_ _5901_/A vssd1 vssd1 vccd1 vccd1 _7852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3662_ clkbuf_0__3662_/X vssd1 vssd1 vccd1 vccd1 _7540__25/A sky130_fd_sc_hd__clkbuf_4
X_6881_ _7834_/A _7563_/B vssd1 vssd1 vccd1 vccd1 _6881_/X sky130_fd_sc_hd__xor2_1
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5832_ _7925_/Q _4435_/A _5836_/S vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__mux2_1
X_8620_ _8622_/CLK _8620_/D vssd1 vssd1 vccd1 vccd1 _8620_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5763_ _5763_/A vssd1 vssd1 vccd1 vccd1 _8004_/D sky130_fd_sc_hd__clkbuf_1
X_8551_ _8554_/CLK _8551_/D vssd1 vssd1 vccd1 vccd1 _8551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4714_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4714_/X sky130_fd_sc_hd__buf_2
X_8482_ _8482_/CLK _8482_/D vssd1 vssd1 vccd1 vccd1 _8482_/Q sky130_fd_sc_hd__dfxtp_1
X_5694_ _8034_/Q _5636_/X _5698_/S vssd1 vssd1 vccd1 vccd1 _5695_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4645_ _4645_/A vssd1 vssd1 vccd1 vccd1 _8279_/D sky130_fd_sc_hd__clkbuf_1
X_7433_ _7433_/A vssd1 vssd1 vccd1 vccd1 _8452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4576_ _4576_/A vssd1 vssd1 vccd1 vccd1 _8310_/D sky130_fd_sc_hd__clkbuf_1
X_7364_ _8428_/Q _7352_/X _7360_/X _7286_/B vssd1 vssd1 vccd1 vccd1 _7365_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_115_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6315_ _8416_/Q _8415_/Q vssd1 vssd1 vccd1 vccd1 _7358_/A sky130_fd_sc_hd__nor2_2
X_7295_ _7288_/X _7289_/Y _7292_/Y _7293_/Y _7294_/X vssd1 vssd1 vccd1 vccd1 _7331_/D
+ sky130_fd_sc_hd__o2111a_1
X_6246_ _6240_/X _8081_/Q _6245_/X _6238_/X _7870_/Q vssd1 vssd1 vccd1 vccd1 _7870_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6177_ _6177_/A vssd1 vssd1 vccd1 vccd1 _6186_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_97_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5128_ _5095_/X _5119_/X _5127_/X vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3312_ clkbuf_0__3312_/X vssd1 vssd1 vccd1 vccd1 _6782__338/A sky130_fd_sc_hd__clkbuf_4
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _8224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7156__543 _7157__544/A vssd1 vssd1 vccd1 vccd1 _8352_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7748__46 _7751__49/A vssd1 vssd1 vccd1 vccd1 _8597_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7057__463 _7058__464/A vssd1 vssd1 vccd1 vccd1 _8272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6591__243 _6591__243/A vssd1 vssd1 vccd1 vccd1 _8003_/CLK sky130_fd_sc_hd__inv_2
X_4430_ _4427_/X _8358_/Q _4442_/S vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4115_/X _8388_/Q _4365_/S vssd1 vssd1 vccd1 vccd1 _4362_/A sky130_fd_sc_hd__mux2_1
X_6100_ _7866_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__or2_1
XFILLER_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4292_ _4292_/A vssd1 vssd1 vccd1 vccd1 _8420_/D sky130_fd_sc_hd__clkbuf_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7982_ _8612_/CLK _7982_/D vssd1 vssd1 vccd1 vccd1 _7982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3645_ clkbuf_0__3645_/X vssd1 vssd1 vccd1 vccd1 _7467_/A sky130_fd_sc_hd__clkbuf_4
X_8637__253 vssd1 vssd1 vccd1 vccd1 partID[4] _8637__253/LO sky130_fd_sc_hd__conb_1
X_6864_ _8627_/Q _6864_/B vssd1 vssd1 vccd1 vccd1 _6864_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5815_ _5815_/A vssd1 vssd1 vccd1 vccd1 _7933_/D sky130_fd_sc_hd__clkbuf_1
X_7468__141 _7471__144/A vssd1 vssd1 vccd1 vccd1 _8480_/CLK sky130_fd_sc_hd__inv_2
X_8603_ _8612_/CLK _8603_/D vssd1 vssd1 vccd1 vccd1 _8603_/Q sky130_fd_sc_hd__dfxtp_1
X_5746_ _8011_/Q _5633_/X _5746_/S vssd1 vssd1 vccd1 vccd1 _5747_/A sky130_fd_sc_hd__mux2_1
X_8534_ _8534_/CLK _8534_/D vssd1 vssd1 vccd1 vccd1 _8534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8465_ _8465_/CLK _8465_/D vssd1 vssd1 vccd1 vccd1 _8465_/Q sky130_fd_sc_hd__dfxtp_1
X_5677_ _5677_/A vssd1 vssd1 vccd1 vccd1 _8042_/D sky130_fd_sc_hd__clkbuf_1
X_4628_ _5700_/A _5000_/A vssd1 vssd1 vccd1 vccd1 _4644_/S sky130_fd_sc_hd__or2_2
X_7416_ _8207_/Q _7756_/B _7413_/X _7415_/X _7336_/X vssd1 vssd1 vccd1 vccd1 _8444_/D
+ sky130_fd_sc_hd__o311a_1
X_8396_ _8396_/CLK _8396_/D vssd1 vssd1 vccd1 vccd1 _8396_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3475_ _7198_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3475_/X sky130_fd_sc_hd__clkbuf_16
X_4559_ _8317_/Q _4513_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__mux2_1
X_7278_ _7330_/A _7331_/A _7330_/B _7331_/B vssd1 vssd1 vccd1 vccd1 _7297_/C sky130_fd_sc_hd__and4_1
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6229_ _6247_/A vssd1 vssd1 vccd1 vccd1 _6229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3310_ clkbuf_0__3310_/X vssd1 vssd1 vccd1 vccd1 _6769__327/A sky130_fd_sc_hd__clkbuf_16
XFILLER_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _3930_/A vssd1 vssd1 vccd1 vccd1 _8601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5600_ _5600_/A vssd1 vssd1 vccd1 vccd1 _8078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5531_ _8131_/Q _4441_/A _5531_/S vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8250_ _8250_/CLK _8250_/D vssd1 vssd1 vccd1 vccd1 _8250_/Q sky130_fd_sc_hd__dfxtp_1
X_5462_ _5462_/A vssd1 vssd1 vccd1 vccd1 _8166_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3260_ _6644_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3260_/X sky130_fd_sc_hd__clkbuf_16
X_4413_ _4111_/X _8365_/Q _4419_/S vssd1 vssd1 vccd1 vccd1 _4414_/A sky130_fd_sc_hd__mux2_1
X_8181_ _8181_/CLK _8181_/D vssd1 vssd1 vccd1 vccd1 _8181_/Q sky130_fd_sc_hd__dfxtp_1
X_5393_ _5393_/A _5393_/B vssd1 vssd1 vccd1 vccd1 _5393_/Y sky130_fd_sc_hd__nand2_1
X_4344_ _4344_/A vssd1 vssd1 vccd1 vccd1 _8396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _6014_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _6015_/A sky130_fd_sc_hd__and2_1
XFILLER_100_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _4275_/A vssd1 vssd1 vccd1 vccd1 _8455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8674__239 vssd1 vssd1 vccd1 vccd1 _8674__239/HI partID[1] sky130_fd_sc_hd__conb_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7965_ _8570_/CLK _7965_/D vssd1 vssd1 vccd1 vccd1 _7965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6916_ _6916_/A vssd1 vssd1 vccd1 vccd1 _6916_/X sky130_fd_sc_hd__buf_1
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6598__249 _6599__250/A vssd1 vssd1 vccd1 vccd1 _8009_/CLK sky130_fd_sc_hd__inv_2
X_7896_ _8436_/CLK _7896_/D vssd1 vssd1 vccd1 vccd1 _7896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6847_ _6847_/A _7586_/A _6847_/C vssd1 vssd1 vccd1 vccd1 _6909_/A sky130_fd_sc_hd__and3_1
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5729_ _5729_/A vssd1 vssd1 vccd1 vccd1 _8019_/D sky130_fd_sc_hd__clkbuf_1
X_8517_ _8517_/CLK _8517_/D vssd1 vssd1 vccd1 vccd1 _8517_/Q sky130_fd_sc_hd__dfxtp_1
X_8448_ _8604_/CLK _8448_/D vssd1 vssd1 vccd1 vccd1 _8448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8379_ _8379_/CLK _8379_/D vssd1 vssd1 vccd1 vccd1 _8379_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3458_ _7116_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3458_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7193__72 _7194__73/A vssd1 vssd1 vccd1 vccd1 _8381_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4060_ _3974_/X _8518_/Q _4062_/S vssd1 vssd1 vccd1 vccd1 _4061_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4962_ _4478_/X _4669_/A _4961_/X _4903_/X vssd1 vssd1 vccd1 vccd1 _8261_/D sky130_fd_sc_hd__o211a_1
X_4893_ _4996_/B _4891_/X _4892_/X vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__o21a_1
X_6701_ _6701_/A vssd1 vssd1 vccd1 vccd1 _8081_/D sky130_fd_sc_hd__clkbuf_1
X_7681_ _7681_/A _7681_/B _7681_/C vssd1 vssd1 vccd1 vccd1 _7681_/X sky130_fd_sc_hd__or3_1
X_3913_ _7981_/Q vssd1 vssd1 vccd1 vccd1 _6368_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1_0__3413_ clkbuf_0__3413_/X vssd1 vssd1 vccd1 vccd1 _6932__383/A sky130_fd_sc_hd__clkbuf_4
X_6632_ _6674_/A vssd1 vssd1 vccd1 vccd1 _6632_/X sky130_fd_sc_hd__buf_1
XFILLER_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6563_ _7760_/A _6563_/B _6563_/C _6563_/D vssd1 vssd1 vccd1 vccd1 _6564_/A sky130_fd_sc_hd__and4_1
Xclkbuf_1_1_0__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6693__310/A sky130_fd_sc_hd__clkbuf_4
X_5514_ _5514_/A vssd1 vssd1 vccd1 vccd1 _8139_/D sky130_fd_sc_hd__clkbuf_1
X_8302_ _8302_/CLK _8302_/D vssd1 vssd1 vccd1 vccd1 _8302_/Q sky130_fd_sc_hd__dfxtp_1
X_6494_ _8613_/Q _6494_/B _8146_/Q vssd1 vssd1 vccd1 vccd1 _6494_/X sky130_fd_sc_hd__and3_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3312_ _6779_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3312_/X sky130_fd_sc_hd__clkbuf_16
X_5445_ _5424_/X _8173_/Q _5447_/S vssd1 vssd1 vccd1 vccd1 _5446_/A sky130_fd_sc_hd__mux2_1
X_8233_ _8233_/CLK _8233_/D vssd1 vssd1 vccd1 vccd1 _8233_/Q sky130_fd_sc_hd__dfxtp_1
X_8164_ _8164_/CLK _8164_/D vssd1 vssd1 vccd1 vccd1 _8164_/Q sky130_fd_sc_hd__dfxtp_1
X_5376_ _5376_/A _5376_/B vssd1 vssd1 vccd1 vccd1 _5377_/C sky130_fd_sc_hd__or2_1
X_4327_ _4327_/A vssd1 vssd1 vccd1 vccd1 _8403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8095_ _8556_/CLK _8095_/D vssd1 vssd1 vccd1 vccd1 _8095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4258_ _4258_/A vssd1 vssd1 vccd1 vccd1 _8461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4189_ _5790_/A vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _8623_/CLK _7948_/D vssd1 vssd1 vccd1 vccd1 _7948_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7879_ _8630_/CLK _7879_/D vssd1 vssd1 vccd1 vccd1 _7879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5230_ _8589_/Q _5230_/B vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__or2_1
XFILLER_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5161_ _5095_/A _5158_/X _5160_/X vssd1 vssd1 vccd1 vccd1 _5161_/X sky130_fd_sc_hd__a21o_1
X_4112_ _4111_/X _8499_/Q _4124_/S vssd1 vssd1 vccd1 vccd1 _4113_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5092_ _5134_/A vssd1 vssd1 vccd1 vccd1 _5239_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4043_ _4043_/A vssd1 vssd1 vccd1 vccd1 _8526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5994_ _5994_/A vssd1 vssd1 vccd1 vccd1 _5994_/X sky130_fd_sc_hd__clkbuf_1
X_7802_ _8620_/Q _7811_/B vssd1 vssd1 vccd1 vccd1 _7802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4945_ _8016_/Q _4807_/A _4796_/A _4944_/X vssd1 vssd1 vccd1 vccd1 _4946_/C sky130_fd_sc_hd__o211a_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7037__450 _7037__450/A vssd1 vssd1 vccd1 vccd1 _8257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7150__538 _7152__540/A vssd1 vssd1 vccd1 vccd1 _8347_/CLK sky130_fd_sc_hd__inv_2
X_4876_ _8419_/Q _4855_/X _8227_/Q _4856_/X _4834_/X vssd1 vssd1 vccd1 vccd1 _4876_/X
+ sky130_fd_sc_hd__o221a_1
X_7664_ _8558_/Q _7664_/B _7664_/C vssd1 vssd1 vccd1 vccd1 _7664_/X sky130_fd_sc_hd__and3_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7595_ _7578_/X _7647_/A _7664_/C vssd1 vssd1 vccd1 vccd1 _7596_/C sky130_fd_sc_hd__a21o_1
X_6546_ _8092_/Q _7977_/Q _6548_/S vssd1 vssd1 vccd1 vccd1 _6547_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3258_ clkbuf_0__3258_/X vssd1 vssd1 vccd1 vccd1 _6636__279/A sky130_fd_sc_hd__clkbuf_4
X_6477_ _6494_/B vssd1 vssd1 vccd1 vccd1 _6490_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6612__260 _6612__260/A vssd1 vssd1 vccd1 vccd1 _8020_/CLK sky130_fd_sc_hd__inv_2
X_5428_ _5616_/A vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__clkbuf_2
X_8216_ _8604_/CLK _8216_/D vssd1 vssd1 vccd1 vccd1 _8216_/Q sky130_fd_sc_hd__dfxtp_1
X_8147_ _8147_/CLK _8147_/D vssd1 vssd1 vccd1 vccd1 _8147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5359_ _8517_/Q _5359_/B vssd1 vssd1 vccd1 vccd1 _5359_/X sky130_fd_sc_hd__or2_1
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8078_ _8078_/CLK _8078_/D vssd1 vssd1 vccd1 vccd1 _8078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_2 _3940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3474_ clkbuf_0__3474_/X vssd1 vssd1 vccd1 vccd1 _7210_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6693__310 _6693__310/A vssd1 vssd1 vccd1 vccd1 _8078_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _8232_/Q _8187_/Q _8079_/Q _8424_/Q _4710_/A _4729_/X vssd1 vssd1 vccd1 vccd1
+ _4730_/X sky130_fd_sc_hd__mux4_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ _4661_/A vssd1 vssd1 vccd1 vccd1 _8272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7462__136 _7463__137/A vssd1 vssd1 vccd1 vccd1 _8475_/CLK sky130_fd_sc_hd__inv_2
X_7380_ _8433_/Q _7368_/X _7376_/X _7379_/Y vssd1 vssd1 vccd1 vccd1 _7381_/B sky130_fd_sc_hd__o2bb2a_1
X_6400_ _6416_/A _6400_/B _6400_/C vssd1 vssd1 vccd1 vccd1 _6400_/Y sky130_fd_sc_hd__nor3_2
X_4592_ _4607_/S vssd1 vssd1 vccd1 vccd1 _4601_/S sky130_fd_sc_hd__buf_2
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6262_ _6257_/X _8091_/Q _6261_/X _6255_/X _7880_/Q vssd1 vssd1 vccd1 vccd1 _7880_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5213_ _5087_/X _5199_/X _5203_/X _5212_/X vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__a31o_2
X_8001_ _8001_/CLK _8001_/D vssd1 vssd1 vccd1 vccd1 _8001_/Q sky130_fd_sc_hd__dfxtp_1
X_6193_ _6193_/A vssd1 vssd1 vccd1 vccd1 _6280_/A sky130_fd_sc_hd__buf_2
XFILLER_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5144_ _8200_/Q _5144_/B vssd1 vssd1 vccd1 vccd1 _5217_/A sky130_fd_sc_hd__xnor2_4
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5075_/A _5075_/B _5074_/X vssd1 vssd1 vccd1 vccd1 _6986_/C sky130_fd_sc_hd__or3b_2
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4026_ _8204_/Q vssd1 vssd1 vccd1 vccd1 _4336_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _5977_/A vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _8173_/Q _4865_/X _4713_/A _4927_/X vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__o211a_1
X_7527__14 _7528__15/A vssd1 vssd1 vccd1 vccd1 _8528_/CLK sky130_fd_sc_hd__inv_2
X_7716_ _7716_/A _7716_/B _7723_/C vssd1 vssd1 vccd1 vccd1 _7717_/A sky130_fd_sc_hd__and3_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7647_ _7647_/A vssd1 vssd1 vccd1 vccd1 _7647_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4859_ _4844_/X _4851_/X _4683_/A _4858_/X vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7578_ _7681_/A _7681_/B _7575_/X _7642_/A _7577_/X vssd1 vssd1 vccd1 vccd1 _7578_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6529_ _6036_/A _7969_/Q _6537_/S vssd1 vssd1 vccd1 vccd1 _6530_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3457_ clkbuf_0__3457_/X vssd1 vssd1 vccd1 vccd1 _7115__510/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5900_ _4156_/X _7852_/Q _5908_/S vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3661_ clkbuf_0__3661_/X vssd1 vssd1 vccd1 vccd1 _7534__20/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6880_ _6891_/C _6880_/B vssd1 vssd1 vccd1 vccd1 _7563_/B sky130_fd_sc_hd__nand2_2
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5831_ _5831_/A vssd1 vssd1 vccd1 vccd1 _7926_/D sky130_fd_sc_hd__clkbuf_1
X_5762_ _8004_/Q _5630_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8550_ _8554_/CLK _8550_/D vssd1 vssd1 vccd1 vccd1 _8550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4713_ _4713_/A vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8481_ _8481_/CLK _8481_/D vssd1 vssd1 vccd1 vccd1 _8481_/Q sky130_fd_sc_hd__dfxtp_1
X_5693_ _5693_/A vssd1 vssd1 vccd1 vccd1 _8035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4644_ _4478_/X _8279_/Q _4644_/S vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__mux2_1
X_7432_ _8452_/Q _7413_/A _7432_/S vssd1 vssd1 vccd1 vccd1 _7433_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4575_ _4427_/X _8310_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__mux2_1
X_7363_ _7371_/A _7363_/B vssd1 vssd1 vccd1 vccd1 _8427_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7294_ _8633_/Q _7294_/B vssd1 vssd1 vccd1 vccd1 _7294_/X sky130_fd_sc_hd__or2_1
X_6314_ _8443_/Q _6310_/X _6312_/X _7318_/A vssd1 vssd1 vccd1 vccd1 _6314_/X sky130_fd_sc_hd__a211o_1
X_6245_ _6306_/A vssd1 vssd1 vccd1 vccd1 _6245_/X sky130_fd_sc_hd__clkbuf_2
X_6176_ _6176_/A vssd1 vssd1 vccd1 vccd1 _6176_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5127_ _5121_/X _5124_/X _5333_/A vssd1 vssd1 vccd1 vccd1 _5127_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3311_ clkbuf_0__3311_/X vssd1 vssd1 vccd1 vccd1 _6778__335/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5058_ _4453_/X _8224_/Q _5066_/S vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4009_ _8540_/Q _3872_/X _4017_/S vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6794__348 _6794__348/A vssd1 vssd1 vccd1 vccd1 _8140_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ _4360_/A vssd1 vssd1 vccd1 vccd1 _8389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4291_ _8420_/Q _4203_/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__mux2_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6030_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__and2_1
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7981_ _8570_/CLK _7981_/D vssd1 vssd1 vccd1 vccd1 _7981_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3644_ clkbuf_0__3644_/X vssd1 vssd1 vccd1 vccd1 _7443__121/A sky130_fd_sc_hd__clkbuf_4
X_6863_ _7566_/B _7566_/C vssd1 vssd1 vccd1 vccd1 _6864_/B sky130_fd_sc_hd__nand2_1
X_5814_ _5601_/X _7933_/Q _5818_/S vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__mux2_1
X_8602_ _8608_/CLK _8602_/D vssd1 vssd1 vccd1 vccd1 _8602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5745_ _5745_/A vssd1 vssd1 vccd1 vccd1 _8012_/D sky130_fd_sc_hd__clkbuf_1
X_8533_ _8533_/CLK _8533_/D vssd1 vssd1 vccd1 vccd1 _8533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8464_ _8464_/CLK _8464_/D vssd1 vssd1 vccd1 vccd1 _8464_/Q sky130_fd_sc_hd__dfxtp_1
X_5676_ _5610_/X _8042_/Q _5680_/S vssd1 vssd1 vccd1 vccd1 _5677_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3474_ _7197_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3474_/X sky130_fd_sc_hd__clkbuf_16
X_4627_ _5880_/A vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__buf_2
X_7415_ _8444_/Q _7424_/B vssd1 vssd1 vccd1 vccd1 _7415_/X sky130_fd_sc_hd__or2_1
X_8395_ _8395_/CLK _8395_/D vssd1 vssd1 vccd1 vccd1 _8395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4558_ _4558_/A vssd1 vssd1 vccd1 vccd1 _8318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4489_ _8575_/Q vssd1 vssd1 vccd1 vccd1 _4489_/X sky130_fd_sc_hd__buf_2
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7277_ _8628_/Q _7369_/A _7369_/B vssd1 vssd1 vccd1 vccd1 _7331_/B sky130_fd_sc_hd__nand3b_1
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6228_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__buf_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6175_/A vssd1 vssd1 vccd1 vccd1 _6159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6208__182 _6209__183/A vssd1 vssd1 vccd1 vccd1 _7851_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6818__362 _6819__363/A vssd1 vssd1 vccd1 vccd1 _8157_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5530_ _5530_/A vssd1 vssd1 vccd1 vccd1 _8132_/D sky130_fd_sc_hd__clkbuf_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7031__445 _7031__445/A vssd1 vssd1 vccd1 vccd1 _8252_/CLK sky130_fd_sc_hd__inv_2
X_5461_ _5420_/X _8166_/Q _5465_/S vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4412_ _4412_/A vssd1 vssd1 vccd1 vccd1 _8366_/D sky130_fd_sc_hd__clkbuf_1
X_8180_ _8180_/CLK _8180_/D vssd1 vssd1 vccd1 vccd1 _8180_/Q sky130_fd_sc_hd__dfxtp_1
X_5392_ _5236_/X _5385_/X _5391_/Y _5374_/X vssd1 vssd1 vccd1 vccd1 _8198_/D sky130_fd_sc_hd__o211a_1
X_4343_ _4115_/X _8396_/Q _4347_/S vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__mux2_1
X_4274_ _8455_/Q _4206_/X _4278_/S vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__mux2_1
X_6013_ _6013_/A vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7964_ _8570_/CLK _7964_/D vssd1 vssd1 vccd1 vccd1 _7964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7114__509 _7114__509/A vssd1 vssd1 vccd1 vccd1 _8318_/CLK sky130_fd_sc_hd__inv_2
X_7895_ _8436_/CLK _7895_/D vssd1 vssd1 vccd1 vccd1 _7895_/Q sky130_fd_sc_hd__dfxtp_1
X_6846_ _7798_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6847_/C sky130_fd_sc_hd__or2_1
XFILLER_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8516_ _8516_/CLK _8516_/D vssd1 vssd1 vccd1 vccd1 _8516_/Q sky130_fd_sc_hd__dfxtp_1
X_5728_ _8019_/Q _5633_/X _5728_/S vssd1 vssd1 vccd1 vccd1 _5729_/A sky130_fd_sc_hd__mux2_1
X_3989_ _3989_/A vssd1 vssd1 vccd1 vccd1 _8584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5659_ _5613_/X _8057_/Q _5661_/S vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__mux2_1
X_8447_ _8604_/CLK _8447_/D vssd1 vssd1 vccd1 vccd1 _8447_/Q sky130_fd_sc_hd__dfxtp_1
X_8378_ _8378_/CLK _8378_/D vssd1 vssd1 vccd1 vccd1 _8378_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3457_ _7110_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3457_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6351__219 _6351__219/A vssd1 vssd1 vccd1 vccd1 _7931_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7329_ _7394_/A _7394_/B _7798_/A vssd1 vssd1 vccd1 vccd1 _7329_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7513__2 _7513__2/A vssd1 vssd1 vccd1 vccd1 _8516_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8091_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _4672_/A _8261_/Q _4989_/A _4960_/X _4741_/A vssd1 vssd1 vccd1 vccd1 _4961_/X
+ sky130_fd_sc_hd__a221o_1
X_4892_ _8313_/Q _4815_/X _4838_/X _8297_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4892_/X
+ sky130_fd_sc_hd__o221a_1
X_6700_ _7815_/A _8081_/Q _6706_/S vssd1 vssd1 vccd1 vccd1 _6701_/A sky130_fd_sc_hd__mux2_1
X_7680_ _8560_/Q _7672_/A _8561_/Q vssd1 vssd1 vccd1 vccd1 _7681_/C sky130_fd_sc_hd__a21oi_1
XFILLER_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3912_ _7982_/Q vssd1 vssd1 vccd1 vccd1 _6454_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1_0__3412_ clkbuf_0__3412_/X vssd1 vssd1 vccd1 vccd1 _6928__380/A sky130_fd_sc_hd__clkbuf_4
X_6631_ _6631_/A vssd1 vssd1 vccd1 vccd1 _6631_/X sky130_fd_sc_hd__buf_1
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8301_ _8301_/CLK _8301_/D vssd1 vssd1 vccd1 vccd1 _8301_/Q sky130_fd_sc_hd__dfxtp_1
X_6751__313 _6753__315/A vssd1 vssd1 vccd1 vccd1 _8105_/CLK sky130_fd_sc_hd__inv_2
X_6562_ _6562_/A _6562_/B vssd1 vssd1 vccd1 vccd1 _6563_/D sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6685__303/A sky130_fd_sc_hd__clkbuf_4
X_5513_ _8139_/Q _4495_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__mux2_1
X_6493_ _7955_/Q _6483_/X _6452_/A _6492_/X _6472_/A vssd1 vssd1 vccd1 vccd1 _7955_/D
+ sky130_fd_sc_hd__a221o_1
X_8232_ _8232_/CLK _8232_/D vssd1 vssd1 vccd1 vccd1 _8232_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3311_ _6773_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3311_/X sky130_fd_sc_hd__clkbuf_16
X_5444_ _5444_/A vssd1 vssd1 vccd1 vccd1 _8174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8163_ _8554_/CLK _8163_/D vssd1 vssd1 vccd1 vccd1 _8163_/Q sky130_fd_sc_hd__dfxtp_1
X_5375_ _5373_/A _5377_/B _5373_/Y _5374_/X vssd1 vssd1 vccd1 vccd1 _8204_/D sky130_fd_sc_hd__o211a_1
X_4326_ _8403_/Q _4226_/X _4328_/S vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8094_ _8270_/CLK _8094_/D vssd1 vssd1 vccd1 vccd1 _8094_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_113_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4257_ _8461_/Q _4238_/X _4257_/S vssd1 vssd1 vccd1 vccd1 _4258_/A sky130_fd_sc_hd__mux2_1
X_7045_ _7051_/A vssd1 vssd1 vccd1 vccd1 _7045_/X sky130_fd_sc_hd__buf_1
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4188_ _4454_/A _4985_/A _4970_/C vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__or3_4
XFILLER_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7947_ _8622_/CLK _7947_/D vssd1 vssd1 vccd1 vccd1 _7947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _8622_/CLK _7878_/D vssd1 vssd1 vccd1 vccd1 _7878_/Q sky130_fd_sc_hd__dfxtp_1
X_6829_ _8546_/Q _8545_/Q _8544_/Q _8543_/Q vssd1 vssd1 vccd1 vccd1 _6850_/A sky130_fd_sc_hd__and4_2
XFILLER_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5160_ _5121_/X _5159_/X _5344_/A vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4111_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__buf_2
X_5091_ _5112_/B _5103_/B vssd1 vssd1 vccd1 vccd1 _5134_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4042_ _3974_/X _8526_/Q _4044_/S vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7801_ _7798_/Y _7799_/Y _7800_/X vssd1 vssd1 vccd1 vccd1 _8619_/D sky130_fd_sc_hd__a21oi_1
X_5993_ _5993_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__or2_4
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4944_ _8327_/Q _4817_/A _4861_/A _4943_/X vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4875_ _4874_/X _8182_/Q _8074_/Q _4853_/X vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__a22o_1
X_7663_ _7663_/A vssd1 vssd1 vccd1 vccd1 _8557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7594_ _7581_/X _7573_/X _7688_/B _7681_/A vssd1 vssd1 vccd1 vccd1 _7647_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6545_ _6545_/A vssd1 vssd1 vccd1 vccd1 _7976_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3257_ clkbuf_0__3257_/X vssd1 vssd1 vccd1 vccd1 _6674_/A sky130_fd_sc_hd__clkbuf_4
X_6476_ _7588_/A vssd1 vssd1 vccd1 vccd1 _7798_/A sky130_fd_sc_hd__clkbuf_4
X_8215_ _8570_/CLK _8215_/D vssd1 vssd1 vccd1 vccd1 _8215_/Q sky130_fd_sc_hd__dfxtp_1
X_5427_ _8188_/Q vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _7912_/Q _8509_/Q _5358_/S vssd1 vssd1 vccd1 vccd1 _5358_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8146_ _8617_/CLK _8146_/D vssd1 vssd1 vccd1 vccd1 _8146_/Q sky130_fd_sc_hd__dfxtp_1
X_7044__455 _7044__455/A vssd1 vssd1 vccd1 vccd1 _8262_/CLK sky130_fd_sc_hd__inv_2
X_8077_ _8077_/CLK _8077_/D vssd1 vssd1 vccd1 vccd1 _8077_/Q sky130_fd_sc_hd__dfxtp_1
X_4309_ _4309_/A vssd1 vssd1 vccd1 vccd1 _8411_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_3 _4156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5289_ _5269_/X _5287_/X _5288_/X _5209_/A vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__o211a_1
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3473_ clkbuf_0__3473_/X vssd1 vssd1 vccd1 vccd1 _7196__75/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6758__319 _6758__319/A vssd1 vssd1 vccd1 vccd1 _8111_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3809_ clkbuf_0__3809_/X vssd1 vssd1 vccd1 vccd1 _7734__35/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4660_ _8272_/Q _4501_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4591_ _5862_/A _5000_/A vssd1 vssd1 vccd1 vccd1 _4607_/S sky130_fd_sc_hd__or2_2
XFILLER_115_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6261_ _6306_/A vssd1 vssd1 vccd1 vccd1 _6261_/X sky130_fd_sc_hd__clkbuf_2
X_5212_ _5351_/A _5207_/X _5209_/X _5211_/X _5217_/A vssd1 vssd1 vccd1 vccd1 _5212_/X
+ sky130_fd_sc_hd__o221a_1
X_8000_ _8000_/CLK _8000_/D vssd1 vssd1 vccd1 vccd1 _8000_/Q sky130_fd_sc_hd__dfxtp_1
X_6192_ _6088_/B _7983_/Q _6190_/X _6191_/X _6101_/A vssd1 vssd1 vccd1 vccd1 _6192_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5143_ _5204_/A vssd1 vssd1 vccd1 vccd1 _5247_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5074_ _5074_/A _5074_/B _5074_/C _5074_/D vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__and4_1
XFILLER_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4025_ _5467_/A vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__buf_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ _5976_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5977_/A sky130_fd_sc_hd__or2_1
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4927_ _8234_/Q _4821_/A _4926_/X _4861_/A vssd1 vssd1 vccd1 vccd1 _4927_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7715_ _7715_/A vssd1 vssd1 vccd1 vccd1 _8573_/D sky130_fd_sc_hd__clkbuf_1
X_4858_ _4845_/X _4854_/X _4857_/X vssd1 vssd1 vccd1 vccd1 _4858_/X sky130_fd_sc_hd__o21a_1
X_7646_ _8553_/Q vssd1 vssd1 vccd1 vccd1 _7646_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3309_ clkbuf_0__3309_/X vssd1 vssd1 vccd1 vccd1 _6791_/A sky130_fd_sc_hd__clkbuf_4
X_4789_ _4758_/X _4788_/X _4946_/A vssd1 vssd1 vccd1 vccd1 _4789_/X sky130_fd_sc_hd__a21o_1
X_7577_ _7581_/A _7579_/A _7575_/X vssd1 vssd1 vccd1 vccd1 _7577_/X sky130_fd_sc_hd__or3b_1
X_6202__177 _6204__179/A vssd1 vssd1 vccd1 vccd1 _7846_/CLK sky130_fd_sc_hd__inv_2
X_8647__212 vssd1 vssd1 vccd1 vccd1 _8647__212/HI caravel_irq[3] sky130_fd_sc_hd__conb_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _6550_/A vssd1 vssd1 vccd1 vccd1 _6537_/S sky130_fd_sc_hd__buf_2
XFILLER_109_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6459_ _6472_/A vssd1 vssd1 vccd1 vccd1 _6459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8129_ _8129_/CLK _8129_/D vssd1 vssd1 vccd1 vccd1 _8129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3456_ clkbuf_0__3456_/X vssd1 vssd1 vccd1 vccd1 _7109__505/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7231__102 _7231__102/A vssd1 vssd1 vccd1 vccd1 _8411_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6812__357 _6813__358/A vssd1 vssd1 vccd1 vccd1 _8152_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3660_ clkbuf_0__3660_/X vssd1 vssd1 vccd1 vccd1 _7526__13/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5830_ _7926_/Q _4432_/A _5836_/S vssd1 vssd1 vccd1 vccd1 _5831_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5761_ _5761_/A vssd1 vssd1 vccd1 vccd1 _8005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8480_ _8480_/CLK _8480_/D vssd1 vssd1 vccd1 vccd1 _8480_/Q sky130_fd_sc_hd__dfxtp_1
X_4712_ _4733_/A vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__clkbuf_4
X_5692_ _8035_/Q _5633_/X _5692_/S vssd1 vssd1 vccd1 vccd1 _5693_/A sky130_fd_sc_hd__mux2_1
X_7431_ _8214_/Q _7411_/A _7413_/A _7430_/X _7420_/A vssd1 vssd1 vccd1 vccd1 _8451_/D
+ sky130_fd_sc_hd__o311a_1
X_4643_ _4643_/A vssd1 vssd1 vccd1 vccd1 _8280_/D sky130_fd_sc_hd__clkbuf_1
X_4574_ _4589_/S vssd1 vssd1 vccd1 vccd1 _4583_/S sky130_fd_sc_hd__clkbuf_4
X_7362_ _8427_/Q _7352_/X _7360_/X _7361_/Y vssd1 vssd1 vccd1 vccd1 _7363_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7293_ _8633_/Q _7294_/B vssd1 vssd1 vccd1 vccd1 _7293_/Y sky130_fd_sc_hd__nand2_1
X_6313_ _8415_/Q vssd1 vssd1 vccd1 vccd1 _7318_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6244_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6306_/A sky130_fd_sc_hd__buf_4
X_6175_ _6175_/A vssd1 vssd1 vccd1 vccd1 _6175_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5126_ _5204_/A vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5057_ _5072_/S vssd1 vssd1 vccd1 vccd1 _5066_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4008_ _4023_/S vssd1 vssd1 vccd1 vccd1 _4017_/S sky130_fd_sc_hd__buf_2
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7220__94 _7221__95/A vssd1 vssd1 vccd1 vccd1 _8403_/CLK sky130_fd_sc_hd__inv_2
X_6915__370 _6915__370/A vssd1 vssd1 vccd1 vccd1 _8166_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7629_ _7629_/A vssd1 vssd1 vccd1 vccd1 _8548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7163__549 _7164__550/A vssd1 vssd1 vccd1 vccd1 _8358_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3439_ clkbuf_0__3439_/X vssd1 vssd1 vccd1 vccd1 _7023__438/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4290_ _4290_/A vssd1 vssd1 vccd1 vccd1 _8421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7064__469 _7065__470/A vssd1 vssd1 vccd1 vccd1 _8278_/CLK sky130_fd_sc_hd__inv_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7980_ _8270_/CLK _7980_/D vssd1 vssd1 vccd1 vccd1 _7980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3643_ clkbuf_0__3643_/X vssd1 vssd1 vccd1 vccd1 _7441__120/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6862_ _6842_/C _6852_/B _8549_/Q vssd1 vssd1 vccd1 vccd1 _7566_/C sky130_fd_sc_hd__a21o_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8601_ _8601_/CLK _8601_/D vssd1 vssd1 vccd1 vccd1 _8601_/Q sky130_fd_sc_hd__dfxtp_1
X_5813_ _5813_/A vssd1 vssd1 vccd1 vccd1 _7934_/D sky130_fd_sc_hd__clkbuf_1
X_8532_ _8532_/CLK _8532_/D vssd1 vssd1 vccd1 vccd1 _8532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5744_ _8012_/Q _5630_/X _5746_/S vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__mux2_1
X_8463_ _8463_/CLK _8463_/D vssd1 vssd1 vccd1 vccd1 _8463_/Q sky130_fd_sc_hd__dfxtp_1
X_5675_ _5675_/A vssd1 vssd1 vccd1 vccd1 _8043_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3473_ _7191_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3473_/X sky130_fd_sc_hd__clkbuf_16
X_8394_ _8394_/CLK _8394_/D vssd1 vssd1 vccd1 vccd1 _8394_/Q sky130_fd_sc_hd__dfxtp_1
X_4626_ _4626_/A vssd1 vssd1 vccd1 vccd1 _8287_/D sky130_fd_sc_hd__clkbuf_1
X_7414_ _7430_/B vssd1 vssd1 vccd1 vccd1 _7424_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4557_ _8318_/Q _4507_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4488_ _4488_/A vssd1 vssd1 vccd1 vccd1 _8341_/D sky130_fd_sc_hd__clkbuf_1
X_7276_ _7369_/A _7369_/B _8628_/Q vssd1 vssd1 vccd1 vccd1 _7330_/B sky130_fd_sc_hd__a21bo_1
XFILLER_103_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6227_ _6280_/A _6306_/B vssd1 vssd1 vccd1 vccd1 _6272_/A sky130_fd_sc_hd__or2_4
X_6568__225 _6568__225/A vssd1 vssd1 vccd1 vccd1 _7985_/CLK sky130_fd_sc_hd__inv_2
X_7475__147 _7477__149/A vssd1 vssd1 vccd1 vccd1 _8486_/CLK sky130_fd_sc_hd__inv_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6136_/A _6155_/X _6156_/X _6157_/X vssd1 vssd1 vccd1 vccd1 _6158_/X sky130_fd_sc_hd__o211a_1
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5109_ _5221_/A vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__buf_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6073_/X _6087_/X _6088_/X _6082_/X vssd1 vssd1 vccd1 vccd1 _6089_/X sky130_fd_sc_hd__o211a_1
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3809_ _7729_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3809_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7727__29 _7728__30/A vssd1 vssd1 vccd1 vccd1 _8580_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5460_ _5460_/A vssd1 vssd1 vccd1 vccd1 _8167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4411_ _4104_/X _8366_/Q _4419_/S vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5391_ _5393_/A _5391_/B vssd1 vssd1 vccd1 vccd1 _5391_/Y sky130_fd_sc_hd__nand2_1
X_4342_ _4342_/A vssd1 vssd1 vccd1 vccd1 _8397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4273_ _4273_/A vssd1 vssd1 vccd1 vccd1 _8456_/D sky130_fd_sc_hd__clkbuf_1
X_6012_ _6012_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _6013_/A sky130_fd_sc_hd__and2_1
XFILLER_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
.ends

