// This is the unpowered netlist.
module WishboneInterconnect (master0_wb_ack_i,
    master0_wb_cyc_o,
    master0_wb_error_i,
    master0_wb_stall_i,
    master0_wb_stb_o,
    master0_wb_we_o,
    master1_wb_ack_i,
    master1_wb_cyc_o,
    master1_wb_error_i,
    master1_wb_stall_i,
    master1_wb_stb_o,
    master1_wb_we_o,
    master2_wb_ack_i,
    master2_wb_cyc_o,
    master2_wb_error_i,
    master2_wb_stall_i,
    master2_wb_stb_o,
    master2_wb_we_o,
    slave0_wb_ack_o,
    slave0_wb_cyc_i,
    slave0_wb_error_o,
    slave0_wb_stall_o,
    slave0_wb_stb_i,
    slave0_wb_we_i,
    slave1_wb_ack_o,
    slave1_wb_cyc_i,
    slave1_wb_error_o,
    slave1_wb_stall_o,
    slave1_wb_stb_i,
    slave1_wb_we_i,
    slave2_wb_ack_o,
    slave2_wb_cyc_i,
    slave2_wb_error_o,
    slave2_wb_stall_o,
    slave2_wb_stb_i,
    slave2_wb_we_i,
    slave3_wb_ack_o,
    slave3_wb_cyc_i,
    slave3_wb_error_o,
    slave3_wb_stall_o,
    slave3_wb_stb_i,
    slave3_wb_we_i,
    slave4_wb_ack_o,
    slave4_wb_cyc_i,
    slave4_wb_error_o,
    slave4_wb_stall_o,
    slave4_wb_stb_i,
    slave4_wb_we_i,
    wb_clk_i,
    wb_rst_i,
    master0_wb_adr_o,
    master0_wb_data_i,
    master0_wb_data_o,
    master0_wb_sel_o,
    master1_wb_adr_o,
    master1_wb_data_i,
    master1_wb_data_o,
    master1_wb_sel_o,
    master2_wb_adr_o,
    master2_wb_data_i,
    master2_wb_data_o,
    master2_wb_sel_o,
    probe_master0_currentSlave,
    probe_master1_currentSlave,
    probe_master2_currentSlave,
    probe_master3_currentSlave,
    probe_slave0_currentMaster,
    probe_slave1_currentMaster,
    probe_slave2_currentMaster,
    probe_slave3_currentMaster,
    slave0_wb_adr_i,
    slave0_wb_data_i,
    slave0_wb_data_o,
    slave0_wb_sel_i,
    slave1_wb_adr_i,
    slave1_wb_data_i,
    slave1_wb_data_o,
    slave1_wb_sel_i,
    slave2_wb_adr_i,
    slave2_wb_data_i,
    slave2_wb_data_o,
    slave2_wb_sel_i,
    slave3_wb_adr_i,
    slave3_wb_data_i,
    slave3_wb_data_o,
    slave3_wb_sel_i,
    slave4_wb_adr_i,
    slave4_wb_data_i,
    slave4_wb_data_o,
    slave4_wb_sel_i);
 output master0_wb_ack_i;
 input master0_wb_cyc_o;
 output master0_wb_error_i;
 output master0_wb_stall_i;
 input master0_wb_stb_o;
 input master0_wb_we_o;
 output master1_wb_ack_i;
 input master1_wb_cyc_o;
 output master1_wb_error_i;
 output master1_wb_stall_i;
 input master1_wb_stb_o;
 input master1_wb_we_o;
 output master2_wb_ack_i;
 input master2_wb_cyc_o;
 output master2_wb_error_i;
 output master2_wb_stall_i;
 input master2_wb_stb_o;
 input master2_wb_we_o;
 input slave0_wb_ack_o;
 output slave0_wb_cyc_i;
 input slave0_wb_error_o;
 input slave0_wb_stall_o;
 output slave0_wb_stb_i;
 output slave0_wb_we_i;
 input slave1_wb_ack_o;
 output slave1_wb_cyc_i;
 input slave1_wb_error_o;
 input slave1_wb_stall_o;
 output slave1_wb_stb_i;
 output slave1_wb_we_i;
 input slave2_wb_ack_o;
 output slave2_wb_cyc_i;
 input slave2_wb_error_o;
 input slave2_wb_stall_o;
 output slave2_wb_stb_i;
 output slave2_wb_we_i;
 input slave3_wb_ack_o;
 output slave3_wb_cyc_i;
 input slave3_wb_error_o;
 input slave3_wb_stall_o;
 output slave3_wb_stb_i;
 output slave3_wb_we_i;
 input slave4_wb_ack_o;
 output slave4_wb_cyc_i;
 input slave4_wb_error_o;
 input slave4_wb_stall_o;
 output slave4_wb_stb_i;
 output slave4_wb_we_i;
 input wb_clk_i;
 input wb_rst_i;
 input [27:0] master0_wb_adr_o;
 output [31:0] master0_wb_data_i;
 input [31:0] master0_wb_data_o;
 input [3:0] master0_wb_sel_o;
 input [27:0] master1_wb_adr_o;
 output [31:0] master1_wb_data_i;
 input [31:0] master1_wb_data_o;
 input [3:0] master1_wb_sel_o;
 input [27:0] master2_wb_adr_o;
 output [31:0] master2_wb_data_i;
 input [31:0] master2_wb_data_o;
 input [3:0] master2_wb_sel_o;
 output [1:0] probe_master0_currentSlave;
 output [1:0] probe_master1_currentSlave;
 output [1:0] probe_master2_currentSlave;
 output [1:0] probe_master3_currentSlave;
 output [1:0] probe_slave0_currentMaster;
 output [1:0] probe_slave1_currentMaster;
 output [1:0] probe_slave2_currentMaster;
 output [1:0] probe_slave3_currentMaster;
 output [23:0] slave0_wb_adr_i;
 output [31:0] slave0_wb_data_i;
 input [31:0] slave0_wb_data_o;
 output [3:0] slave0_wb_sel_i;
 output [23:0] slave1_wb_adr_i;
 output [31:0] slave1_wb_data_i;
 input [31:0] slave1_wb_data_o;
 output [3:0] slave1_wb_sel_i;
 output [23:0] slave2_wb_adr_i;
 output [31:0] slave2_wb_data_i;
 input [31:0] slave2_wb_data_o;
 output [3:0] slave2_wb_sel_i;
 output [23:0] slave3_wb_adr_i;
 output [31:0] slave3_wb_data_i;
 input [31:0] slave3_wb_data_o;
 output [3:0] slave3_wb_sel_i;
 output [23:0] slave4_wb_adr_i;
 output [31:0] slave4_wb_data_i;
 input [31:0] slave4_wb_data_o;
 output [3:0] slave4_wb_sel_i;

 wire net1017;
 wire net1018;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \slave0MultiMaster.arbiter.currentMaster[0] ;
 wire \slave0MultiMaster.arbiter.currentMaster[1] ;
 wire \slave1MultiMaster.arbiter.currentMaster[0] ;
 wire \slave1MultiMaster.arbiter.currentMaster[1] ;
 wire \slave2MultiMaster.arbiter.currentMaster[0] ;
 wire \slave2MultiMaster.arbiter.currentMaster[1] ;
 wire \slave3MultiMaster.arbiter.currentMaster[0] ;
 wire \slave3MultiMaster.arbiter.currentMaster[1] ;
 wire \slave4MultiMaster.arbiter.currentMaster[0] ;
 wire \slave4MultiMaster.arbiter.currentMaster[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_475 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_476 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_477 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_478 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_479 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_480 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_481 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_482 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_483 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_484 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_485 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_486 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_487 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_488 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_489 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_490 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_491 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_492 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_493 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_494 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_495 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_496 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_497 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_498 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_499 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_500 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_501 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_502 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_503 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_504 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_505 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_506 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_507 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_508 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_509 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_510 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_511 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_512 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_513 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_514 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_515 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_516 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_517 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_518 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_519 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_520 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_521 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_522 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_523 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_524 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_525 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_526 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_527 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_528 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_529 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_530 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_531 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_532 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_533 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_534 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_535 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_536 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_537 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_538 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_539 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_540 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_541 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_542 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_543 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_544 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_545 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_546 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_547 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_548 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_549 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_550 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_551 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_552 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_553 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_554 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_555 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_556 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_557 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_558 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_559 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_560 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_561 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_562 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_563 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_564 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_565 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_566 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_567 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_568 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_569 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_570 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_571 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_572 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_573 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_574 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_575 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_576 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_577 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_578 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_579 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_580 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_581 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_582 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_583 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_584 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_585 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_586 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_587 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_588 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_589 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_590 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_591 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_592 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_593 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_594 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_595 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_596 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_597 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_598 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_599 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_600 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_601 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_602 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_603 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_604 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_605 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_606 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_607 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_608 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_609 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_610 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_611 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_612 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_613 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_614 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_615 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_616 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_617 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_618 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_619 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_620 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_621 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_622 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_623 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_624 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_625 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_626 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_627 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_628 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_629 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_630 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_631 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_632 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_633 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_634 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_635 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_636 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_637 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_638 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_639 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_640 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_641 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_642 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_643 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_644 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_645 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_646 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_647 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_648 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_649 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_650 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_651 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_652 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_653 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_654 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_655 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_656 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net53));
 sky130_fd_sc_hd__decap_4 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_290_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_292_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_293_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_293_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_296_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_296_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_296_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_296_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_296_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_296_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_296_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_296_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_296_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_296_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_296_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_296_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_297_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_298_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_298_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_298_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_298_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_298_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_298_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_298_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_298_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_298_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_298_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_298_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_298_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_298_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_298_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_298_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_299_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_299_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_299_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_302_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_303_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_303_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_304_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_304_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_304_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_306_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_306_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_306_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_306_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_306_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_307_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_307_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_308_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_308_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_310_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_314_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_314_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_314_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_314_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_314_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_314_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_314_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_314_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_314_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_316_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_316_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_316_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_316_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_318_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_320_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_320_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_320_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_320_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_322_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_322_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_324_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_324_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_326_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_326_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_326_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_326_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_326_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_326_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_326_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_326_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_328_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_328_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_328_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_328_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_328_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_328_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_330_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_332_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_332_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_332_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_333_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_333_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_333_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_334_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_334_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_339_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_339_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_339_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_343_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_343_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_344_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_344_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_344_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_344_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_345_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_346_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_346_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_346_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_348_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_348_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_348_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_349_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_350_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_350_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_350_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_352_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_352_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_352_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_354_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_354_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_354_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_354_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_354_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_354_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_355_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_355_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_356_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_356_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_356_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_356_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_356_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_356_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_356_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_357_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_357_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_357_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_357_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_357_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_357_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_359_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_359_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_360_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_360_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_360_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_360_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_360_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_361_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_361_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_361_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_361_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_362_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_362_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_363_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_364_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_364_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_364_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_364_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_366_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_366_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_366_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_366_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_366_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_367_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_368_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_368_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_368_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_369_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_369_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_369_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_369_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_370_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_370_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_370_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_370_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_371_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_371_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_371_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_372_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_372_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_372_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_372_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_372_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_373_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_373_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_376_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_376_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_376_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_379_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_380_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_380_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_380_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_380_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_381_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_381_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_381_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_382_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_382_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_384_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_384_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_385_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_385_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_385_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_385_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_385_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_386_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_386_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_387_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_387_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_387_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_387_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_387_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_387_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_388_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_388_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_389_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_389_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_389_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_391_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_391_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_391_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_391_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_392_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_392_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__conb_1 WishboneInterconnect_1017 (.LO(net1017));
 sky130_fd_sc_hd__conb_1 WishboneInterconnect_1018 (.LO(net1018));
 sky130_fd_sc_hd__clkinv_8 _0728_ (.A(net1006),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_6 _0729_ (.A(net1009),
    .Y(_0589_));
 sky130_fd_sc_hd__inv_6 _0730_ (.A(net29),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_2 _0731_ (.A(\slave1MultiMaster.arbiter.currentMaster[1] ),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(\slave2MultiMaster.arbiter.currentMaster[0] ),
    .Y(_0592_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(\slave0MultiMaster.arbiter.currentMaster[1] ),
    .Y(_0593_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(\slave4MultiMaster.arbiter.currentMaster[1] ),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(net340),
    .Y(_0595_));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(net341),
    .Y(_0596_));
 sky130_fd_sc_hd__nor4b_4 _0737_ (.A(net1007),
    .B(net87),
    .C(net86),
    .D_N(net1008),
    .Y(_0597_));
 sky130_fd_sc_hd__or4b_4 _0738_ (.A(net1007),
    .B(net87),
    .C(net86),
    .D_N(net1008),
    .X(_0598_));
 sky130_fd_sc_hd__or4b_1 _0739_ (.A(_0588_),
    .B(\slave1MultiMaster.arbiter.currentMaster[1] ),
    .C(net1000),
    .D_N(\slave1MultiMaster.arbiter.currentMaster[0] ),
    .X(_0599_));
 sky130_fd_sc_hd__or3_4 _0740_ (.A(net152),
    .B(net1010),
    .C(net1012),
    .X(_0600_));
 sky130_fd_sc_hd__clkinv_4 _0741_ (.A(net999),
    .Y(_0601_));
 sky130_fd_sc_hd__nor4b_4 _0742_ (.A(net152),
    .B(net1010),
    .C(net1012),
    .D_N(net1014),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_8 _0743_ (.A(net1014),
    .B(_0601_),
    .Y(_0603_));
 sky130_fd_sc_hd__and4b_2 _0744_ (.A_N(\slave1MultiMaster.arbiter.currentMaster[0] ),
    .B(\slave1MultiMaster.arbiter.currentMaster[1] ),
    .C(net997),
    .D(net1009),
    .X(_0604_));
 sky130_fd_sc_hd__nor4b_4 _0745_ (.A(net18),
    .B(net20),
    .C(net19),
    .D_N(net17),
    .Y(_0605_));
 sky130_fd_sc_hd__or4b_4 _0746_ (.A(net18),
    .B(net20),
    .C(net19),
    .D_N(net17),
    .X(_0606_));
 sky130_fd_sc_hd__nor2_4 _0747_ (.A(net1005),
    .B(net993),
    .Y(_0607_));
 sky130_fd_sc_hd__a21oi_1 _0748_ (.A1(net1006),
    .A2(_0597_),
    .B1(\slave1MultiMaster.arbiter.currentMaster[0] ),
    .Y(_0608_));
 sky130_fd_sc_hd__o211a_1 _0749_ (.A1(_0588_),
    .A2(net1000),
    .B1(net997),
    .C1(net1009),
    .X(_0609_));
 sky130_fd_sc_hd__o41a_4 _0750_ (.A1(_0604_),
    .A2(_0607_),
    .A3(_0608_),
    .A4(_0609_),
    .B1(_0599_),
    .X(_0610_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(net934),
    .Y(net491));
 sky130_fd_sc_hd__o221a_1 _0752_ (.A1(_0588_),
    .A2(net1000),
    .B1(net993),
    .B2(net1005),
    .C1(\slave1MultiMaster.arbiter.currentMaster[1] ),
    .X(_0611_));
 sky130_fd_sc_hd__a211o_1 _0753_ (.A1(\slave1MultiMaster.arbiter.currentMaster[0] ),
    .A2(_0591_),
    .B1(net993),
    .C1(net1005),
    .X(_0612_));
 sky130_fd_sc_hd__a211o_4 _0754_ (.A1(_0609_),
    .A2(_0612_),
    .B1(_0611_),
    .C1(_0604_),
    .X(net492));
 sky130_fd_sc_hd__or3b_4 _0755_ (.A(net1010),
    .B(net1012),
    .C_N(net152),
    .X(_0613_));
 sky130_fd_sc_hd__nor4b_4 _0756_ (.A(net1014),
    .B(net1010),
    .C(net1012),
    .D_N(net152),
    .Y(_0614_));
 sky130_fd_sc_hd__or2_4 _0757_ (.A(net1014),
    .B(net990),
    .X(_0615_));
 sky130_fd_sc_hd__and4_2 _0758_ (.A(net1009),
    .B(\slave2MultiMaster.arbiter.currentMaster[1] ),
    .C(_0592_),
    .D(net985),
    .X(_0616_));
 sky130_fd_sc_hd__a21o_1 _0759_ (.A1(net1009),
    .A2(net985),
    .B1(\slave2MultiMaster.arbiter.currentMaster[1] ),
    .X(_0617_));
 sky130_fd_sc_hd__nor4b_4 _0760_ (.A(net1008),
    .B(net87),
    .C(net86),
    .D_N(net1007),
    .Y(_0618_));
 sky130_fd_sc_hd__or4b_4 _0761_ (.A(net1008),
    .B(net87),
    .C(net86),
    .D_N(net1007),
    .X(_0619_));
 sky130_fd_sc_hd__nand2_8 _0762_ (.A(net1006),
    .B(_0618_),
    .Y(_0620_));
 sky130_fd_sc_hd__and2b_1 _0763_ (.A_N(\slave2MultiMaster.arbiter.currentMaster[1] ),
    .B(\slave2MultiMaster.arbiter.currentMaster[0] ),
    .X(_0621_));
 sky130_fd_sc_hd__nor4b_4 _0764_ (.A(net17),
    .B(net20),
    .C(net19),
    .D_N(net18),
    .Y(_0622_));
 sky130_fd_sc_hd__or4b_4 _0765_ (.A(net17),
    .B(net20),
    .C(net19),
    .D_N(net18),
    .X(_0623_));
 sky130_fd_sc_hd__and3b_1 _0766_ (.A_N(_0621_),
    .B(_0622_),
    .C(net29),
    .X(_0624_));
 sky130_fd_sc_hd__or3_1 _0767_ (.A(net1005),
    .B(_0621_),
    .C(net977),
    .X(_0625_));
 sky130_fd_sc_hd__a31o_4 _0768_ (.A1(_0617_),
    .A2(_0620_),
    .A3(_0625_),
    .B1(_0616_),
    .X(net494));
 sky130_fd_sc_hd__a221o_1 _0769_ (.A1(net1009),
    .A2(net985),
    .B1(_0622_),
    .B2(net29),
    .C1(_0592_),
    .X(_0626_));
 sky130_fd_sc_hd__o31a_4 _0770_ (.A1(_0616_),
    .A2(_0620_),
    .A3(_0624_),
    .B1(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(_0627_),
    .Y(net493));
 sky130_fd_sc_hd__and2b_2 _0772_ (.A_N(\slave3MultiMaster.arbiter.currentMaster[1] ),
    .B(\slave3MultiMaster.arbiter.currentMaster[0] ),
    .X(_0628_));
 sky130_fd_sc_hd__or4bb_4 _0773_ (.A(net20),
    .B(net19),
    .C_N(net18),
    .D_N(net17),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _0774_ (.A(_0590_),
    .B(net973),
    .Y(_0630_));
 sky130_fd_sc_hd__and4bb_2 _0775_ (.A_N(net1010),
    .B_N(net1012),
    .C(net152),
    .D(net1014),
    .X(_0631_));
 sky130_fd_sc_hd__or4bb_4 _0776_ (.A(net1010),
    .B(net1012),
    .C_N(net152),
    .D_N(net1014),
    .X(_0632_));
 sky130_fd_sc_hd__a21o_1 _0777_ (.A1(net1009),
    .A2(net969),
    .B1(\slave3MultiMaster.arbiter.currentMaster[1] ),
    .X(_0633_));
 sky130_fd_sc_hd__and4bb_4 _0778_ (.A_N(net87),
    .B_N(net86),
    .C(net1007),
    .D(net1008),
    .X(_0634_));
 sky130_fd_sc_hd__or4bb_4 _0779_ (.A(net87),
    .B(net86),
    .C_N(net1007),
    .D_N(net1008),
    .X(_0635_));
 sky130_fd_sc_hd__o32a_1 _0780_ (.A1(net1005),
    .A2(_0628_),
    .A3(net974),
    .B1(net965),
    .B2(_0588_),
    .X(_0636_));
 sky130_fd_sc_hd__or4b_4 _0781_ (.A(_0589_),
    .B(\slave3MultiMaster.arbiter.currentMaster[0] ),
    .C(_0632_),
    .D_N(\slave3MultiMaster.arbiter.currentMaster[1] ),
    .X(_0637_));
 sky130_fd_sc_hd__a21bo_4 _0782_ (.A1(_0633_),
    .A2(_0636_),
    .B1_N(_0637_),
    .X(net496));
 sky130_fd_sc_hd__o221a_2 _0783_ (.A1(net1005),
    .A2(net974),
    .B1(_0632_),
    .B2(_0589_),
    .C1(\slave3MultiMaster.arbiter.currentMaster[0] ),
    .X(_0638_));
 sky130_fd_sc_hd__o311a_2 _0784_ (.A1(net1005),
    .A2(_0628_),
    .A3(net974),
    .B1(_0634_),
    .C1(net1006),
    .X(_0639_));
 sky130_fd_sc_hd__a21oi_4 _0785_ (.A1(_0637_),
    .A2(_0639_),
    .B1(_0638_),
    .Y(_0640_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(_0640_),
    .Y(net495));
 sky130_fd_sc_hd__nor4_4 _0787_ (.A(net1007),
    .B(net1008),
    .C(net87),
    .D(net86),
    .Y(_0641_));
 sky130_fd_sc_hd__or4_4 _0788_ (.A(net1007),
    .B(net1008),
    .C(net87),
    .D(net86),
    .X(_0642_));
 sky130_fd_sc_hd__or4b_1 _0789_ (.A(_0588_),
    .B(\slave0MultiMaster.arbiter.currentMaster[1] ),
    .C(net961),
    .D_N(\slave0MultiMaster.arbiter.currentMaster[0] ),
    .X(_0643_));
 sky130_fd_sc_hd__nor4_4 _0790_ (.A(net152),
    .B(net1014),
    .C(net1010),
    .D(net1012),
    .Y(_0644_));
 sky130_fd_sc_hd__or2_4 _0791_ (.A(net1014),
    .B(net999),
    .X(_0645_));
 sky130_fd_sc_hd__o211a_1 _0792_ (.A1(_0588_),
    .A2(net961),
    .B1(net957),
    .C1(net1009),
    .X(_0646_));
 sky130_fd_sc_hd__a21oi_1 _0793_ (.A1(net1006),
    .A2(_0641_),
    .B1(\slave0MultiMaster.arbiter.currentMaster[0] ),
    .Y(_0647_));
 sky130_fd_sc_hd__and4b_2 _0794_ (.A_N(\slave0MultiMaster.arbiter.currentMaster[0] ),
    .B(\slave0MultiMaster.arbiter.currentMaster[1] ),
    .C(net957),
    .D(net1009),
    .X(_0648_));
 sky130_fd_sc_hd__nor4_4 _0795_ (.A(net18),
    .B(net17),
    .C(net20),
    .D(net19),
    .Y(_0649_));
 sky130_fd_sc_hd__or4_4 _0796_ (.A(net18),
    .B(net17),
    .C(net20),
    .D(net19),
    .X(_0650_));
 sky130_fd_sc_hd__nor2_2 _0797_ (.A(_0590_),
    .B(net953),
    .Y(_0651_));
 sky130_fd_sc_hd__o41a_4 _0798_ (.A1(_0646_),
    .A2(_0647_),
    .A3(_0648_),
    .A4(_0651_),
    .B1(_0643_),
    .X(_0652_));
 sky130_fd_sc_hd__inv_2 _0799_ (.A(_0652_),
    .Y(net489));
 sky130_fd_sc_hd__o221a_1 _0800_ (.A1(_0588_),
    .A2(net961),
    .B1(net953),
    .B2(net1005),
    .C1(\slave0MultiMaster.arbiter.currentMaster[1] ),
    .X(_0653_));
 sky130_fd_sc_hd__a211o_1 _0801_ (.A1(\slave0MultiMaster.arbiter.currentMaster[0] ),
    .A2(_0593_),
    .B1(net953),
    .C1(net1005),
    .X(_0654_));
 sky130_fd_sc_hd__a211o_4 _0802_ (.A1(_0646_),
    .A2(_0654_),
    .B1(_0653_),
    .C1(_0648_),
    .X(net490));
 sky130_fd_sc_hd__nor4b_4 _0803_ (.A(net1007),
    .B(net1008),
    .C(net87),
    .D_N(net86),
    .Y(_0655_));
 sky130_fd_sc_hd__or4b_4 _0804_ (.A(net85),
    .B(net84),
    .C(net87),
    .D_N(net86),
    .X(_0656_));
 sky130_fd_sc_hd__or2_1 _0805_ (.A(net343),
    .B(net950),
    .X(_0657_));
 sky130_fd_sc_hd__o221a_1 _0806_ (.A1(net273),
    .A2(net982),
    .B1(net965),
    .B2(net308),
    .C1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__or2_1 _0807_ (.A(net238),
    .B(net1001),
    .X(_0659_));
 sky130_fd_sc_hd__o211a_1 _0808_ (.A1(net203),
    .A2(net962),
    .B1(_0658_),
    .C1(_0659_),
    .X(net414));
 sky130_fd_sc_hd__o22a_1 _0809_ (.A1(net284),
    .A2(net982),
    .B1(net951),
    .B2(net354),
    .X(_0660_));
 sky130_fd_sc_hd__o221a_2 _0810_ (.A1(net249),
    .A2(net1000),
    .B1(net966),
    .B2(net319),
    .C1(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_2 _0811_ (.A0(net214),
    .A1(_0661_),
    .S(net962),
    .X(net425));
 sky130_fd_sc_hd__or2_1 _0812_ (.A(net365),
    .B(net950),
    .X(_0662_));
 sky130_fd_sc_hd__o221a_1 _0813_ (.A1(net295),
    .A2(net982),
    .B1(net968),
    .B2(net330),
    .C1(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__or2_1 _0814_ (.A(net260),
    .B(net1001),
    .X(_0664_));
 sky130_fd_sc_hd__o211a_1 _0815_ (.A1(net225),
    .A2(net962),
    .B1(_0663_),
    .C1(_0664_),
    .X(net436));
 sky130_fd_sc_hd__o22a_1 _0816_ (.A1(net298),
    .A2(net981),
    .B1(net948),
    .B2(net368),
    .X(_0665_));
 sky130_fd_sc_hd__o221a_2 _0817_ (.A1(net263),
    .A2(net1000),
    .B1(net965),
    .B2(net333),
    .C1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_2 _0818_ (.A0(net228),
    .A1(_0666_),
    .S(net962),
    .X(net439));
 sky130_fd_sc_hd__or2_1 _0819_ (.A(net369),
    .B(net950),
    .X(_0667_));
 sky130_fd_sc_hd__o221a_1 _0820_ (.A1(net299),
    .A2(net984),
    .B1(net968),
    .B2(net334),
    .C1(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__or2_1 _0821_ (.A(net264),
    .B(net1001),
    .X(_0669_));
 sky130_fd_sc_hd__o211a_2 _0822_ (.A1(net229),
    .A2(net962),
    .B1(_0668_),
    .C1(_0669_),
    .X(net440));
 sky130_fd_sc_hd__or2_1 _0823_ (.A(net370),
    .B(net949),
    .X(_0670_));
 sky130_fd_sc_hd__o221a_1 _0824_ (.A1(net300),
    .A2(net983),
    .B1(net967),
    .B2(net335),
    .C1(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__or2_1 _0825_ (.A(net265),
    .B(net1002),
    .X(_0672_));
 sky130_fd_sc_hd__o211a_4 _0826_ (.A1(net230),
    .A2(net963),
    .B1(_0671_),
    .C1(_0672_),
    .X(net441));
 sky130_fd_sc_hd__or2_1 _0827_ (.A(net371),
    .B(net951),
    .X(_0673_));
 sky130_fd_sc_hd__o221a_1 _0828_ (.A1(net301),
    .A2(net983),
    .B1(net967),
    .B2(net336),
    .C1(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__or2_1 _0829_ (.A(net266),
    .B(net1003),
    .X(_0675_));
 sky130_fd_sc_hd__o211a_4 _0830_ (.A1(net231),
    .A2(net963),
    .B1(_0674_),
    .C1(_0675_),
    .X(net442));
 sky130_fd_sc_hd__or2_1 _0831_ (.A(net372),
    .B(net949),
    .X(_0676_));
 sky130_fd_sc_hd__o221a_1 _0832_ (.A1(net302),
    .A2(net983),
    .B1(net967),
    .B2(net337),
    .C1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__or2_1 _0833_ (.A(net267),
    .B(net1002),
    .X(_0678_));
 sky130_fd_sc_hd__o211a_4 _0834_ (.A1(net232),
    .A2(net964),
    .B1(_0677_),
    .C1(_0678_),
    .X(net443));
 sky130_fd_sc_hd__o22a_1 _0835_ (.A1(net303),
    .A2(net981),
    .B1(net948),
    .B2(net373),
    .X(_0679_));
 sky130_fd_sc_hd__o221a_1 _0836_ (.A1(net268),
    .A2(net1000),
    .B1(net965),
    .B2(net338),
    .C1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_8 _0837_ (.A0(net233),
    .A1(_0680_),
    .S(_0642_),
    .X(net444));
 sky130_fd_sc_hd__o22a_1 _0838_ (.A1(net304),
    .A2(net982),
    .B1(net950),
    .B2(net374),
    .X(_0681_));
 sky130_fd_sc_hd__o221a_1 _0839_ (.A1(net269),
    .A2(net1001),
    .B1(net968),
    .B2(net339),
    .C1(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_2 _0840_ (.A0(net234),
    .A1(_0682_),
    .S(net964),
    .X(net445));
 sky130_fd_sc_hd__or2_1 _0841_ (.A(net344),
    .B(net950),
    .X(_0683_));
 sky130_fd_sc_hd__o221a_1 _0842_ (.A1(net274),
    .A2(net984),
    .B1(net968),
    .B2(net309),
    .C1(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__or2_1 _0843_ (.A(net239),
    .B(net1001),
    .X(_0685_));
 sky130_fd_sc_hd__o211a_2 _0844_ (.A1(net204),
    .A2(net962),
    .B1(_0684_),
    .C1(_0685_),
    .X(net415));
 sky130_fd_sc_hd__o22a_1 _0845_ (.A1(net275),
    .A2(net984),
    .B1(net968),
    .B2(net310),
    .X(_0686_));
 sky130_fd_sc_hd__o221a_1 _0846_ (.A1(net240),
    .A2(net1001),
    .B1(net950),
    .B2(net345),
    .C1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__o21a_2 _0847_ (.A1(net205),
    .A2(net964),
    .B1(_0687_),
    .X(net416));
 sky130_fd_sc_hd__or2_1 _0848_ (.A(net346),
    .B(net948),
    .X(_0688_));
 sky130_fd_sc_hd__o221a_1 _0849_ (.A1(net276),
    .A2(net981),
    .B1(net965),
    .B2(net311),
    .C1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__or2_1 _0850_ (.A(net241),
    .B(net1000),
    .X(_0690_));
 sky130_fd_sc_hd__o211a_4 _0851_ (.A1(net206),
    .A2(net961),
    .B1(_0689_),
    .C1(_0690_),
    .X(net417));
 sky130_fd_sc_hd__or2_1 _0852_ (.A(net347),
    .B(net949),
    .X(_0691_));
 sky130_fd_sc_hd__o221a_1 _0853_ (.A1(net277),
    .A2(net984),
    .B1(net967),
    .B2(net312),
    .C1(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__or2_1 _0854_ (.A(net242),
    .B(net1002),
    .X(_0693_));
 sky130_fd_sc_hd__o211a_4 _0855_ (.A1(net207),
    .A2(net963),
    .B1(_0692_),
    .C1(_0693_),
    .X(net418));
 sky130_fd_sc_hd__or2_1 _0856_ (.A(net348),
    .B(net949),
    .X(_0694_));
 sky130_fd_sc_hd__o221a_1 _0857_ (.A1(net278),
    .A2(net983),
    .B1(net967),
    .B2(net313),
    .C1(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__or2_1 _0858_ (.A(net243),
    .B(net1002),
    .X(_0696_));
 sky130_fd_sc_hd__o211a_4 _0859_ (.A1(net208),
    .A2(net964),
    .B1(_0695_),
    .C1(_0696_),
    .X(net419));
 sky130_fd_sc_hd__or2_1 _0860_ (.A(net349),
    .B(net948),
    .X(_0697_));
 sky130_fd_sc_hd__o221a_1 _0861_ (.A1(net279),
    .A2(net981),
    .B1(net965),
    .B2(net314),
    .C1(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__or2_1 _0862_ (.A(net244),
    .B(net1000),
    .X(_0699_));
 sky130_fd_sc_hd__o211a_4 _0863_ (.A1(net209),
    .A2(net961),
    .B1(_0698_),
    .C1(_0699_),
    .X(net420));
 sky130_fd_sc_hd__or2_1 _0864_ (.A(net350),
    .B(net948),
    .X(_0700_));
 sky130_fd_sc_hd__o221a_1 _0865_ (.A1(net280),
    .A2(net981),
    .B1(net966),
    .B2(net315),
    .C1(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__or2_1 _0866_ (.A(net245),
    .B(net1004),
    .X(_0702_));
 sky130_fd_sc_hd__o211a_4 _0867_ (.A1(net210),
    .A2(net961),
    .B1(_0701_),
    .C1(_0702_),
    .X(net421));
 sky130_fd_sc_hd__o22a_1 _0868_ (.A1(net281),
    .A2(net981),
    .B1(net951),
    .B2(net351),
    .X(_0703_));
 sky130_fd_sc_hd__o221a_4 _0869_ (.A1(net246),
    .A2(net1004),
    .B1(net965),
    .B2(net316),
    .C1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_8 _0870_ (.A0(net211),
    .A1(_0704_),
    .S(net961),
    .X(net422));
 sky130_fd_sc_hd__or2_1 _0871_ (.A(net352),
    .B(net948),
    .X(_0705_));
 sky130_fd_sc_hd__o221a_1 _0872_ (.A1(net282),
    .A2(net981),
    .B1(net966),
    .B2(net317),
    .C1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__or2_1 _0873_ (.A(net247),
    .B(net1004),
    .X(_0707_));
 sky130_fd_sc_hd__o211a_4 _0874_ (.A1(net212),
    .A2(net961),
    .B1(_0706_),
    .C1(_0707_),
    .X(net423));
 sky130_fd_sc_hd__or2_1 _0875_ (.A(net353),
    .B(net949),
    .X(_0708_));
 sky130_fd_sc_hd__o221a_1 _0876_ (.A1(net283),
    .A2(net983),
    .B1(net967),
    .B2(net318),
    .C1(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__or2_1 _0877_ (.A(net248),
    .B(net1002),
    .X(_0710_));
 sky130_fd_sc_hd__o211a_4 _0878_ (.A1(net213),
    .A2(net963),
    .B1(_0709_),
    .C1(_0710_),
    .X(net424));
 sky130_fd_sc_hd__or2_1 _0879_ (.A(net355),
    .B(net950),
    .X(_0711_));
 sky130_fd_sc_hd__o221a_1 _0880_ (.A1(net285),
    .A2(net981),
    .B1(net968),
    .B2(net320),
    .C1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__or2_1 _0881_ (.A(net250),
    .B(net1001),
    .X(_0713_));
 sky130_fd_sc_hd__o211a_4 _0882_ (.A1(net215),
    .A2(net962),
    .B1(_0712_),
    .C1(_0713_),
    .X(net426));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(net356),
    .B(net948),
    .X(_0714_));
 sky130_fd_sc_hd__o221a_1 _0884_ (.A1(net286),
    .A2(net982),
    .B1(net966),
    .B2(net321),
    .C1(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__or2_1 _0885_ (.A(net251),
    .B(net1000),
    .X(_0716_));
 sky130_fd_sc_hd__o211a_4 _0886_ (.A1(net216),
    .A2(net961),
    .B1(_0715_),
    .C1(_0716_),
    .X(net427));
 sky130_fd_sc_hd__or2_1 _0887_ (.A(net357),
    .B(net950),
    .X(_0717_));
 sky130_fd_sc_hd__o221a_1 _0888_ (.A1(net287),
    .A2(net981),
    .B1(net968),
    .B2(net322),
    .C1(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__or2_1 _0889_ (.A(net252),
    .B(net1003),
    .X(_0719_));
 sky130_fd_sc_hd__o211a_4 _0890_ (.A1(net217),
    .A2(net962),
    .B1(_0718_),
    .C1(_0719_),
    .X(net428));
 sky130_fd_sc_hd__or2_1 _0891_ (.A(net358),
    .B(net951),
    .X(_0720_));
 sky130_fd_sc_hd__o221a_2 _0892_ (.A1(net288),
    .A2(net984),
    .B1(net968),
    .B2(net323),
    .C1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(net253),
    .B(net1003),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_2 _0894_ (.A1(net218),
    .A2(net963),
    .B1(_0721_),
    .C1(_0722_),
    .X(net429));
 sky130_fd_sc_hd__o22a_1 _0895_ (.A1(net289),
    .A2(net982),
    .B1(net948),
    .B2(net359),
    .X(_0723_));
 sky130_fd_sc_hd__o221a_4 _0896_ (.A1(net254),
    .A2(net1001),
    .B1(net966),
    .B2(net324),
    .C1(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_8 _0897_ (.A0(net219),
    .A1(_0724_),
    .S(net962),
    .X(net430));
 sky130_fd_sc_hd__or2_1 _0898_ (.A(net360),
    .B(net949),
    .X(_0725_));
 sky130_fd_sc_hd__o221a_1 _0899_ (.A1(net290),
    .A2(net983),
    .B1(net967),
    .B2(net325),
    .C1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__or2_1 _0900_ (.A(net255),
    .B(net1002),
    .X(_0727_));
 sky130_fd_sc_hd__o211a_4 _0901_ (.A1(net220),
    .A2(net964),
    .B1(_0726_),
    .C1(_0727_),
    .X(net431));
 sky130_fd_sc_hd__or2_1 _0902_ (.A(net361),
    .B(net949),
    .X(_0010_));
 sky130_fd_sc_hd__o221a_1 _0903_ (.A1(net291),
    .A2(net983),
    .B1(net967),
    .B2(net326),
    .C1(_0010_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _0904_ (.A(net256),
    .B(net1002),
    .X(_0012_));
 sky130_fd_sc_hd__o211a_4 _0905_ (.A1(net221),
    .A2(net963),
    .B1(_0011_),
    .C1(_0012_),
    .X(net432));
 sky130_fd_sc_hd__or2_1 _0906_ (.A(net362),
    .B(net949),
    .X(_0013_));
 sky130_fd_sc_hd__o221a_1 _0907_ (.A1(net292),
    .A2(net983),
    .B1(net967),
    .B2(net327),
    .C1(_0013_),
    .X(_0014_));
 sky130_fd_sc_hd__or2_1 _0908_ (.A(net257),
    .B(net1002),
    .X(_0015_));
 sky130_fd_sc_hd__o211a_2 _0909_ (.A1(net222),
    .A2(net963),
    .B1(_0014_),
    .C1(_0015_),
    .X(net433));
 sky130_fd_sc_hd__o22a_1 _0910_ (.A1(net293),
    .A2(net982),
    .B1(net948),
    .B2(net363),
    .X(_0016_));
 sky130_fd_sc_hd__o221a_4 _0911_ (.A1(net258),
    .A2(net1001),
    .B1(net965),
    .B2(net328),
    .C1(_0016_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_2 _0912_ (.A0(net223),
    .A1(_0017_),
    .S(net963),
    .X(net434));
 sky130_fd_sc_hd__o22a_1 _0913_ (.A1(net294),
    .A2(net982),
    .B1(net966),
    .B2(net329),
    .X(_0018_));
 sky130_fd_sc_hd__o221a_4 _0914_ (.A1(net259),
    .A2(net1001),
    .B1(net950),
    .B2(net364),
    .C1(_0018_),
    .X(_0019_));
 sky130_fd_sc_hd__o21a_2 _0915_ (.A1(net224),
    .A2(net963),
    .B1(_0019_),
    .X(net435));
 sky130_fd_sc_hd__or2_1 _0916_ (.A(net366),
    .B(net949),
    .X(_0020_));
 sky130_fd_sc_hd__o221a_1 _0917_ (.A1(net296),
    .A2(net983),
    .B1(net968),
    .B2(net331),
    .C1(_0020_),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _0918_ (.A(net261),
    .B(net1002),
    .X(_0022_));
 sky130_fd_sc_hd__o211a_2 _0919_ (.A1(net226),
    .A2(net964),
    .B1(_0021_),
    .C1(_0022_),
    .X(net437));
 sky130_fd_sc_hd__or2_1 _0920_ (.A(net367),
    .B(net949),
    .X(_0023_));
 sky130_fd_sc_hd__o221a_1 _0921_ (.A1(net297),
    .A2(net983),
    .B1(net967),
    .B2(net332),
    .C1(_0023_),
    .X(_0024_));
 sky130_fd_sc_hd__or2_1 _0922_ (.A(net262),
    .B(net1002),
    .X(_0025_));
 sky130_fd_sc_hd__o211a_2 _0923_ (.A1(net227),
    .A2(net963),
    .B1(_0024_),
    .C1(_0025_),
    .X(net438));
 sky130_fd_sc_hd__nor2_1 _0924_ (.A(_0595_),
    .B(net965),
    .Y(_0026_));
 sky130_fd_sc_hd__a221o_1 _0925_ (.A1(net305),
    .A2(_0618_),
    .B1(_0655_),
    .B2(net375),
    .C1(_0026_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _0926_ (.A(net270),
    .B(_0597_),
    .X(_0028_));
 sky130_fd_sc_hd__a211o_4 _0927_ (.A1(net235),
    .A2(_0641_),
    .B1(_0027_),
    .C1(_0028_),
    .X(net446));
 sky130_fd_sc_hd__a22o_1 _0928_ (.A1(net306),
    .A2(_0618_),
    .B1(_0655_),
    .B2(net376),
    .X(_0029_));
 sky130_fd_sc_hd__a221o_4 _0929_ (.A1(net271),
    .A2(_0597_),
    .B1(_0634_),
    .B2(net341),
    .C1(_0029_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_2 _0930_ (.A0(net236),
    .A1(_0030_),
    .S(net962),
    .X(net447));
 sky130_fd_sc_hd__nor2_1 _0931_ (.A(_0588_),
    .B(_0655_),
    .Y(_0031_));
 sky130_fd_sc_hd__a211o_1 _0932_ (.A1(net342),
    .A2(_0655_),
    .B1(_0031_),
    .C1(_0634_),
    .X(_0032_));
 sky130_fd_sc_hd__o21a_1 _0933_ (.A1(net307),
    .A2(net965),
    .B1(net981),
    .X(_0033_));
 sky130_fd_sc_hd__a221o_1 _0934_ (.A1(net272),
    .A2(_0618_),
    .B1(_0032_),
    .B2(_0033_),
    .C1(_0597_),
    .X(_0034_));
 sky130_fd_sc_hd__o21a_1 _0935_ (.A1(net237),
    .A2(net1000),
    .B1(net961),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_4 _0936_ (.A1(net202),
    .A2(_0641_),
    .B1(_0034_),
    .B2(_0035_),
    .X(net413));
 sky130_fd_sc_hd__nor4b_4 _0937_ (.A(net18),
    .B(net17),
    .C(net20),
    .D_N(net19),
    .Y(_0036_));
 sky130_fd_sc_hd__or4b_4 _0938_ (.A(net18),
    .B(net17),
    .C(net20),
    .D_N(net19),
    .X(_0037_));
 sky130_fd_sc_hd__or2_1 _0939_ (.A(net343),
    .B(net945),
    .X(_0038_));
 sky130_fd_sc_hd__o221a_2 _0940_ (.A1(net273),
    .A2(net979),
    .B1(net975),
    .B2(net308),
    .C1(_0038_),
    .X(_0039_));
 sky130_fd_sc_hd__or2_1 _0941_ (.A(net238),
    .B(net994),
    .X(_0040_));
 sky130_fd_sc_hd__o211a_4 _0942_ (.A1(net203),
    .A2(net952),
    .B1(_0039_),
    .C1(_0040_),
    .X(net379));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(net354),
    .B(net947),
    .X(_0041_));
 sky130_fd_sc_hd__o221a_1 _0944_ (.A1(net284),
    .A2(net977),
    .B1(net973),
    .B2(net319),
    .C1(_0041_),
    .X(_0042_));
 sky130_fd_sc_hd__or2_1 _0945_ (.A(net249),
    .B(net993),
    .X(_0043_));
 sky130_fd_sc_hd__o211a_4 _0946_ (.A1(net214),
    .A2(net953),
    .B1(_0042_),
    .C1(_0043_),
    .X(net390));
 sky130_fd_sc_hd__or2_1 _0947_ (.A(net365),
    .B(net945),
    .X(_0044_));
 sky130_fd_sc_hd__o221a_1 _0948_ (.A1(net295),
    .A2(net979),
    .B1(net975),
    .B2(net330),
    .C1(_0044_),
    .X(_0045_));
 sky130_fd_sc_hd__or2_1 _0949_ (.A(net260),
    .B(net994),
    .X(_0046_));
 sky130_fd_sc_hd__o211a_4 _0950_ (.A1(net225),
    .A2(net954),
    .B1(_0045_),
    .C1(_0046_),
    .X(net401));
 sky130_fd_sc_hd__or2_1 _0951_ (.A(net368),
    .B(net947),
    .X(_0047_));
 sky130_fd_sc_hd__o221a_1 _0952_ (.A1(net298),
    .A2(net977),
    .B1(net973),
    .B2(net333),
    .C1(_0047_),
    .X(_0048_));
 sky130_fd_sc_hd__or2_1 _0953_ (.A(net263),
    .B(net996),
    .X(_0049_));
 sky130_fd_sc_hd__o211a_4 _0954_ (.A1(net228),
    .A2(net952),
    .B1(_0048_),
    .C1(_0049_),
    .X(net404));
 sky130_fd_sc_hd__or2_1 _0955_ (.A(net369),
    .B(net945),
    .X(_0050_));
 sky130_fd_sc_hd__o221a_1 _0956_ (.A1(net299),
    .A2(net979),
    .B1(net975),
    .B2(net334),
    .C1(_0050_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_1 _0957_ (.A(net264),
    .B(net994),
    .X(_0052_));
 sky130_fd_sc_hd__o211a_4 _0958_ (.A1(net229),
    .A2(net954),
    .B1(_0051_),
    .C1(_0052_),
    .X(net405));
 sky130_fd_sc_hd__or2_1 _0959_ (.A(net370),
    .B(net946),
    .X(_0053_));
 sky130_fd_sc_hd__o221a_1 _0960_ (.A1(net300),
    .A2(net978),
    .B1(net976),
    .B2(net335),
    .C1(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__or2_1 _0961_ (.A(net265),
    .B(net995),
    .X(_0055_));
 sky130_fd_sc_hd__o211a_4 _0962_ (.A1(net230),
    .A2(net955),
    .B1(_0054_),
    .C1(_0055_),
    .X(net406));
 sky130_fd_sc_hd__or2_1 _0963_ (.A(net371),
    .B(net946),
    .X(_0056_));
 sky130_fd_sc_hd__o221a_1 _0964_ (.A1(net301),
    .A2(net980),
    .B1(net976),
    .B2(net336),
    .C1(_0056_),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _0965_ (.A(net266),
    .B(net995),
    .X(_0058_));
 sky130_fd_sc_hd__o211a_4 _0966_ (.A1(net231),
    .A2(net955),
    .B1(_0057_),
    .C1(_0058_),
    .X(net407));
 sky130_fd_sc_hd__or2_1 _0967_ (.A(net372),
    .B(net946),
    .X(_0059_));
 sky130_fd_sc_hd__o221a_1 _0968_ (.A1(net302),
    .A2(net980),
    .B1(net976),
    .B2(net337),
    .C1(_0059_),
    .X(_0060_));
 sky130_fd_sc_hd__or2_1 _0969_ (.A(net267),
    .B(net995),
    .X(_0061_));
 sky130_fd_sc_hd__o211a_4 _0970_ (.A1(net232),
    .A2(net954),
    .B1(_0060_),
    .C1(_0061_),
    .X(net408));
 sky130_fd_sc_hd__or2_1 _0971_ (.A(net373),
    .B(net944),
    .X(_0062_));
 sky130_fd_sc_hd__o221a_1 _0972_ (.A1(net303),
    .A2(net977),
    .B1(net973),
    .B2(net338),
    .C1(_0062_),
    .X(_0063_));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(net268),
    .B(net993),
    .X(_0064_));
 sky130_fd_sc_hd__o211a_4 _0974_ (.A1(net233),
    .A2(net952),
    .B1(_0063_),
    .C1(_0064_),
    .X(net409));
 sky130_fd_sc_hd__or2_1 _0975_ (.A(net374),
    .B(net945),
    .X(_0065_));
 sky130_fd_sc_hd__o221a_1 _0976_ (.A1(net304),
    .A2(net979),
    .B1(net975),
    .B2(net339),
    .C1(_0065_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _0977_ (.A(net269),
    .B(net994),
    .X(_0067_));
 sky130_fd_sc_hd__o211a_4 _0978_ (.A1(net234),
    .A2(net954),
    .B1(_0066_),
    .C1(_0067_),
    .X(net410));
 sky130_fd_sc_hd__or2_1 _0979_ (.A(net344),
    .B(net945),
    .X(_0068_));
 sky130_fd_sc_hd__o221a_1 _0980_ (.A1(net274),
    .A2(net979),
    .B1(net975),
    .B2(net309),
    .C1(_0068_),
    .X(_0069_));
 sky130_fd_sc_hd__or2_1 _0981_ (.A(net239),
    .B(net994),
    .X(_0070_));
 sky130_fd_sc_hd__o211a_4 _0982_ (.A1(net204),
    .A2(net954),
    .B1(_0069_),
    .C1(_0070_),
    .X(net380));
 sky130_fd_sc_hd__or2_1 _0983_ (.A(net345),
    .B(net945),
    .X(_0071_));
 sky130_fd_sc_hd__o221a_2 _0984_ (.A1(net275),
    .A2(net979),
    .B1(net975),
    .B2(net310),
    .C1(_0071_),
    .X(_0072_));
 sky130_fd_sc_hd__or2_1 _0985_ (.A(net240),
    .B(net994),
    .X(_0073_));
 sky130_fd_sc_hd__o211a_4 _0986_ (.A1(net205),
    .A2(net952),
    .B1(_0072_),
    .C1(_0073_),
    .X(net381));
 sky130_fd_sc_hd__or2_1 _0987_ (.A(net346),
    .B(net944),
    .X(_0074_));
 sky130_fd_sc_hd__o221a_1 _0988_ (.A1(net276),
    .A2(net977),
    .B1(net973),
    .B2(net311),
    .C1(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__or2_1 _0989_ (.A(net241),
    .B(net996),
    .X(_0076_));
 sky130_fd_sc_hd__o211a_4 _0990_ (.A1(net206),
    .A2(net952),
    .B1(_0075_),
    .C1(_0076_),
    .X(net382));
 sky130_fd_sc_hd__or2_1 _0991_ (.A(net347),
    .B(net947),
    .X(_0077_));
 sky130_fd_sc_hd__o221a_1 _0992_ (.A1(net277),
    .A2(net978),
    .B1(_0629_),
    .B2(net312),
    .C1(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__or2_1 _0993_ (.A(net242),
    .B(net995),
    .X(_0079_));
 sky130_fd_sc_hd__o211a_4 _0994_ (.A1(net207),
    .A2(net955),
    .B1(_0078_),
    .C1(_0079_),
    .X(net383));
 sky130_fd_sc_hd__or2_1 _0995_ (.A(net348),
    .B(net946),
    .X(_0080_));
 sky130_fd_sc_hd__o221a_1 _0996_ (.A1(net278),
    .A2(net978),
    .B1(net976),
    .B2(net313),
    .C1(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__or2_1 _0997_ (.A(net243),
    .B(net995),
    .X(_0082_));
 sky130_fd_sc_hd__o211a_4 _0998_ (.A1(net208),
    .A2(net954),
    .B1(_0081_),
    .C1(_0082_),
    .X(net384));
 sky130_fd_sc_hd__or2_1 _0999_ (.A(net349),
    .B(net944),
    .X(_0083_));
 sky130_fd_sc_hd__o221a_1 _1000_ (.A1(net279),
    .A2(net977),
    .B1(net974),
    .B2(net314),
    .C1(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__or2_1 _1001_ (.A(net244),
    .B(net993),
    .X(_0085_));
 sky130_fd_sc_hd__o211a_4 _1002_ (.A1(net209),
    .A2(net953),
    .B1(_0084_),
    .C1(_0085_),
    .X(net385));
 sky130_fd_sc_hd__or2_1 _1003_ (.A(net350),
    .B(net944),
    .X(_0086_));
 sky130_fd_sc_hd__o221a_1 _1004_ (.A1(net280),
    .A2(net977),
    .B1(net974),
    .B2(net315),
    .C1(_0086_),
    .X(_0087_));
 sky130_fd_sc_hd__or2_1 _1005_ (.A(net245),
    .B(net996),
    .X(_0088_));
 sky130_fd_sc_hd__o211a_4 _1006_ (.A1(net210),
    .A2(net952),
    .B1(_0087_),
    .C1(_0088_),
    .X(net386));
 sky130_fd_sc_hd__or2_1 _1007_ (.A(net351),
    .B(net947),
    .X(_0089_));
 sky130_fd_sc_hd__o221a_1 _1008_ (.A1(net281),
    .A2(net980),
    .B1(net973),
    .B2(net316),
    .C1(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _1009_ (.A(net246),
    .B(net993),
    .X(_0091_));
 sky130_fd_sc_hd__o211a_4 _1010_ (.A1(net211),
    .A2(net953),
    .B1(_0090_),
    .C1(_0091_),
    .X(net387));
 sky130_fd_sc_hd__or2_1 _1011_ (.A(net352),
    .B(net944),
    .X(_0092_));
 sky130_fd_sc_hd__o221a_1 _1012_ (.A1(net282),
    .A2(net977),
    .B1(net973),
    .B2(net317),
    .C1(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__or2_1 _1013_ (.A(net247),
    .B(net996),
    .X(_0094_));
 sky130_fd_sc_hd__o211a_4 _1014_ (.A1(net212),
    .A2(net952),
    .B1(_0093_),
    .C1(_0094_),
    .X(net388));
 sky130_fd_sc_hd__or2_1 _1015_ (.A(net353),
    .B(net946),
    .X(_0095_));
 sky130_fd_sc_hd__o221a_1 _1016_ (.A1(net283),
    .A2(net978),
    .B1(net976),
    .B2(net318),
    .C1(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__or2_1 _1017_ (.A(net248),
    .B(net995),
    .X(_0097_));
 sky130_fd_sc_hd__o211a_4 _1018_ (.A1(net213),
    .A2(net955),
    .B1(_0096_),
    .C1(_0097_),
    .X(net389));
 sky130_fd_sc_hd__or2_1 _1019_ (.A(net355),
    .B(net945),
    .X(_0098_));
 sky130_fd_sc_hd__o221a_1 _1020_ (.A1(net285),
    .A2(net979),
    .B1(net975),
    .B2(net320),
    .C1(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__or2_1 _1021_ (.A(net250),
    .B(net994),
    .X(_0100_));
 sky130_fd_sc_hd__o211a_4 _1022_ (.A1(net215),
    .A2(net954),
    .B1(_0099_),
    .C1(_0100_),
    .X(net391));
 sky130_fd_sc_hd__or2_1 _1023_ (.A(net356),
    .B(net944),
    .X(_0101_));
 sky130_fd_sc_hd__o221a_1 _1024_ (.A1(net286),
    .A2(net977),
    .B1(net973),
    .B2(net321),
    .C1(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__or2_1 _1025_ (.A(net251),
    .B(net993),
    .X(_0103_));
 sky130_fd_sc_hd__o211a_4 _1026_ (.A1(net216),
    .A2(net953),
    .B1(_0102_),
    .C1(_0103_),
    .X(net392));
 sky130_fd_sc_hd__or2_1 _1027_ (.A(net357),
    .B(net945),
    .X(_0104_));
 sky130_fd_sc_hd__o221a_1 _1028_ (.A1(net287),
    .A2(net979),
    .B1(net975),
    .B2(net322),
    .C1(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _1029_ (.A(net252),
    .B(net994),
    .X(_0106_));
 sky130_fd_sc_hd__o211a_4 _1030_ (.A1(net217),
    .A2(net954),
    .B1(_0105_),
    .C1(_0106_),
    .X(net393));
 sky130_fd_sc_hd__or2_1 _1031_ (.A(net358),
    .B(net947),
    .X(_0107_));
 sky130_fd_sc_hd__o221a_1 _1032_ (.A1(net288),
    .A2(net978),
    .B1(_0629_),
    .B2(net323),
    .C1(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__or2_1 _1033_ (.A(net253),
    .B(net995),
    .X(_0109_));
 sky130_fd_sc_hd__o211a_4 _1034_ (.A1(net218),
    .A2(net955),
    .B1(_0108_),
    .C1(_0109_),
    .X(net394));
 sky130_fd_sc_hd__or2_1 _1035_ (.A(net359),
    .B(net944),
    .X(_0110_));
 sky130_fd_sc_hd__o221a_1 _1036_ (.A1(net289),
    .A2(net979),
    .B1(net973),
    .B2(net324),
    .C1(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__or2_1 _1037_ (.A(net254),
    .B(net994),
    .X(_0112_));
 sky130_fd_sc_hd__o211a_4 _1038_ (.A1(net219),
    .A2(net952),
    .B1(_0111_),
    .C1(_0112_),
    .X(net395));
 sky130_fd_sc_hd__or2_1 _1039_ (.A(net360),
    .B(net945),
    .X(_0113_));
 sky130_fd_sc_hd__o221a_1 _1040_ (.A1(net290),
    .A2(net978),
    .B1(net975),
    .B2(net325),
    .C1(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__or2_1 _1041_ (.A(net255),
    .B(net995),
    .X(_0115_));
 sky130_fd_sc_hd__o211a_4 _1042_ (.A1(net220),
    .A2(net954),
    .B1(_0114_),
    .C1(_0115_),
    .X(net396));
 sky130_fd_sc_hd__or2_1 _1043_ (.A(net361),
    .B(net946),
    .X(_0116_));
 sky130_fd_sc_hd__o221a_1 _1044_ (.A1(net291),
    .A2(net978),
    .B1(net976),
    .B2(net326),
    .C1(_0116_),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _1045_ (.A(net256),
    .B(net996),
    .X(_0118_));
 sky130_fd_sc_hd__o211a_4 _1046_ (.A1(net221),
    .A2(net954),
    .B1(_0117_),
    .C1(_0118_),
    .X(net397));
 sky130_fd_sc_hd__or2_1 _1047_ (.A(net362),
    .B(net946),
    .X(_0119_));
 sky130_fd_sc_hd__o221a_1 _1048_ (.A1(net292),
    .A2(net978),
    .B1(net976),
    .B2(net327),
    .C1(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__or2_1 _1049_ (.A(net257),
    .B(net995),
    .X(_0121_));
 sky130_fd_sc_hd__o211a_4 _1050_ (.A1(net222),
    .A2(net955),
    .B1(_0120_),
    .C1(_0121_),
    .X(net398));
 sky130_fd_sc_hd__or2_1 _1051_ (.A(net363),
    .B(net944),
    .X(_0122_));
 sky130_fd_sc_hd__o221a_1 _1052_ (.A1(net293),
    .A2(net980),
    .B1(net973),
    .B2(net328),
    .C1(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _1053_ (.A(net258),
    .B(net993),
    .X(_0124_));
 sky130_fd_sc_hd__o211a_4 _1054_ (.A1(net223),
    .A2(net952),
    .B1(_0123_),
    .C1(_0124_),
    .X(net399));
 sky130_fd_sc_hd__or2_1 _1055_ (.A(net364),
    .B(net945),
    .X(_0125_));
 sky130_fd_sc_hd__o221a_1 _1056_ (.A1(net294),
    .A2(net979),
    .B1(net975),
    .B2(net329),
    .C1(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__or2_1 _1057_ (.A(net259),
    .B(net994),
    .X(_0127_));
 sky130_fd_sc_hd__o211a_4 _1058_ (.A1(net224),
    .A2(net952),
    .B1(_0126_),
    .C1(_0127_),
    .X(net400));
 sky130_fd_sc_hd__or2_1 _1059_ (.A(net366),
    .B(net946),
    .X(_0128_));
 sky130_fd_sc_hd__o221a_1 _1060_ (.A1(net296),
    .A2(net978),
    .B1(net976),
    .B2(net331),
    .C1(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _1061_ (.A(net261),
    .B(net996),
    .X(_0130_));
 sky130_fd_sc_hd__o211a_4 _1062_ (.A1(net226),
    .A2(net955),
    .B1(_0129_),
    .C1(_0130_),
    .X(net402));
 sky130_fd_sc_hd__or2_1 _1063_ (.A(net367),
    .B(net946),
    .X(_0131_));
 sky130_fd_sc_hd__o221a_1 _1064_ (.A1(net297),
    .A2(net978),
    .B1(net976),
    .B2(net332),
    .C1(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _1065_ (.A(net262),
    .B(net995),
    .X(_0133_));
 sky130_fd_sc_hd__o211a_4 _1066_ (.A1(net227),
    .A2(net955),
    .B1(_0132_),
    .C1(_0133_),
    .X(net403));
 sky130_fd_sc_hd__nor2_1 _1067_ (.A(_0595_),
    .B(net974),
    .Y(_0134_));
 sky130_fd_sc_hd__a221o_1 _1068_ (.A1(net305),
    .A2(_0622_),
    .B1(_0036_),
    .B2(net375),
    .C1(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _1069_ (.A(net270),
    .B(_0605_),
    .X(_0136_));
 sky130_fd_sc_hd__a211o_2 _1070_ (.A1(net235),
    .A2(_0649_),
    .B1(_0135_),
    .C1(_0136_),
    .X(net411));
 sky130_fd_sc_hd__nor2_1 _1071_ (.A(_0596_),
    .B(net974),
    .Y(_0137_));
 sky130_fd_sc_hd__a221o_1 _1072_ (.A1(net306),
    .A2(_0622_),
    .B1(_0036_),
    .B2(net376),
    .C1(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__and2_1 _1073_ (.A(net271),
    .B(_0605_),
    .X(_0139_));
 sky130_fd_sc_hd__a211o_2 _1074_ (.A1(net236),
    .A2(_0649_),
    .B1(_0138_),
    .C1(_0139_),
    .X(net412));
 sky130_fd_sc_hd__a21bo_1 _1075_ (.A1(net342),
    .A2(_0036_),
    .B1_N(net974),
    .X(_0140_));
 sky130_fd_sc_hd__a21o_1 _1076_ (.A1(net29),
    .A2(net944),
    .B1(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__o21a_1 _1077_ (.A1(net307),
    .A2(net974),
    .B1(net977),
    .X(_0142_));
 sky130_fd_sc_hd__a221o_1 _1078_ (.A1(net272),
    .A2(_0622_),
    .B1(_0141_),
    .B2(_0142_),
    .C1(_0605_),
    .X(_0143_));
 sky130_fd_sc_hd__o21a_1 _1079_ (.A1(net237),
    .A2(net993),
    .B1(net953),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_2 _1080_ (.A1(net202),
    .A2(_0649_),
    .B1(_0143_),
    .B2(_0144_),
    .X(net378));
 sky130_fd_sc_hd__nor2_1 _1081_ (.A(net919),
    .B(net867),
    .Y(_0145_));
 sky130_fd_sc_hd__mux2_1 _1082_ (.A0(net1),
    .A1(net135),
    .S(net867),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_2 _1083_ (.A1(net68),
    .A2(net845),
    .B1(_0146_),
    .B2(net919),
    .X(net497));
 sky130_fd_sc_hd__mux2_1 _1084_ (.A0(net12),
    .A1(net146),
    .S(net867),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_2 _1085_ (.A1(net79),
    .A2(net848),
    .B1(_0147_),
    .B2(net919),
    .X(net508));
 sky130_fd_sc_hd__mux2_1 _1086_ (.A0(net21),
    .A1(net155),
    .S(net867),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_4 _1087_ (.A1(net88),
    .A2(net845),
    .B1(_0148_),
    .B2(net919),
    .X(net513));
 sky130_fd_sc_hd__mux2_1 _1088_ (.A0(net22),
    .A1(net156),
    .S(net868),
    .X(_0149_));
 sky130_fd_sc_hd__a22o_4 _1089_ (.A1(net89),
    .A2(net845),
    .B1(_0149_),
    .B2(net920),
    .X(net514));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(net23),
    .A1(net157),
    .S(net869),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_2 _1091_ (.A1(net90),
    .A2(net845),
    .B1(_0150_),
    .B2(net920),
    .X(net515));
 sky130_fd_sc_hd__mux2_1 _1092_ (.A0(net24),
    .A1(net158),
    .S(net869),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_2 _1093_ (.A1(net91),
    .A2(net845),
    .B1(_0151_),
    .B2(net921),
    .X(net516));
 sky130_fd_sc_hd__mux2_1 _1094_ (.A0(net25),
    .A1(net159),
    .S(net869),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_1 _1095_ (.A1(net92),
    .A2(net846),
    .B1(_0152_),
    .B2(net921),
    .X(net517));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(net26),
    .A1(net160),
    .S(net869),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_1 _1097_ (.A1(net93),
    .A2(net846),
    .B1(_0153_),
    .B2(net921),
    .X(net518));
 sky130_fd_sc_hd__mux2_1 _1098_ (.A0(net27),
    .A1(net161),
    .S(net867),
    .X(_0154_));
 sky130_fd_sc_hd__a22o_2 _1099_ (.A1(net94),
    .A2(net845),
    .B1(_0154_),
    .B2(net919),
    .X(net519));
 sky130_fd_sc_hd__mux2_1 _1100_ (.A0(net28),
    .A1(net162),
    .S(net869),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_2 _1101_ (.A1(net95),
    .A2(net848),
    .B1(_0155_),
    .B2(net919),
    .X(net520));
 sky130_fd_sc_hd__mux2_1 _1102_ (.A0(net2),
    .A1(net136),
    .S(net869),
    .X(_0156_));
 sky130_fd_sc_hd__a22o_1 _1103_ (.A1(net69),
    .A2(net846),
    .B1(_0156_),
    .B2(net922),
    .X(net498));
 sky130_fd_sc_hd__mux2_1 _1104_ (.A0(net3),
    .A1(net137),
    .S(net870),
    .X(_0157_));
 sky130_fd_sc_hd__a22o_1 _1105_ (.A1(net70),
    .A2(net846),
    .B1(_0157_),
    .B2(net922),
    .X(net499));
 sky130_fd_sc_hd__mux2_1 _1106_ (.A0(net4),
    .A1(net138),
    .S(net871),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _1107_ (.A1(net71),
    .A2(net847),
    .B1(_0158_),
    .B2(net923),
    .X(net500));
 sky130_fd_sc_hd__mux2_1 _1108_ (.A0(net5),
    .A1(net139),
    .S(net871),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _1109_ (.A1(net72),
    .A2(net847),
    .B1(_0159_),
    .B2(net923),
    .X(net501));
 sky130_fd_sc_hd__mux2_1 _1110_ (.A0(net6),
    .A1(net140),
    .S(net871),
    .X(_0160_));
 sky130_fd_sc_hd__a22o_1 _1111_ (.A1(net73),
    .A2(net846),
    .B1(_0160_),
    .B2(net923),
    .X(net502));
 sky130_fd_sc_hd__mux2_1 _1112_ (.A0(net7),
    .A1(net141),
    .S(net871),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_1 _1113_ (.A1(net74),
    .A2(net847),
    .B1(_0161_),
    .B2(net923),
    .X(net503));
 sky130_fd_sc_hd__mux2_1 _1114_ (.A0(net8),
    .A1(net142),
    .S(net872),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _1115_ (.A1(net75),
    .A2(net847),
    .B1(_0162_),
    .B2(net925),
    .X(net504));
 sky130_fd_sc_hd__mux2_1 _1116_ (.A0(net9),
    .A1(net143),
    .S(net870),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_2 _1117_ (.A1(net76),
    .A2(net846),
    .B1(_0163_),
    .B2(net921),
    .X(net505));
 sky130_fd_sc_hd__mux2_1 _1118_ (.A0(net10),
    .A1(net144),
    .S(net874),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _1119_ (.A1(net77),
    .A2(net846),
    .B1(_0164_),
    .B2(net925),
    .X(net506));
 sky130_fd_sc_hd__mux2_1 _1120_ (.A0(net11),
    .A1(net145),
    .S(net871),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _1121_ (.A1(net78),
    .A2(net846),
    .B1(_0165_),
    .B2(net923),
    .X(net507));
 sky130_fd_sc_hd__mux2_1 _1122_ (.A0(net13),
    .A1(net147),
    .S(net872),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _1123_ (.A1(net80),
    .A2(net846),
    .B1(_0166_),
    .B2(net925),
    .X(net509));
 sky130_fd_sc_hd__mux2_1 _1124_ (.A0(net14),
    .A1(net148),
    .S(net872),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _1125_ (.A1(net81),
    .A2(net847),
    .B1(_0167_),
    .B2(net925),
    .X(net510));
 sky130_fd_sc_hd__mux2_1 _1126_ (.A0(net15),
    .A1(net149),
    .S(net872),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _1127_ (.A1(net82),
    .A2(net847),
    .B1(_0168_),
    .B2(net925),
    .X(net511));
 sky130_fd_sc_hd__mux2_1 _1128_ (.A0(net16),
    .A1(net150),
    .S(net872),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _1129_ (.A1(net83),
    .A2(net846),
    .B1(_0169_),
    .B2(net925),
    .X(net512));
 sky130_fd_sc_hd__nand2_8 _1130_ (.A(net925),
    .B(net872),
    .Y(_0170_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(net97),
    .A1(net30),
    .S(net919),
    .X(_0171_));
 sky130_fd_sc_hd__o22a_2 _1132_ (.A1(net164),
    .A2(net844),
    .B1(_0171_),
    .B2(net867),
    .X(net522));
 sky130_fd_sc_hd__mux2_1 _1133_ (.A0(net108),
    .A1(net41),
    .S(net920),
    .X(_0172_));
 sky130_fd_sc_hd__o22a_2 _1134_ (.A1(net175),
    .A2(net844),
    .B1(_0172_),
    .B2(net867),
    .X(net533));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(net119),
    .A1(net52),
    .S(net919),
    .X(_0173_));
 sky130_fd_sc_hd__o22a_2 _1136_ (.A1(net186),
    .A2(net844),
    .B1(_0173_),
    .B2(net867),
    .X(net544));
 sky130_fd_sc_hd__mux2_1 _1137_ (.A0(net122),
    .A1(net55),
    .S(net921),
    .X(_0174_));
 sky130_fd_sc_hd__o22a_1 _1138_ (.A1(net189),
    .A2(net844),
    .B1(_0174_),
    .B2(net869),
    .X(net547));
 sky130_fd_sc_hd__mux2_1 _1139_ (.A0(net123),
    .A1(net56),
    .S(net922),
    .X(_0175_));
 sky130_fd_sc_hd__o22a_1 _1140_ (.A1(net190),
    .A2(net844),
    .B1(_0175_),
    .B2(net870),
    .X(net548));
 sky130_fd_sc_hd__mux2_1 _1141_ (.A0(net124),
    .A1(net57),
    .S(net922),
    .X(_0176_));
 sky130_fd_sc_hd__o22a_1 _1142_ (.A1(net191),
    .A2(net844),
    .B1(_0176_),
    .B2(net870),
    .X(net549));
 sky130_fd_sc_hd__mux2_1 _1143_ (.A0(net125),
    .A1(net58),
    .S(net922),
    .X(_0177_));
 sky130_fd_sc_hd__o22a_1 _1144_ (.A1(net192),
    .A2(net843),
    .B1(_0177_),
    .B2(net870),
    .X(net550));
 sky130_fd_sc_hd__mux2_1 _1145_ (.A0(net126),
    .A1(net59),
    .S(net922),
    .X(_0178_));
 sky130_fd_sc_hd__o22a_1 _1146_ (.A1(net193),
    .A2(net843),
    .B1(_0178_),
    .B2(net870),
    .X(net551));
 sky130_fd_sc_hd__mux2_1 _1147_ (.A0(net127),
    .A1(net60),
    .S(net921),
    .X(_0179_));
 sky130_fd_sc_hd__o22a_1 _1148_ (.A1(net194),
    .A2(net843),
    .B1(_0179_),
    .B2(net871),
    .X(net552));
 sky130_fd_sc_hd__mux2_1 _1149_ (.A0(net128),
    .A1(net61),
    .S(net921),
    .X(_0180_));
 sky130_fd_sc_hd__o22a_1 _1150_ (.A1(net195),
    .A2(net843),
    .B1(_0180_),
    .B2(net870),
    .X(net553));
 sky130_fd_sc_hd__mux2_1 _1151_ (.A0(net98),
    .A1(net31),
    .S(net923),
    .X(_0181_));
 sky130_fd_sc_hd__o22a_1 _1152_ (.A1(net165),
    .A2(net843),
    .B1(_0181_),
    .B2(net871),
    .X(net523));
 sky130_fd_sc_hd__mux2_1 _1153_ (.A0(net99),
    .A1(net32),
    .S(net923),
    .X(_0182_));
 sky130_fd_sc_hd__o22a_1 _1154_ (.A1(net166),
    .A2(net843),
    .B1(_0182_),
    .B2(net871),
    .X(net524));
 sky130_fd_sc_hd__mux2_1 _1155_ (.A0(net100),
    .A1(net33),
    .S(net923),
    .X(_0183_));
 sky130_fd_sc_hd__o22a_1 _1156_ (.A1(net167),
    .A2(net842),
    .B1(_0183_),
    .B2(net871),
    .X(net525));
 sky130_fd_sc_hd__mux2_1 _1157_ (.A0(net101),
    .A1(net34),
    .S(net923),
    .X(_0184_));
 sky130_fd_sc_hd__o22a_1 _1158_ (.A1(net168),
    .A2(net843),
    .B1(_0184_),
    .B2(net875),
    .X(net526));
 sky130_fd_sc_hd__mux2_1 _1159_ (.A0(net102),
    .A1(net35),
    .S(net924),
    .X(_0185_));
 sky130_fd_sc_hd__o22a_1 _1160_ (.A1(net169),
    .A2(net842),
    .B1(_0185_),
    .B2(net874),
    .X(net527));
 sky130_fd_sc_hd__mux2_1 _1161_ (.A0(net103),
    .A1(net36),
    .S(net924),
    .X(_0186_));
 sky130_fd_sc_hd__o22a_1 _1162_ (.A1(net170),
    .A2(net842),
    .B1(_0186_),
    .B2(net874),
    .X(net528));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(net104),
    .A1(net37),
    .S(net924),
    .X(_0187_));
 sky130_fd_sc_hd__o22a_1 _1164_ (.A1(net171),
    .A2(net842),
    .B1(_0187_),
    .B2(net874),
    .X(net529));
 sky130_fd_sc_hd__mux2_1 _1165_ (.A0(net105),
    .A1(net38),
    .S(net924),
    .X(_0188_));
 sky130_fd_sc_hd__o22a_1 _1166_ (.A1(net172),
    .A2(net842),
    .B1(_0188_),
    .B2(net872),
    .X(net530));
 sky130_fd_sc_hd__mux2_1 _1167_ (.A0(net106),
    .A1(net39),
    .S(net925),
    .X(_0189_));
 sky130_fd_sc_hd__o22a_1 _1168_ (.A1(net173),
    .A2(_0170_),
    .B1(_0189_),
    .B2(net872),
    .X(net531));
 sky130_fd_sc_hd__mux2_1 _1169_ (.A0(net107),
    .A1(net40),
    .S(net926),
    .X(_0190_));
 sky130_fd_sc_hd__o22a_2 _1170_ (.A1(net174),
    .A2(net843),
    .B1(_0190_),
    .B2(net875),
    .X(net532));
 sky130_fd_sc_hd__mux2_1 _1171_ (.A0(net109),
    .A1(net42),
    .S(net924),
    .X(_0191_));
 sky130_fd_sc_hd__o22a_1 _1172_ (.A1(net176),
    .A2(_0170_),
    .B1(_0191_),
    .B2(net872),
    .X(net534));
 sky130_fd_sc_hd__mux2_2 _1173_ (.A0(net110),
    .A1(net43),
    .S(net923),
    .X(_0192_));
 sky130_fd_sc_hd__o22a_1 _1174_ (.A1(net177),
    .A2(_0170_),
    .B1(_0192_),
    .B2(net873),
    .X(net535));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(net111),
    .A1(net44),
    .S(net924),
    .X(_0193_));
 sky130_fd_sc_hd__o22a_1 _1176_ (.A1(net178),
    .A2(net842),
    .B1(_0193_),
    .B2(net873),
    .X(net536));
 sky130_fd_sc_hd__mux2_1 _1177_ (.A0(net112),
    .A1(net45),
    .S(net924),
    .X(_0194_));
 sky130_fd_sc_hd__o22a_1 _1178_ (.A1(net179),
    .A2(net842),
    .B1(_0194_),
    .B2(net872),
    .X(net537));
 sky130_fd_sc_hd__mux2_1 _1179_ (.A0(net113),
    .A1(net46),
    .S(net924),
    .X(_0195_));
 sky130_fd_sc_hd__o22a_1 _1180_ (.A1(net180),
    .A2(net842),
    .B1(_0195_),
    .B2(net873),
    .X(net538));
 sky130_fd_sc_hd__mux2_1 _1181_ (.A0(net114),
    .A1(net47),
    .S(net921),
    .X(_0196_));
 sky130_fd_sc_hd__o22a_4 _1182_ (.A1(net181),
    .A2(net844),
    .B1(_0196_),
    .B2(net869),
    .X(net539));
 sky130_fd_sc_hd__mux2_1 _1183_ (.A0(net115),
    .A1(net48),
    .S(net924),
    .X(_0197_));
 sky130_fd_sc_hd__o22a_1 _1184_ (.A1(net182),
    .A2(net842),
    .B1(_0197_),
    .B2(net873),
    .X(net540));
 sky130_fd_sc_hd__mux2_1 _1185_ (.A0(net116),
    .A1(net49),
    .S(net924),
    .X(_0198_));
 sky130_fd_sc_hd__o22a_1 _1186_ (.A1(net183),
    .A2(net842),
    .B1(_0198_),
    .B2(net873),
    .X(net541));
 sky130_fd_sc_hd__mux2_1 _1187_ (.A0(net117),
    .A1(net50),
    .S(net921),
    .X(_0199_));
 sky130_fd_sc_hd__o22a_4 _1188_ (.A1(net184),
    .A2(net844),
    .B1(_0199_),
    .B2(net869),
    .X(net542));
 sky130_fd_sc_hd__mux2_1 _1189_ (.A0(net118),
    .A1(net51),
    .S(net920),
    .X(_0200_));
 sky130_fd_sc_hd__o22a_4 _1190_ (.A1(net185),
    .A2(net844),
    .B1(_0200_),
    .B2(net868),
    .X(net543));
 sky130_fd_sc_hd__mux2_1 _1191_ (.A0(net120),
    .A1(net53),
    .S(net926),
    .X(_0201_));
 sky130_fd_sc_hd__o22a_2 _1192_ (.A1(net187),
    .A2(net843),
    .B1(_0201_),
    .B2(net871),
    .X(net545));
 sky130_fd_sc_hd__mux2_1 _1193_ (.A0(net121),
    .A1(net54),
    .S(net921),
    .X(_0202_));
 sky130_fd_sc_hd__o22a_4 _1194_ (.A1(net188),
    .A2(net844),
    .B1(_0202_),
    .B2(net869),
    .X(net546));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(net62),
    .A1(net196),
    .S(net868),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_4 _1196_ (.A1(net129),
    .A2(net845),
    .B1(_0203_),
    .B2(net920),
    .X(net554));
 sky130_fd_sc_hd__mux2_1 _1197_ (.A0(net63),
    .A1(net197),
    .S(net868),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_4 _1198_ (.A1(net130),
    .A2(net845),
    .B1(_0204_),
    .B2(net920),
    .X(net555));
 sky130_fd_sc_hd__mux2_1 _1199_ (.A0(net64),
    .A1(net198),
    .S(net868),
    .X(_0205_));
 sky130_fd_sc_hd__a22o_4 _1200_ (.A1(net131),
    .A2(net845),
    .B1(_0205_),
    .B2(net920),
    .X(net556));
 sky130_fd_sc_hd__mux2_1 _1201_ (.A0(net65),
    .A1(net199),
    .S(net868),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_2 _1202_ (.A1(net132),
    .A2(net848),
    .B1(_0206_),
    .B2(net920),
    .X(net557));
 sky130_fd_sc_hd__mux2_1 _1203_ (.A0(net67),
    .A1(net201),
    .S(net867),
    .X(_0207_));
 sky130_fd_sc_hd__a22o_2 _1204_ (.A1(net134),
    .A2(net848),
    .B1(_0207_),
    .B2(net919),
    .X(net559));
 sky130_fd_sc_hd__mux2_1 _1205_ (.A0(net66),
    .A1(net200),
    .S(net867),
    .X(_0208_));
 sky130_fd_sc_hd__a22o_2 _1206_ (.A1(net133),
    .A2(net845),
    .B1(_0208_),
    .B2(net919),
    .X(net558));
 sky130_fd_sc_hd__a221o_4 _1207_ (.A1(net1006),
    .A2(_0641_),
    .B1(net957),
    .B2(net1009),
    .C1(_0651_),
    .X(net521));
 sky130_fd_sc_hd__nor2_1 _1208_ (.A(net927),
    .B(net911),
    .Y(_0209_));
 sky130_fd_sc_hd__mux2_1 _1209_ (.A0(net1),
    .A1(net135),
    .S(net913),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_1 _1210_ (.A1(net68),
    .A2(net838),
    .B1(_0210_),
    .B2(net928),
    .X(net560));
 sky130_fd_sc_hd__mux2_1 _1211_ (.A0(net12),
    .A1(net146),
    .S(net911),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _1212_ (.A1(net79),
    .A2(net838),
    .B1(_0211_),
    .B2(net928),
    .X(net571));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(net21),
    .A1(net155),
    .S(net911),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_2 _1214_ (.A1(net88),
    .A2(net838),
    .B1(_0212_),
    .B2(net927),
    .X(net576));
 sky130_fd_sc_hd__mux2_1 _1215_ (.A0(net22),
    .A1(net156),
    .S(net911),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_2 _1216_ (.A1(net89),
    .A2(net838),
    .B1(_0213_),
    .B2(net927),
    .X(net577));
 sky130_fd_sc_hd__mux2_1 _1217_ (.A0(net23),
    .A1(net157),
    .S(net913),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_1 _1218_ (.A1(net90),
    .A2(net841),
    .B1(_0214_),
    .B2(net929),
    .X(net578));
 sky130_fd_sc_hd__mux2_1 _1219_ (.A0(net24),
    .A1(net158),
    .S(net913),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _1220_ (.A1(net91),
    .A2(net841),
    .B1(_0215_),
    .B2(net929),
    .X(net579));
 sky130_fd_sc_hd__mux2_1 _1221_ (.A0(net25),
    .A1(net159),
    .S(net914),
    .X(_0216_));
 sky130_fd_sc_hd__a22o_1 _1222_ (.A1(net92),
    .A2(net838),
    .B1(_0216_),
    .B2(net929),
    .X(net580));
 sky130_fd_sc_hd__mux2_1 _1223_ (.A0(net26),
    .A1(net160),
    .S(net914),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _1224_ (.A1(net93),
    .A2(net839),
    .B1(_0217_),
    .B2(net929),
    .X(net581));
 sky130_fd_sc_hd__mux2_1 _1225_ (.A0(net27),
    .A1(net161),
    .S(net914),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _1226_ (.A1(net94),
    .A2(net839),
    .B1(_0218_),
    .B2(net929),
    .X(net582));
 sky130_fd_sc_hd__mux2_1 _1227_ (.A0(net28),
    .A1(net162),
    .S(net914),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_1 _1228_ (.A1(net95),
    .A2(net839),
    .B1(_0219_),
    .B2(net929),
    .X(net583));
 sky130_fd_sc_hd__mux2_1 _1229_ (.A0(net2),
    .A1(net136),
    .S(net914),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _1230_ (.A1(net69),
    .A2(net839),
    .B1(_0220_),
    .B2(net929),
    .X(net561));
 sky130_fd_sc_hd__mux2_1 _1231_ (.A0(net3),
    .A1(net137),
    .S(net914),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_1 _1232_ (.A1(net70),
    .A2(net839),
    .B1(_0221_),
    .B2(net930),
    .X(net562));
 sky130_fd_sc_hd__mux2_1 _1233_ (.A0(net4),
    .A1(net138),
    .S(net915),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _1234_ (.A1(net71),
    .A2(net839),
    .B1(_0222_),
    .B2(net930),
    .X(net563));
 sky130_fd_sc_hd__mux2_1 _1235_ (.A0(net5),
    .A1(net139),
    .S(net915),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_1 _1236_ (.A1(net72),
    .A2(net839),
    .B1(_0223_),
    .B2(net930),
    .X(net564));
 sky130_fd_sc_hd__mux2_1 _1237_ (.A0(net6),
    .A1(net140),
    .S(net915),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_1 _1238_ (.A1(net73),
    .A2(net839),
    .B1(_0224_),
    .B2(net930),
    .X(net565));
 sky130_fd_sc_hd__mux2_1 _1239_ (.A0(net7),
    .A1(net141),
    .S(net915),
    .X(_0225_));
 sky130_fd_sc_hd__a22o_1 _1240_ (.A1(net74),
    .A2(net840),
    .B1(_0225_),
    .B2(net930),
    .X(net566));
 sky130_fd_sc_hd__mux2_1 _1241_ (.A0(net8),
    .A1(net142),
    .S(net918),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_1 _1242_ (.A1(net75),
    .A2(net839),
    .B1(_0226_),
    .B2(net932),
    .X(net567));
 sky130_fd_sc_hd__mux2_1 _1243_ (.A0(net9),
    .A1(net143),
    .S(net916),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_1 _1244_ (.A1(net76),
    .A2(net840),
    .B1(_0227_),
    .B2(net932),
    .X(net568));
 sky130_fd_sc_hd__mux2_1 _1245_ (.A0(net10),
    .A1(net144),
    .S(net915),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_1 _1246_ (.A1(net77),
    .A2(net840),
    .B1(_0228_),
    .B2(net932),
    .X(net569));
 sky130_fd_sc_hd__mux2_1 _1247_ (.A0(net11),
    .A1(net145),
    .S(net916),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_1 _1248_ (.A1(net78),
    .A2(net839),
    .B1(_0229_),
    .B2(net932),
    .X(net570));
 sky130_fd_sc_hd__mux2_1 _1249_ (.A0(net13),
    .A1(net147),
    .S(net916),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _1250_ (.A1(net80),
    .A2(net840),
    .B1(_0230_),
    .B2(net932),
    .X(net572));
 sky130_fd_sc_hd__mux2_1 _1251_ (.A0(net14),
    .A1(net148),
    .S(net916),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _1252_ (.A1(net81),
    .A2(net840),
    .B1(_0231_),
    .B2(net932),
    .X(net573));
 sky130_fd_sc_hd__mux2_1 _1253_ (.A0(net15),
    .A1(net149),
    .S(net916),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _1254_ (.A1(net82),
    .A2(net840),
    .B1(_0232_),
    .B2(net932),
    .X(net574));
 sky130_fd_sc_hd__mux2_1 _1255_ (.A0(net16),
    .A1(net150),
    .S(net916),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _1256_ (.A1(net83),
    .A2(net840),
    .B1(_0233_),
    .B2(net932),
    .X(net575));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(net927),
    .B(net911),
    .Y(_0234_));
 sky130_fd_sc_hd__mux2_1 _1258_ (.A0(net97),
    .A1(net30),
    .S(net928),
    .X(_0235_));
 sky130_fd_sc_hd__o22a_1 _1259_ (.A1(net164),
    .A2(net834),
    .B1(_0235_),
    .B2(net911),
    .X(net585));
 sky130_fd_sc_hd__mux2_1 _1260_ (.A0(net108),
    .A1(net41),
    .S(net927),
    .X(_0236_));
 sky130_fd_sc_hd__o22a_2 _1261_ (.A1(net175),
    .A2(net834),
    .B1(_0236_),
    .B2(net911),
    .X(net596));
 sky130_fd_sc_hd__mux2_1 _1262_ (.A0(net119),
    .A1(net52),
    .S(net927),
    .X(_0237_));
 sky130_fd_sc_hd__o22a_2 _1263_ (.A1(net186),
    .A2(net834),
    .B1(_0237_),
    .B2(net911),
    .X(net607));
 sky130_fd_sc_hd__mux2_1 _1264_ (.A0(net122),
    .A1(net55),
    .S(net927),
    .X(_0238_));
 sky130_fd_sc_hd__o22a_2 _1265_ (.A1(net189),
    .A2(net834),
    .B1(_0238_),
    .B2(net911),
    .X(net610));
 sky130_fd_sc_hd__mux2_1 _1266_ (.A0(net123),
    .A1(net56),
    .S(net927),
    .X(_0239_));
 sky130_fd_sc_hd__o22a_2 _1267_ (.A1(net190),
    .A2(net834),
    .B1(_0239_),
    .B2(net912),
    .X(net611));
 sky130_fd_sc_hd__mux2_1 _1268_ (.A0(net124),
    .A1(net57),
    .S(net928),
    .X(_0240_));
 sky130_fd_sc_hd__o22a_2 _1269_ (.A1(net191),
    .A2(net834),
    .B1(_0240_),
    .B2(net913),
    .X(net612));
 sky130_fd_sc_hd__mux2_1 _1270_ (.A0(net125),
    .A1(net58),
    .S(net928),
    .X(_0241_));
 sky130_fd_sc_hd__o22a_2 _1271_ (.A1(net192),
    .A2(net834),
    .B1(_0241_),
    .B2(net913),
    .X(net613));
 sky130_fd_sc_hd__mux2_1 _1272_ (.A0(net126),
    .A1(net59),
    .S(net931),
    .X(_0242_));
 sky130_fd_sc_hd__o22a_1 _1273_ (.A1(net193),
    .A2(net834),
    .B1(_0242_),
    .B2(net913),
    .X(net614));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(net127),
    .A1(net60),
    .S(net928),
    .X(_0243_));
 sky130_fd_sc_hd__o22a_2 _1275_ (.A1(net194),
    .A2(net834),
    .B1(_0243_),
    .B2(net912),
    .X(net615));
 sky130_fd_sc_hd__mux2_1 _1276_ (.A0(net128),
    .A1(net61),
    .S(net929),
    .X(_0244_));
 sky130_fd_sc_hd__o22a_2 _1277_ (.A1(net195),
    .A2(net837),
    .B1(_0244_),
    .B2(net913),
    .X(net616));
 sky130_fd_sc_hd__mux2_1 _1278_ (.A0(net98),
    .A1(net31),
    .S(net929),
    .X(_0245_));
 sky130_fd_sc_hd__o22a_2 _1279_ (.A1(net165),
    .A2(net834),
    .B1(_0245_),
    .B2(net914),
    .X(net586));
 sky130_fd_sc_hd__mux2_1 _1280_ (.A0(net99),
    .A1(net32),
    .S(net931),
    .X(_0246_));
 sky130_fd_sc_hd__o22a_1 _1281_ (.A1(net166),
    .A2(net837),
    .B1(_0246_),
    .B2(net914),
    .X(net587));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(net100),
    .A1(net33),
    .S(net929),
    .X(_0247_));
 sky130_fd_sc_hd__o22a_1 _1283_ (.A1(net167),
    .A2(net836),
    .B1(_0247_),
    .B2(net914),
    .X(net588));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(net101),
    .A1(net34),
    .S(net931),
    .X(_0248_));
 sky130_fd_sc_hd__o22a_1 _1285_ (.A1(net168),
    .A2(net836),
    .B1(_0248_),
    .B2(net915),
    .X(net589));
 sky130_fd_sc_hd__mux2_1 _1286_ (.A0(net102),
    .A1(net35),
    .S(net930),
    .X(_0249_));
 sky130_fd_sc_hd__o22a_1 _1287_ (.A1(net169),
    .A2(net836),
    .B1(_0249_),
    .B2(net915),
    .X(net590));
 sky130_fd_sc_hd__mux2_1 _1288_ (.A0(net103),
    .A1(net36),
    .S(net930),
    .X(_0250_));
 sky130_fd_sc_hd__o22a_1 _1289_ (.A1(net170),
    .A2(net836),
    .B1(_0250_),
    .B2(net915),
    .X(net591));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(net104),
    .A1(net37),
    .S(net931),
    .X(_0251_));
 sky130_fd_sc_hd__o22a_1 _1291_ (.A1(net171),
    .A2(net836),
    .B1(_0251_),
    .B2(net915),
    .X(net592));
 sky130_fd_sc_hd__mux2_1 _1292_ (.A0(net105),
    .A1(net38),
    .S(net930),
    .X(_0252_));
 sky130_fd_sc_hd__o22a_1 _1293_ (.A1(net172),
    .A2(net836),
    .B1(_0252_),
    .B2(net915),
    .X(net593));
 sky130_fd_sc_hd__mux2_1 _1294_ (.A0(net106),
    .A1(net39),
    .S(net930),
    .X(_0253_));
 sky130_fd_sc_hd__o22a_1 _1295_ (.A1(net173),
    .A2(net836),
    .B1(_0253_),
    .B2(net918),
    .X(net594));
 sky130_fd_sc_hd__mux2_1 _1296_ (.A0(net107),
    .A1(net40),
    .S(net933),
    .X(_0254_));
 sky130_fd_sc_hd__o22a_2 _1297_ (.A1(net174),
    .A2(net836),
    .B1(_0254_),
    .B2(net916),
    .X(net595));
 sky130_fd_sc_hd__mux2_2 _1298_ (.A0(net109),
    .A1(net42),
    .S(net933),
    .X(_0255_));
 sky130_fd_sc_hd__o22a_1 _1299_ (.A1(net176),
    .A2(net835),
    .B1(_0255_),
    .B2(net917),
    .X(net597));
 sky130_fd_sc_hd__mux2_1 _1300_ (.A0(net110),
    .A1(net43),
    .S(net930),
    .X(_0256_));
 sky130_fd_sc_hd__o22a_1 _1301_ (.A1(net177),
    .A2(net837),
    .B1(_0256_),
    .B2(net918),
    .X(net598));
 sky130_fd_sc_hd__mux2_1 _1302_ (.A0(net111),
    .A1(net44),
    .S(net932),
    .X(_0257_));
 sky130_fd_sc_hd__o22a_1 _1303_ (.A1(net178),
    .A2(net835),
    .B1(_0257_),
    .B2(net918),
    .X(net599));
 sky130_fd_sc_hd__mux2_1 _1304_ (.A0(net112),
    .A1(net45),
    .S(net932),
    .X(_0258_));
 sky130_fd_sc_hd__o22a_1 _1305_ (.A1(net179),
    .A2(net835),
    .B1(_0258_),
    .B2(net918),
    .X(net600));
 sky130_fd_sc_hd__mux2_1 _1306_ (.A0(net113),
    .A1(net46),
    .S(net933),
    .X(_0259_));
 sky130_fd_sc_hd__o22a_1 _1307_ (.A1(net180),
    .A2(net835),
    .B1(_0259_),
    .B2(net917),
    .X(net601));
 sky130_fd_sc_hd__mux2_1 _1308_ (.A0(net114),
    .A1(net47),
    .S(net933),
    .X(_0260_));
 sky130_fd_sc_hd__o22a_1 _1309_ (.A1(net181),
    .A2(net835),
    .B1(_0260_),
    .B2(net916),
    .X(net602));
 sky130_fd_sc_hd__mux2_1 _1310_ (.A0(net115),
    .A1(net48),
    .S(net934),
    .X(_0261_));
 sky130_fd_sc_hd__o22a_1 _1311_ (.A1(net182),
    .A2(net836),
    .B1(_0261_),
    .B2(net916),
    .X(net603));
 sky130_fd_sc_hd__mux2_1 _1312_ (.A0(net116),
    .A1(net49),
    .S(net933),
    .X(_0262_));
 sky130_fd_sc_hd__o22a_1 _1313_ (.A1(net183),
    .A2(net835),
    .B1(_0262_),
    .B2(net917),
    .X(net604));
 sky130_fd_sc_hd__mux2_1 _1314_ (.A0(net117),
    .A1(net50),
    .S(net933),
    .X(_0263_));
 sky130_fd_sc_hd__o22a_1 _1315_ (.A1(net184),
    .A2(net835),
    .B1(_0263_),
    .B2(net917),
    .X(net605));
 sky130_fd_sc_hd__mux2_1 _1316_ (.A0(net118),
    .A1(net51),
    .S(net933),
    .X(_0264_));
 sky130_fd_sc_hd__o22a_1 _1317_ (.A1(net185),
    .A2(net835),
    .B1(_0264_),
    .B2(net916),
    .X(net606));
 sky130_fd_sc_hd__mux2_1 _1318_ (.A0(net120),
    .A1(net53),
    .S(net933),
    .X(_0265_));
 sky130_fd_sc_hd__o22a_1 _1319_ (.A1(net187),
    .A2(net835),
    .B1(_0265_),
    .B2(net917),
    .X(net608));
 sky130_fd_sc_hd__mux2_2 _1320_ (.A0(net121),
    .A1(net54),
    .S(net933),
    .X(_0266_));
 sky130_fd_sc_hd__o22a_1 _1321_ (.A1(net188),
    .A2(net835),
    .B1(_0266_),
    .B2(net917),
    .X(net609));
 sky130_fd_sc_hd__mux2_1 _1322_ (.A0(net62),
    .A1(net196),
    .S(net913),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _1323_ (.A1(net129),
    .A2(net838),
    .B1(_0267_),
    .B2(net928),
    .X(net617));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(net63),
    .A1(net197),
    .S(net911),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_2 _1325_ (.A1(net130),
    .A2(net838),
    .B1(_0268_),
    .B2(net927),
    .X(net618));
 sky130_fd_sc_hd__mux2_1 _1326_ (.A0(net64),
    .A1(net198),
    .S(net913),
    .X(_0269_));
 sky130_fd_sc_hd__a22o_1 _1327_ (.A1(net131),
    .A2(net841),
    .B1(_0269_),
    .B2(net928),
    .X(net619));
 sky130_fd_sc_hd__mux2_1 _1328_ (.A0(net65),
    .A1(net199),
    .S(net913),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _1329_ (.A1(net132),
    .A2(net838),
    .B1(_0270_),
    .B2(net928),
    .X(net620));
 sky130_fd_sc_hd__mux2_1 _1330_ (.A0(net67),
    .A1(net201),
    .S(net912),
    .X(_0271_));
 sky130_fd_sc_hd__a22o_1 _1331_ (.A1(net134),
    .A2(net838),
    .B1(_0271_),
    .B2(net928),
    .X(net622));
 sky130_fd_sc_hd__mux2_1 _1332_ (.A0(net66),
    .A1(net200),
    .S(net912),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _1333_ (.A1(net133),
    .A2(net838),
    .B1(_0272_),
    .B2(net927),
    .X(net621));
 sky130_fd_sc_hd__a221o_4 _1334_ (.A1(net96),
    .A2(_0597_),
    .B1(net997),
    .B2(net163),
    .C1(_0607_),
    .X(net584));
 sky130_fd_sc_hd__nor2_8 _1335_ (.A(net904),
    .B(net895),
    .Y(_0273_));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(net1),
    .A1(net135),
    .S(net902),
    .X(_0274_));
 sky130_fd_sc_hd__a22o_4 _1337_ (.A1(net68),
    .A2(net833),
    .B1(_0274_),
    .B2(net894),
    .X(net623));
 sky130_fd_sc_hd__mux2_1 _1338_ (.A0(net12),
    .A1(net146),
    .S(net902),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_4 _1339_ (.A1(net79),
    .A2(net833),
    .B1(_0275_),
    .B2(net893),
    .X(net634));
 sky130_fd_sc_hd__mux2_1 _1340_ (.A0(net21),
    .A1(net155),
    .S(net902),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_4 _1341_ (.A1(net88),
    .A2(net833),
    .B1(_0276_),
    .B2(net894),
    .X(net639));
 sky130_fd_sc_hd__mux2_1 _1342_ (.A0(net22),
    .A1(net156),
    .S(net902),
    .X(_0277_));
 sky130_fd_sc_hd__a22o_4 _1343_ (.A1(net89),
    .A2(net833),
    .B1(_0277_),
    .B2(net893),
    .X(net640));
 sky130_fd_sc_hd__mux2_1 _1344_ (.A0(net23),
    .A1(net157),
    .S(net909),
    .X(_0278_));
 sky130_fd_sc_hd__a22o_4 _1345_ (.A1(net90),
    .A2(net832),
    .B1(_0278_),
    .B2(net901),
    .X(net641));
 sky130_fd_sc_hd__mux2_1 _1346_ (.A0(net24),
    .A1(net158),
    .S(net903),
    .X(_0279_));
 sky130_fd_sc_hd__a22o_2 _1347_ (.A1(net91),
    .A2(net832),
    .B1(_0279_),
    .B2(net897),
    .X(net642));
 sky130_fd_sc_hd__mux2_1 _1348_ (.A0(net25),
    .A1(net159),
    .S(net903),
    .X(_0280_));
 sky130_fd_sc_hd__a22o_1 _1349_ (.A1(net92),
    .A2(net832),
    .B1(_0280_),
    .B2(net897),
    .X(net643));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(net26),
    .A1(net160),
    .S(net903),
    .X(_0281_));
 sky130_fd_sc_hd__a22o_1 _1351_ (.A1(net93),
    .A2(net832),
    .B1(_0281_),
    .B2(net895),
    .X(net644));
 sky130_fd_sc_hd__mux2_1 _1352_ (.A0(net27),
    .A1(net161),
    .S(net903),
    .X(_0282_));
 sky130_fd_sc_hd__a22o_2 _1353_ (.A1(net94),
    .A2(net832),
    .B1(_0282_),
    .B2(net896),
    .X(net645));
 sky130_fd_sc_hd__mux2_1 _1354_ (.A0(net28),
    .A1(net162),
    .S(net903),
    .X(_0283_));
 sky130_fd_sc_hd__a22o_2 _1355_ (.A1(net95),
    .A2(net832),
    .B1(_0283_),
    .B2(net895),
    .X(net646));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(net2),
    .A1(net136),
    .S(net903),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_2 _1357_ (.A1(net69),
    .A2(net832),
    .B1(_0284_),
    .B2(net896),
    .X(net624));
 sky130_fd_sc_hd__mux2_1 _1358_ (.A0(net3),
    .A1(net137),
    .S(net903),
    .X(_0285_));
 sky130_fd_sc_hd__a22o_2 _1359_ (.A1(net70),
    .A2(net832),
    .B1(_0285_),
    .B2(net896),
    .X(net625));
 sky130_fd_sc_hd__mux2_1 _1360_ (.A0(net4),
    .A1(net138),
    .S(net903),
    .X(_0286_));
 sky130_fd_sc_hd__a22o_1 _1361_ (.A1(net71),
    .A2(net831),
    .B1(_0286_),
    .B2(net895),
    .X(net626));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(net5),
    .A1(net139),
    .S(net904),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_1 _1363_ (.A1(net72),
    .A2(net831),
    .B1(_0287_),
    .B2(net896),
    .X(net627));
 sky130_fd_sc_hd__mux2_1 _1364_ (.A0(net6),
    .A1(net140),
    .S(net903),
    .X(_0288_));
 sky130_fd_sc_hd__a22o_2 _1365_ (.A1(net73),
    .A2(net831),
    .B1(_0288_),
    .B2(net898),
    .X(net628));
 sky130_fd_sc_hd__mux2_1 _1366_ (.A0(net7),
    .A1(net141),
    .S(net907),
    .X(_0289_));
 sky130_fd_sc_hd__a22o_2 _1367_ (.A1(net74),
    .A2(net831),
    .B1(_0289_),
    .B2(net898),
    .X(net629));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(net8),
    .A1(net142),
    .S(net905),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_1 _1369_ (.A1(net75),
    .A2(net831),
    .B1(_0290_),
    .B2(net898),
    .X(net630));
 sky130_fd_sc_hd__mux2_1 _1370_ (.A0(net9),
    .A1(net143),
    .S(net909),
    .X(_0291_));
 sky130_fd_sc_hd__a22o_2 _1371_ (.A1(net76),
    .A2(_0273_),
    .B1(_0291_),
    .B2(net900),
    .X(net631));
 sky130_fd_sc_hd__mux2_1 _1372_ (.A0(net10),
    .A1(net144),
    .S(net907),
    .X(_0292_));
 sky130_fd_sc_hd__a22o_2 _1373_ (.A1(net77),
    .A2(net831),
    .B1(_0292_),
    .B2(net898),
    .X(net632));
 sky130_fd_sc_hd__mux2_1 _1374_ (.A0(net11),
    .A1(net145),
    .S(net907),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_2 _1375_ (.A1(net78),
    .A2(net831),
    .B1(_0293_),
    .B2(net898),
    .X(net633));
 sky130_fd_sc_hd__mux2_1 _1376_ (.A0(net13),
    .A1(net147),
    .S(net905),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_1 _1377_ (.A1(net80),
    .A2(net831),
    .B1(_0294_),
    .B2(net898),
    .X(net635));
 sky130_fd_sc_hd__mux2_1 _1378_ (.A0(net14),
    .A1(net148),
    .S(net905),
    .X(_0295_));
 sky130_fd_sc_hd__a22o_1 _1379_ (.A1(net81),
    .A2(net831),
    .B1(_0295_),
    .B2(net899),
    .X(net636));
 sky130_fd_sc_hd__mux2_1 _1380_ (.A0(net15),
    .A1(net149),
    .S(net905),
    .X(_0296_));
 sky130_fd_sc_hd__a22o_1 _1381_ (.A1(net82),
    .A2(net831),
    .B1(_0296_),
    .B2(net899),
    .X(net637));
 sky130_fd_sc_hd__mux2_1 _1382_ (.A0(net16),
    .A1(net150),
    .S(net906),
    .X(_0297_));
 sky130_fd_sc_hd__a22o_1 _1383_ (.A1(net83),
    .A2(net832),
    .B1(_0297_),
    .B2(net899),
    .X(net638));
 sky130_fd_sc_hd__nand2_1 _1384_ (.A(net904),
    .B(net895),
    .Y(_0298_));
 sky130_fd_sc_hd__mux2_1 _1385_ (.A0(net97),
    .A1(net30),
    .S(net893),
    .X(_0299_));
 sky130_fd_sc_hd__o22a_4 _1386_ (.A1(net164),
    .A2(net830),
    .B1(_0299_),
    .B2(net902),
    .X(net648));
 sky130_fd_sc_hd__mux2_1 _1387_ (.A0(net108),
    .A1(net41),
    .S(net893),
    .X(_0300_));
 sky130_fd_sc_hd__o22a_4 _1388_ (.A1(net175),
    .A2(net830),
    .B1(_0300_),
    .B2(net902),
    .X(net659));
 sky130_fd_sc_hd__mux2_1 _1389_ (.A0(net119),
    .A1(net52),
    .S(net893),
    .X(_0301_));
 sky130_fd_sc_hd__o22a_4 _1390_ (.A1(net186),
    .A2(net830),
    .B1(_0301_),
    .B2(net910),
    .X(net670));
 sky130_fd_sc_hd__mux2_1 _1391_ (.A0(net122),
    .A1(net55),
    .S(net901),
    .X(_0302_));
 sky130_fd_sc_hd__o22a_4 _1392_ (.A1(net189),
    .A2(net830),
    .B1(_0302_),
    .B2(net909),
    .X(net673));
 sky130_fd_sc_hd__mux2_1 _1393_ (.A0(net123),
    .A1(net56),
    .S(net897),
    .X(_0303_));
 sky130_fd_sc_hd__o22a_2 _1394_ (.A1(net190),
    .A2(net827),
    .B1(_0303_),
    .B2(net903),
    .X(net674));
 sky130_fd_sc_hd__mux2_1 _1395_ (.A0(net124),
    .A1(net57),
    .S(net897),
    .X(_0304_));
 sky130_fd_sc_hd__o22a_1 _1396_ (.A1(net191),
    .A2(net827),
    .B1(_0304_),
    .B2(net904),
    .X(net675));
 sky130_fd_sc_hd__mux2_1 _1397_ (.A0(net125),
    .A1(net58),
    .S(net895),
    .X(_0305_));
 sky130_fd_sc_hd__o22a_1 _1398_ (.A1(net192),
    .A2(net827),
    .B1(_0305_),
    .B2(net904),
    .X(net676));
 sky130_fd_sc_hd__mux2_1 _1399_ (.A0(net126),
    .A1(net59),
    .S(net895),
    .X(_0306_));
 sky130_fd_sc_hd__o22a_1 _1400_ (.A1(net193),
    .A2(net827),
    .B1(_0306_),
    .B2(net904),
    .X(net677));
 sky130_fd_sc_hd__mux2_1 _1401_ (.A0(net127),
    .A1(net60),
    .S(net895),
    .X(_0307_));
 sky130_fd_sc_hd__o22a_1 _1402_ (.A1(net194),
    .A2(net827),
    .B1(_0307_),
    .B2(net904),
    .X(net678));
 sky130_fd_sc_hd__mux2_1 _1403_ (.A0(net128),
    .A1(net61),
    .S(net896),
    .X(_0308_));
 sky130_fd_sc_hd__o22a_1 _1404_ (.A1(net195),
    .A2(net827),
    .B1(_0308_),
    .B2(net904),
    .X(net679));
 sky130_fd_sc_hd__mux2_1 _1405_ (.A0(net98),
    .A1(net31),
    .S(net895),
    .X(_0309_));
 sky130_fd_sc_hd__o22a_1 _1406_ (.A1(net165),
    .A2(net827),
    .B1(_0309_),
    .B2(net904),
    .X(net649));
 sky130_fd_sc_hd__mux2_1 _1407_ (.A0(net99),
    .A1(net32),
    .S(net896),
    .X(_0310_));
 sky130_fd_sc_hd__o22a_1 _1408_ (.A1(net166),
    .A2(net827),
    .B1(_0310_),
    .B2(net904),
    .X(net650));
 sky130_fd_sc_hd__mux2_1 _1409_ (.A0(net100),
    .A1(net33),
    .S(net895),
    .X(_0311_));
 sky130_fd_sc_hd__o22a_1 _1410_ (.A1(net167),
    .A2(net827),
    .B1(_0311_),
    .B2(net908),
    .X(net651));
 sky130_fd_sc_hd__mux2_1 _1411_ (.A0(net101),
    .A1(net34),
    .S(net898),
    .X(_0312_));
 sky130_fd_sc_hd__o22a_2 _1412_ (.A1(net168),
    .A2(net827),
    .B1(_0312_),
    .B2(net908),
    .X(net652));
 sky130_fd_sc_hd__mux2_1 _1413_ (.A0(net102),
    .A1(net35),
    .S(net899),
    .X(_0313_));
 sky130_fd_sc_hd__o22a_1 _1414_ (.A1(net169),
    .A2(net829),
    .B1(_0313_),
    .B2(net905),
    .X(net653));
 sky130_fd_sc_hd__mux2_1 _1415_ (.A0(net103),
    .A1(net36),
    .S(net899),
    .X(_0314_));
 sky130_fd_sc_hd__o22a_1 _1416_ (.A1(net170),
    .A2(net828),
    .B1(_0314_),
    .B2(net905),
    .X(net654));
 sky130_fd_sc_hd__mux2_1 _1417_ (.A0(net104),
    .A1(net37),
    .S(net899),
    .X(_0315_));
 sky130_fd_sc_hd__o22a_1 _1418_ (.A1(net171),
    .A2(net828),
    .B1(_0315_),
    .B2(net905),
    .X(net655));
 sky130_fd_sc_hd__mux2_1 _1419_ (.A0(net105),
    .A1(net38),
    .S(net898),
    .X(_0316_));
 sky130_fd_sc_hd__o22a_1 _1420_ (.A1(net172),
    .A2(net828),
    .B1(_0316_),
    .B2(net905),
    .X(net656));
 sky130_fd_sc_hd__mux2_1 _1421_ (.A0(net106),
    .A1(net39),
    .S(net898),
    .X(_0317_));
 sky130_fd_sc_hd__o22a_1 _1422_ (.A1(net173),
    .A2(net828),
    .B1(_0317_),
    .B2(net905),
    .X(net657));
 sky130_fd_sc_hd__mux2_1 _1423_ (.A0(net107),
    .A1(net40),
    .S(net900),
    .X(_0318_));
 sky130_fd_sc_hd__o22a_2 _1424_ (.A1(net174),
    .A2(net829),
    .B1(_0318_),
    .B2(net907),
    .X(net658));
 sky130_fd_sc_hd__mux2_1 _1425_ (.A0(net109),
    .A1(net42),
    .S(net898),
    .X(_0319_));
 sky130_fd_sc_hd__o22a_1 _1426_ (.A1(net176),
    .A2(net828),
    .B1(_0319_),
    .B2(net905),
    .X(net660));
 sky130_fd_sc_hd__mux2_1 _1427_ (.A0(net110),
    .A1(net43),
    .S(net899),
    .X(_0320_));
 sky130_fd_sc_hd__o22a_2 _1428_ (.A1(net177),
    .A2(net828),
    .B1(_0320_),
    .B2(net907),
    .X(net661));
 sky130_fd_sc_hd__mux2_1 _1429_ (.A0(net111),
    .A1(net44),
    .S(net899),
    .X(_0321_));
 sky130_fd_sc_hd__o22a_1 _1430_ (.A1(net178),
    .A2(net828),
    .B1(_0321_),
    .B2(net906),
    .X(net662));
 sky130_fd_sc_hd__mux2_1 _1431_ (.A0(net112),
    .A1(net45),
    .S(net899),
    .X(_0322_));
 sky130_fd_sc_hd__o22a_1 _1432_ (.A1(net179),
    .A2(net828),
    .B1(_0322_),
    .B2(net906),
    .X(net663));
 sky130_fd_sc_hd__mux2_1 _1433_ (.A0(net113),
    .A1(net46),
    .S(net900),
    .X(_0323_));
 sky130_fd_sc_hd__o22a_1 _1434_ (.A1(net180),
    .A2(net828),
    .B1(_0323_),
    .B2(net906),
    .X(net664));
 sky130_fd_sc_hd__mux2_1 _1435_ (.A0(net114),
    .A1(net47),
    .S(net900),
    .X(_0324_));
 sky130_fd_sc_hd__o22a_4 _1436_ (.A1(net181),
    .A2(net830),
    .B1(_0324_),
    .B2(net909),
    .X(net665));
 sky130_fd_sc_hd__mux2_1 _1437_ (.A0(net115),
    .A1(net48),
    .S(net900),
    .X(_0325_));
 sky130_fd_sc_hd__o22a_1 _1438_ (.A1(net182),
    .A2(net829),
    .B1(_0325_),
    .B2(net906),
    .X(net666));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(net116),
    .A1(net49),
    .S(net900),
    .X(_0326_));
 sky130_fd_sc_hd__o22a_1 _1440_ (.A1(net183),
    .A2(net828),
    .B1(_0326_),
    .B2(net906),
    .X(net667));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(net117),
    .A1(net50),
    .S(net900),
    .X(_0327_));
 sky130_fd_sc_hd__o22a_4 _1442_ (.A1(net184),
    .A2(net830),
    .B1(_0327_),
    .B2(net909),
    .X(net668));
 sky130_fd_sc_hd__mux2_1 _1443_ (.A0(net118),
    .A1(net51),
    .S(net894),
    .X(_0328_));
 sky130_fd_sc_hd__o22a_4 _1444_ (.A1(net185),
    .A2(net830),
    .B1(_0328_),
    .B2(net910),
    .X(net669));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(net120),
    .A1(net53),
    .S(net900),
    .X(_0329_));
 sky130_fd_sc_hd__o22a_2 _1446_ (.A1(net187),
    .A2(net829),
    .B1(_0329_),
    .B2(net909),
    .X(net671));
 sky130_fd_sc_hd__mux2_1 _1447_ (.A0(net121),
    .A1(net54),
    .S(net900),
    .X(_0330_));
 sky130_fd_sc_hd__o22a_4 _1448_ (.A1(net188),
    .A2(net830),
    .B1(_0330_),
    .B2(net909),
    .X(net672));
 sky130_fd_sc_hd__mux2_1 _1449_ (.A0(net62),
    .A1(net196),
    .S(net902),
    .X(_0331_));
 sky130_fd_sc_hd__a22o_4 _1450_ (.A1(net129),
    .A2(net833),
    .B1(_0331_),
    .B2(net893),
    .X(net680));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(net63),
    .A1(net197),
    .S(net902),
    .X(_0332_));
 sky130_fd_sc_hd__a22o_4 _1452_ (.A1(net130),
    .A2(net833),
    .B1(_0332_),
    .B2(net893),
    .X(net681));
 sky130_fd_sc_hd__mux2_1 _1453_ (.A0(net64),
    .A1(net198),
    .S(net902),
    .X(_0333_));
 sky130_fd_sc_hd__a22o_4 _1454_ (.A1(net131),
    .A2(net833),
    .B1(_0333_),
    .B2(net893),
    .X(net682));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(net65),
    .A1(net199),
    .S(net910),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_4 _1456_ (.A1(net132),
    .A2(net833),
    .B1(_0334_),
    .B2(net893),
    .X(net683));
 sky130_fd_sc_hd__mux2_1 _1457_ (.A0(net67),
    .A1(net201),
    .S(net910),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_4 _1458_ (.A1(net134),
    .A2(net833),
    .B1(_0335_),
    .B2(net894),
    .X(net685));
 sky130_fd_sc_hd__mux2_1 _1459_ (.A0(net66),
    .A1(net200),
    .S(net902),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_4 _1460_ (.A1(net133),
    .A2(net833),
    .B1(_0336_),
    .B2(net893),
    .X(net684));
 sky130_fd_sc_hd__o221ai_4 _1461_ (.A1(_0589_),
    .A2(_0615_),
    .B1(net980),
    .B2(_0590_),
    .C1(_0620_),
    .Y(net647));
 sky130_fd_sc_hd__nor2_1 _1462_ (.A(net889),
    .B(net881),
    .Y(_0337_));
 sky130_fd_sc_hd__mux2_1 _1463_ (.A0(net1),
    .A1(net135),
    .S(net884),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_2 _1464_ (.A1(net68),
    .A2(net823),
    .B1(_0338_),
    .B2(net876),
    .X(net686));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(net12),
    .A1(net146),
    .S(net884),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_2 _1466_ (.A1(net79),
    .A2(net823),
    .B1(_0339_),
    .B2(net876),
    .X(net697));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(net21),
    .A1(net155),
    .S(net884),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_2 _1468_ (.A1(net88),
    .A2(net823),
    .B1(_0340_),
    .B2(net876),
    .X(net702));
 sky130_fd_sc_hd__mux2_1 _1469_ (.A0(net22),
    .A1(net156),
    .S(net884),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_2 _1470_ (.A1(net89),
    .A2(net823),
    .B1(_0341_),
    .B2(net876),
    .X(net703));
 sky130_fd_sc_hd__mux2_1 _1471_ (.A0(net23),
    .A1(net157),
    .S(net885),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_2 _1472_ (.A1(net90),
    .A2(net824),
    .B1(_0342_),
    .B2(net877),
    .X(net704));
 sky130_fd_sc_hd__mux2_1 _1473_ (.A0(net24),
    .A1(net158),
    .S(net885),
    .X(_0343_));
 sky130_fd_sc_hd__a22o_1 _1474_ (.A1(net91),
    .A2(net824),
    .B1(_0343_),
    .B2(net877),
    .X(net705));
 sky130_fd_sc_hd__mux2_1 _1475_ (.A0(net25),
    .A1(net159),
    .S(net889),
    .X(_0344_));
 sky130_fd_sc_hd__a22o_4 _1476_ (.A1(net92),
    .A2(net826),
    .B1(_0344_),
    .B2(net881),
    .X(net706));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(net26),
    .A1(net160),
    .S(net887),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_4 _1478_ (.A1(net93),
    .A2(net825),
    .B1(_0345_),
    .B2(net878),
    .X(net707));
 sky130_fd_sc_hd__mux2_1 _1479_ (.A0(net27),
    .A1(net161),
    .S(net885),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_2 _1480_ (.A1(net94),
    .A2(net824),
    .B1(_0346_),
    .B2(net877),
    .X(net708));
 sky130_fd_sc_hd__mux2_1 _1481_ (.A0(net28),
    .A1(net162),
    .S(net885),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_2 _1482_ (.A1(net95),
    .A2(net824),
    .B1(_0347_),
    .B2(net877),
    .X(net709));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(net2),
    .A1(net136),
    .S(net885),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _1484_ (.A1(net69),
    .A2(net824),
    .B1(_0348_),
    .B2(net877),
    .X(net687));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(net3),
    .A1(net137),
    .S(net885),
    .X(_0349_));
 sky130_fd_sc_hd__a22o_1 _1486_ (.A1(net70),
    .A2(net824),
    .B1(_0349_),
    .B2(net877),
    .X(net688));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(net4),
    .A1(net138),
    .S(net888),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _1488_ (.A1(net71),
    .A2(net825),
    .B1(_0350_),
    .B2(net879),
    .X(net689));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(net5),
    .A1(net139),
    .S(net888),
    .X(_0351_));
 sky130_fd_sc_hd__a22o_1 _1490_ (.A1(net72),
    .A2(net825),
    .B1(_0351_),
    .B2(net879),
    .X(net690));
 sky130_fd_sc_hd__mux2_1 _1491_ (.A0(net6),
    .A1(net140),
    .S(net888),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _1492_ (.A1(net73),
    .A2(net825),
    .B1(_0352_),
    .B2(net879),
    .X(net691));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(net7),
    .A1(net141),
    .S(net887),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_2 _1494_ (.A1(net74),
    .A2(net825),
    .B1(_0353_),
    .B2(net878),
    .X(net692));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(net8),
    .A1(net142),
    .S(net887),
    .X(_0354_));
 sky130_fd_sc_hd__a22o_1 _1496_ (.A1(net75),
    .A2(net825),
    .B1(_0354_),
    .B2(net879),
    .X(net693));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(net9),
    .A1(net143),
    .S(net887),
    .X(_0355_));
 sky130_fd_sc_hd__a22o_1 _1498_ (.A1(net76),
    .A2(net825),
    .B1(_0355_),
    .B2(net878),
    .X(net694));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(net10),
    .A1(net144),
    .S(net889),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_2 _1500_ (.A1(net77),
    .A2(net825),
    .B1(_0356_),
    .B2(net881),
    .X(net695));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(net11),
    .A1(net145),
    .S(net889),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_2 _1502_ (.A1(net78),
    .A2(net825),
    .B1(_0357_),
    .B2(net881),
    .X(net696));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(net13),
    .A1(net147),
    .S(net889),
    .X(_0358_));
 sky130_fd_sc_hd__a22o_1 _1504_ (.A1(net80),
    .A2(net825),
    .B1(_0358_),
    .B2(net881),
    .X(net698));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(net14),
    .A1(net148),
    .S(net890),
    .X(_0359_));
 sky130_fd_sc_hd__a22o_1 _1506_ (.A1(net81),
    .A2(net826),
    .B1(_0359_),
    .B2(net880),
    .X(net699));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(net15),
    .A1(net149),
    .S(net890),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _1508_ (.A1(net82),
    .A2(net826),
    .B1(_0360_),
    .B2(net880),
    .X(net700));
 sky130_fd_sc_hd__mux2_1 _1509_ (.A0(net16),
    .A1(net150),
    .S(net890),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _1510_ (.A1(net83),
    .A2(net826),
    .B1(_0361_),
    .B2(net880),
    .X(net701));
 sky130_fd_sc_hd__nand2_8 _1511_ (.A(net889),
    .B(net881),
    .Y(_0362_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(net97),
    .A1(net30),
    .S(net876),
    .X(_0363_));
 sky130_fd_sc_hd__o22a_2 _1513_ (.A1(net164),
    .A2(net822),
    .B1(_0363_),
    .B2(net884),
    .X(net711));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(net108),
    .A1(net41),
    .S(net883),
    .X(_0364_));
 sky130_fd_sc_hd__o22a_2 _1515_ (.A1(net175),
    .A2(net822),
    .B1(_0364_),
    .B2(net886),
    .X(net722));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(net119),
    .A1(net52),
    .S(net883),
    .X(_0365_));
 sky130_fd_sc_hd__o22a_2 _1517_ (.A1(net186),
    .A2(net822),
    .B1(_0365_),
    .B2(net886),
    .X(net733));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(net122),
    .A1(net55),
    .S(net883),
    .X(_0366_));
 sky130_fd_sc_hd__o22a_2 _1519_ (.A1(net189),
    .A2(net822),
    .B1(_0366_),
    .B2(net886),
    .X(net736));
 sky130_fd_sc_hd__mux2_2 _1520_ (.A0(net123),
    .A1(net56),
    .S(net882),
    .X(_0367_));
 sky130_fd_sc_hd__o22a_4 _1521_ (.A1(net190),
    .A2(net820),
    .B1(_0367_),
    .B2(net889),
    .X(net737));
 sky130_fd_sc_hd__mux2_4 _1522_ (.A0(net124),
    .A1(net57),
    .S(net882),
    .X(_0368_));
 sky130_fd_sc_hd__o22a_4 _1523_ (.A1(net191),
    .A2(net820),
    .B1(_0368_),
    .B2(net889),
    .X(net738));
 sky130_fd_sc_hd__mux2_2 _1524_ (.A0(net125),
    .A1(net58),
    .S(net882),
    .X(_0369_));
 sky130_fd_sc_hd__o22a_4 _1525_ (.A1(net192),
    .A2(net820),
    .B1(_0369_),
    .B2(net891),
    .X(net739));
 sky130_fd_sc_hd__mux2_1 _1526_ (.A0(net126),
    .A1(net59),
    .S(net881),
    .X(_0370_));
 sky130_fd_sc_hd__o22a_4 _1527_ (.A1(net193),
    .A2(net820),
    .B1(_0370_),
    .B2(net891),
    .X(net740));
 sky130_fd_sc_hd__mux2_2 _1528_ (.A0(net127),
    .A1(net60),
    .S(net882),
    .X(_0371_));
 sky130_fd_sc_hd__o22a_4 _1529_ (.A1(net194),
    .A2(net821),
    .B1(_0371_),
    .B2(net887),
    .X(net741));
 sky130_fd_sc_hd__mux2_2 _1530_ (.A0(net128),
    .A1(net61),
    .S(net882),
    .X(_0372_));
 sky130_fd_sc_hd__o22a_4 _1531_ (.A1(net195),
    .A2(net821),
    .B1(_0372_),
    .B2(net889),
    .X(net742));
 sky130_fd_sc_hd__mux2_2 _1532_ (.A0(net98),
    .A1(net31),
    .S(net881),
    .X(_0373_));
 sky130_fd_sc_hd__o22a_2 _1533_ (.A1(net165),
    .A2(net822),
    .B1(_0373_),
    .B2(net887),
    .X(net712));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(net99),
    .A1(net32),
    .S(net881),
    .X(_0374_));
 sky130_fd_sc_hd__o22a_4 _1535_ (.A1(net166),
    .A2(net820),
    .B1(_0374_),
    .B2(net889),
    .X(net713));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(net100),
    .A1(net33),
    .S(net878),
    .X(_0375_));
 sky130_fd_sc_hd__o22a_1 _1537_ (.A1(net167),
    .A2(net822),
    .B1(_0375_),
    .B2(net887),
    .X(net714));
 sky130_fd_sc_hd__mux2_1 _1538_ (.A0(net101),
    .A1(net34),
    .S(net877),
    .X(_0376_));
 sky130_fd_sc_hd__o22a_2 _1539_ (.A1(net168),
    .A2(net822),
    .B1(_0376_),
    .B2(net887),
    .X(net715));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(net102),
    .A1(net35),
    .S(net878),
    .X(_0377_));
 sky130_fd_sc_hd__o22a_1 _1541_ (.A1(net169),
    .A2(net821),
    .B1(_0377_),
    .B2(net887),
    .X(net716));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(net103),
    .A1(net36),
    .S(net878),
    .X(_0378_));
 sky130_fd_sc_hd__o22a_2 _1543_ (.A1(net170),
    .A2(net821),
    .B1(_0378_),
    .B2(net887),
    .X(net717));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(net104),
    .A1(net37),
    .S(net878),
    .X(_0379_));
 sky130_fd_sc_hd__o22a_1 _1545_ (.A1(net171),
    .A2(net821),
    .B1(_0379_),
    .B2(net888),
    .X(net718));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(net105),
    .A1(net38),
    .S(net878),
    .X(_0380_));
 sky130_fd_sc_hd__o22a_1 _1547_ (.A1(net172),
    .A2(net821),
    .B1(_0380_),
    .B2(net888),
    .X(net719));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(net106),
    .A1(net39),
    .S(net878),
    .X(_0381_));
 sky130_fd_sc_hd__o22a_1 _1549_ (.A1(net173),
    .A2(net821),
    .B1(_0381_),
    .B2(net890),
    .X(net720));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(net107),
    .A1(net40),
    .S(net878),
    .X(_0382_));
 sky130_fd_sc_hd__o22a_1 _1551_ (.A1(net174),
    .A2(net821),
    .B1(_0382_),
    .B2(net890),
    .X(net721));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(net109),
    .A1(net42),
    .S(net880),
    .X(_0383_));
 sky130_fd_sc_hd__o22a_1 _1553_ (.A1(net176),
    .A2(net820),
    .B1(_0383_),
    .B2(net890),
    .X(net723));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(net110),
    .A1(net43),
    .S(net880),
    .X(_0384_));
 sky130_fd_sc_hd__o22a_1 _1555_ (.A1(net177),
    .A2(net820),
    .B1(_0384_),
    .B2(net890),
    .X(net724));
 sky130_fd_sc_hd__mux2_1 _1556_ (.A0(net111),
    .A1(net44),
    .S(net880),
    .X(_0385_));
 sky130_fd_sc_hd__o22a_1 _1557_ (.A1(net178),
    .A2(net820),
    .B1(_0385_),
    .B2(net890),
    .X(net725));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(net112),
    .A1(net45),
    .S(net880),
    .X(_0386_));
 sky130_fd_sc_hd__o22a_1 _1559_ (.A1(net179),
    .A2(net820),
    .B1(_0386_),
    .B2(net890),
    .X(net726));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(net113),
    .A1(net46),
    .S(net882),
    .X(_0387_));
 sky130_fd_sc_hd__o22a_1 _1561_ (.A1(net180),
    .A2(_0362_),
    .B1(_0387_),
    .B2(net890),
    .X(net727));
 sky130_fd_sc_hd__mux2_2 _1562_ (.A0(net114),
    .A1(net47),
    .S(net879),
    .X(_0388_));
 sky130_fd_sc_hd__o22a_1 _1563_ (.A1(net181),
    .A2(net820),
    .B1(_0388_),
    .B2(net891),
    .X(net728));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(net115),
    .A1(net48),
    .S(net880),
    .X(_0389_));
 sky130_fd_sc_hd__o22a_1 _1565_ (.A1(net182),
    .A2(_0362_),
    .B1(_0389_),
    .B2(net891),
    .X(net729));
 sky130_fd_sc_hd__mux2_1 _1566_ (.A0(net116),
    .A1(net49),
    .S(net880),
    .X(_0390_));
 sky130_fd_sc_hd__o22a_1 _1567_ (.A1(net183),
    .A2(_0362_),
    .B1(_0390_),
    .B2(net891),
    .X(net730));
 sky130_fd_sc_hd__mux2_1 _1568_ (.A0(net117),
    .A1(net50),
    .S(net879),
    .X(_0391_));
 sky130_fd_sc_hd__o22a_4 _1569_ (.A1(net184),
    .A2(net822),
    .B1(_0391_),
    .B2(net888),
    .X(net731));
 sky130_fd_sc_hd__mux2_1 _1570_ (.A0(net118),
    .A1(net51),
    .S(net877),
    .X(_0392_));
 sky130_fd_sc_hd__o22a_4 _1571_ (.A1(net185),
    .A2(net822),
    .B1(_0392_),
    .B2(net885),
    .X(net732));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(net120),
    .A1(net53),
    .S(net880),
    .X(_0393_));
 sky130_fd_sc_hd__o22a_2 _1573_ (.A1(net187),
    .A2(_0362_),
    .B1(_0393_),
    .B2(net891),
    .X(net734));
 sky130_fd_sc_hd__mux2_1 _1574_ (.A0(net121),
    .A1(net54),
    .S(net879),
    .X(_0394_));
 sky130_fd_sc_hd__o22a_4 _1575_ (.A1(net188),
    .A2(net821),
    .B1(_0394_),
    .B2(net888),
    .X(net735));
 sky130_fd_sc_hd__mux2_1 _1576_ (.A0(net62),
    .A1(net196),
    .S(net884),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_2 _1577_ (.A1(net129),
    .A2(net823),
    .B1(_0395_),
    .B2(net876),
    .X(net743));
 sky130_fd_sc_hd__mux2_1 _1578_ (.A0(net63),
    .A1(net197),
    .S(net884),
    .X(_0396_));
 sky130_fd_sc_hd__a22o_1 _1579_ (.A1(net130),
    .A2(net823),
    .B1(_0396_),
    .B2(net876),
    .X(net744));
 sky130_fd_sc_hd__mux2_1 _1580_ (.A0(net64),
    .A1(net198),
    .S(net885),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_2 _1581_ (.A1(net131),
    .A2(net823),
    .B1(_0397_),
    .B2(net876),
    .X(net745));
 sky130_fd_sc_hd__mux2_1 _1582_ (.A0(net65),
    .A1(net199),
    .S(net884),
    .X(_0398_));
 sky130_fd_sc_hd__a22o_2 _1583_ (.A1(net132),
    .A2(net823),
    .B1(_0398_),
    .B2(net876),
    .X(net746));
 sky130_fd_sc_hd__mux2_1 _1584_ (.A0(net67),
    .A1(net201),
    .S(net884),
    .X(_0399_));
 sky130_fd_sc_hd__a22o_1 _1585_ (.A1(net134),
    .A2(net823),
    .B1(_0399_),
    .B2(net877),
    .X(net748));
 sky130_fd_sc_hd__mux2_1 _1586_ (.A0(net66),
    .A1(net200),
    .S(net884),
    .X(_0400_));
 sky130_fd_sc_hd__a22o_2 _1587_ (.A1(net133),
    .A2(net823),
    .B1(_0400_),
    .B2(net876),
    .X(net747));
 sky130_fd_sc_hd__a221o_4 _1588_ (.A1(net163),
    .A2(net969),
    .B1(_0634_),
    .B2(net96),
    .C1(_0630_),
    .X(net710));
 sky130_fd_sc_hd__nand2_4 _1589_ (.A(net29),
    .B(_0036_),
    .Y(_0401_));
 sky130_fd_sc_hd__a221o_2 _1590_ (.A1(net1006),
    .A2(_0655_),
    .B1(_0036_),
    .B2(net29),
    .C1(_0594_),
    .X(_0402_));
 sky130_fd_sc_hd__a211oi_4 _1591_ (.A1(\slave4MultiMaster.arbiter.currentMaster[0] ),
    .A2(_0594_),
    .B1(net944),
    .C1(net1005),
    .Y(_0403_));
 sky130_fd_sc_hd__or4b_4 _1592_ (.A(net152),
    .B(net1014),
    .C(net1010),
    .D_N(net1012),
    .X(_0404_));
 sky130_fd_sc_hd__inv_2 _1593_ (.A(net939),
    .Y(_0405_));
 sky130_fd_sc_hd__a211o_4 _1594_ (.A1(net1006),
    .A2(_0655_),
    .B1(net939),
    .C1(_0589_),
    .X(_0406_));
 sky130_fd_sc_hd__or4_4 _1595_ (.A(_0589_),
    .B(\slave4MultiMaster.arbiter.currentMaster[0] ),
    .C(_0594_),
    .D(net939),
    .X(_0407_));
 sky130_fd_sc_hd__o211ai_4 _1596_ (.A1(_0403_),
    .A2(_0406_),
    .B1(_0407_),
    .C1(_0402_),
    .Y(_0408_));
 sky130_fd_sc_hd__and4_1 _1597_ (.A(net1006),
    .B(\slave4MultiMaster.arbiter.currentMaster[0] ),
    .C(_0594_),
    .D(_0655_),
    .X(_0409_));
 sky130_fd_sc_hd__a21o_1 _1598_ (.A1(net1006),
    .A2(_0655_),
    .B1(\slave4MultiMaster.arbiter.currentMaster[0] ),
    .X(_0410_));
 sky130_fd_sc_hd__a41oi_4 _1599_ (.A1(_0401_),
    .A2(_0406_),
    .A3(_0407_),
    .A4(_0410_),
    .B1(_0409_),
    .Y(_0411_));
 sky130_fd_sc_hd__nor2_8 _1600_ (.A(net859),
    .B(net849),
    .Y(_0412_));
 sky130_fd_sc_hd__mux2_1 _1601_ (.A0(net1),
    .A1(net135),
    .S(net859),
    .X(_0413_));
 sky130_fd_sc_hd__a22o_1 _1602_ (.A1(net68),
    .A2(net816),
    .B1(_0413_),
    .B2(net849),
    .X(net749));
 sky130_fd_sc_hd__mux2_1 _1603_ (.A0(net12),
    .A1(net146),
    .S(net857),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_2 _1604_ (.A1(net79),
    .A2(net816),
    .B1(_0414_),
    .B2(net849),
    .X(net760));
 sky130_fd_sc_hd__mux2_1 _1605_ (.A0(net21),
    .A1(net155),
    .S(net857),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_2 _1606_ (.A1(net88),
    .A2(net816),
    .B1(_0415_),
    .B2(net849),
    .X(net765));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(net22),
    .A1(net156),
    .S(net857),
    .X(_0416_));
 sky130_fd_sc_hd__a22o_2 _1608_ (.A1(net89),
    .A2(net816),
    .B1(_0416_),
    .B2(net849),
    .X(net766));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(net23),
    .A1(net157),
    .S(net857),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_2 _1610_ (.A1(net90),
    .A2(net816),
    .B1(_0417_),
    .B2(net850),
    .X(net767));
 sky130_fd_sc_hd__mux2_1 _1611_ (.A0(net24),
    .A1(net158),
    .S(net861),
    .X(_0418_));
 sky130_fd_sc_hd__a22o_1 _1612_ (.A1(net91),
    .A2(net817),
    .B1(_0418_),
    .B2(net852),
    .X(net768));
 sky130_fd_sc_hd__mux2_1 _1613_ (.A0(net25),
    .A1(net159),
    .S(net860),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_2 _1614_ (.A1(net92),
    .A2(net817),
    .B1(_0419_),
    .B2(net851),
    .X(net769));
 sky130_fd_sc_hd__mux2_1 _1615_ (.A0(net26),
    .A1(net160),
    .S(net860),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_2 _1616_ (.A1(net93),
    .A2(net818),
    .B1(_0420_),
    .B2(net851),
    .X(net770));
 sky130_fd_sc_hd__mux2_1 _1617_ (.A0(net27),
    .A1(net161),
    .S(net860),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_2 _1618_ (.A1(net94),
    .A2(net817),
    .B1(_0421_),
    .B2(net851),
    .X(net771));
 sky130_fd_sc_hd__mux2_1 _1619_ (.A0(net28),
    .A1(net162),
    .S(net860),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_2 _1620_ (.A1(net95),
    .A2(net817),
    .B1(_0422_),
    .B2(net851),
    .X(net772));
 sky130_fd_sc_hd__mux2_1 _1621_ (.A0(net2),
    .A1(net136),
    .S(net862),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_2 _1622_ (.A1(net69),
    .A2(net818),
    .B1(_0423_),
    .B2(net853),
    .X(net750));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(net3),
    .A1(net137),
    .S(net863),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_2 _1624_ (.A1(net70),
    .A2(net818),
    .B1(_0424_),
    .B2(net853),
    .X(net751));
 sky130_fd_sc_hd__mux2_1 _1625_ (.A0(net4),
    .A1(net138),
    .S(net862),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_2 _1626_ (.A1(net71),
    .A2(net818),
    .B1(_0425_),
    .B2(net853),
    .X(net752));
 sky130_fd_sc_hd__mux2_1 _1627_ (.A0(net5),
    .A1(net139),
    .S(net860),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _1628_ (.A1(net72),
    .A2(net818),
    .B1(_0426_),
    .B2(net852),
    .X(net753));
 sky130_fd_sc_hd__mux2_1 _1629_ (.A0(net6),
    .A1(net140),
    .S(net862),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _1630_ (.A1(net73),
    .A2(net818),
    .B1(_0427_),
    .B2(net853),
    .X(net754));
 sky130_fd_sc_hd__mux2_1 _1631_ (.A0(net7),
    .A1(net141),
    .S(net863),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_2 _1632_ (.A1(net74),
    .A2(net819),
    .B1(_0428_),
    .B2(net853),
    .X(net755));
 sky130_fd_sc_hd__mux2_1 _1633_ (.A0(net8),
    .A1(net142),
    .S(net862),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_2 _1634_ (.A1(net75),
    .A2(net818),
    .B1(_0429_),
    .B2(net854),
    .X(net756));
 sky130_fd_sc_hd__mux2_1 _1635_ (.A0(net9),
    .A1(net143),
    .S(net864),
    .X(_0430_));
 sky130_fd_sc_hd__a22o_4 _1636_ (.A1(net76),
    .A2(net818),
    .B1(_0430_),
    .B2(net855),
    .X(net757));
 sky130_fd_sc_hd__mux2_1 _1637_ (.A0(net10),
    .A1(net144),
    .S(net863),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_2 _1638_ (.A1(net77),
    .A2(net818),
    .B1(_0431_),
    .B2(net853),
    .X(net758));
 sky130_fd_sc_hd__mux2_1 _1639_ (.A0(net11),
    .A1(net145),
    .S(net866),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_2 _1640_ (.A1(net78),
    .A2(net818),
    .B1(_0432_),
    .B2(net855),
    .X(net759));
 sky130_fd_sc_hd__mux2_1 _1641_ (.A0(net13),
    .A1(net147),
    .S(net864),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_2 _1642_ (.A1(net80),
    .A2(net819),
    .B1(_0433_),
    .B2(net855),
    .X(net761));
 sky130_fd_sc_hd__mux2_1 _1643_ (.A0(net14),
    .A1(net148),
    .S(net864),
    .X(_0434_));
 sky130_fd_sc_hd__a22o_1 _1644_ (.A1(net81),
    .A2(net819),
    .B1(_0434_),
    .B2(net854),
    .X(net762));
 sky130_fd_sc_hd__mux2_1 _1645_ (.A0(net15),
    .A1(net149),
    .S(net864),
    .X(_0435_));
 sky130_fd_sc_hd__a22o_1 _1646_ (.A1(net82),
    .A2(net819),
    .B1(_0435_),
    .B2(net855),
    .X(net763));
 sky130_fd_sc_hd__mux2_1 _1647_ (.A0(net16),
    .A1(net150),
    .S(net864),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _1648_ (.A1(net83),
    .A2(net819),
    .B1(_0436_),
    .B2(net856),
    .X(net764));
 sky130_fd_sc_hd__nand2_8 _1649_ (.A(net858),
    .B(net850),
    .Y(_0437_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(net97),
    .A1(net30),
    .S(net850),
    .X(_0438_));
 sky130_fd_sc_hd__o22a_4 _1651_ (.A1(net164),
    .A2(net812),
    .B1(_0438_),
    .B2(net858),
    .X(net774));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(net108),
    .A1(net41),
    .S(net850),
    .X(_0439_));
 sky130_fd_sc_hd__o22a_4 _1653_ (.A1(net175),
    .A2(net812),
    .B1(_0439_),
    .B2(net858),
    .X(net785));
 sky130_fd_sc_hd__mux2_1 _1654_ (.A0(net119),
    .A1(net52),
    .S(net850),
    .X(_0440_));
 sky130_fd_sc_hd__o22a_2 _1655_ (.A1(net186),
    .A2(net812),
    .B1(_0440_),
    .B2(net857),
    .X(net796));
 sky130_fd_sc_hd__mux2_1 _1656_ (.A0(net122),
    .A1(net55),
    .S(net850),
    .X(_0441_));
 sky130_fd_sc_hd__o22a_2 _1657_ (.A1(net189),
    .A2(net812),
    .B1(_0441_),
    .B2(net857),
    .X(net799));
 sky130_fd_sc_hd__mux2_1 _1658_ (.A0(net123),
    .A1(net56),
    .S(net850),
    .X(_0442_));
 sky130_fd_sc_hd__o22a_2 _1659_ (.A1(net190),
    .A2(net812),
    .B1(_0442_),
    .B2(net857),
    .X(net800));
 sky130_fd_sc_hd__mux2_1 _1660_ (.A0(net124),
    .A1(net57),
    .S(net850),
    .X(_0443_));
 sky130_fd_sc_hd__o22a_2 _1661_ (.A1(net191),
    .A2(net812),
    .B1(_0443_),
    .B2(net858),
    .X(net801));
 sky130_fd_sc_hd__mux2_1 _1662_ (.A0(net125),
    .A1(net58),
    .S(net851),
    .X(_0444_));
 sky130_fd_sc_hd__o22a_2 _1663_ (.A1(net192),
    .A2(net812),
    .B1(_0444_),
    .B2(net860),
    .X(net802));
 sky130_fd_sc_hd__mux2_1 _1664_ (.A0(net126),
    .A1(net59),
    .S(net851),
    .X(_0445_));
 sky130_fd_sc_hd__o22a_2 _1665_ (.A1(net193),
    .A2(net812),
    .B1(_0445_),
    .B2(net860),
    .X(net803));
 sky130_fd_sc_hd__mux2_1 _1666_ (.A0(net127),
    .A1(net60),
    .S(net851),
    .X(_0446_));
 sky130_fd_sc_hd__o22a_2 _1667_ (.A1(net194),
    .A2(net812),
    .B1(_0446_),
    .B2(net860),
    .X(net804));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(net128),
    .A1(net61),
    .S(net851),
    .X(_0447_));
 sky130_fd_sc_hd__o22a_2 _1669_ (.A1(net195),
    .A2(net812),
    .B1(_0447_),
    .B2(net860),
    .X(net805));
 sky130_fd_sc_hd__mux2_1 _1670_ (.A0(net98),
    .A1(net31),
    .S(net851),
    .X(_0448_));
 sky130_fd_sc_hd__o22a_2 _1671_ (.A1(net165),
    .A2(net813),
    .B1(_0448_),
    .B2(net861),
    .X(net775));
 sky130_fd_sc_hd__mux2_1 _1672_ (.A0(net99),
    .A1(net32),
    .S(net851),
    .X(_0449_));
 sky130_fd_sc_hd__o22a_2 _1673_ (.A1(net166),
    .A2(net813),
    .B1(_0449_),
    .B2(net860),
    .X(net776));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(net100),
    .A1(net33),
    .S(net853),
    .X(_0450_));
 sky130_fd_sc_hd__o22a_2 _1675_ (.A1(net167),
    .A2(net813),
    .B1(_0450_),
    .B2(net861),
    .X(net777));
 sky130_fd_sc_hd__mux2_1 _1676_ (.A0(net101),
    .A1(net34),
    .S(net853),
    .X(_0451_));
 sky130_fd_sc_hd__o22a_2 _1677_ (.A1(net168),
    .A2(net813),
    .B1(_0451_),
    .B2(net862),
    .X(net778));
 sky130_fd_sc_hd__mux2_2 _1678_ (.A0(net102),
    .A1(net35),
    .S(net853),
    .X(_0452_));
 sky130_fd_sc_hd__o22a_1 _1679_ (.A1(net169),
    .A2(net813),
    .B1(_0452_),
    .B2(net862),
    .X(net779));
 sky130_fd_sc_hd__mux2_2 _1680_ (.A0(net103),
    .A1(net36),
    .S(net854),
    .X(_0453_));
 sky130_fd_sc_hd__o22a_2 _1681_ (.A1(net170),
    .A2(net815),
    .B1(_0453_),
    .B2(net862),
    .X(net780));
 sky130_fd_sc_hd__mux2_1 _1682_ (.A0(net104),
    .A1(net37),
    .S(net854),
    .X(_0454_));
 sky130_fd_sc_hd__o22a_2 _1683_ (.A1(net171),
    .A2(net815),
    .B1(_0454_),
    .B2(net863),
    .X(net781));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(net105),
    .A1(net38),
    .S(net853),
    .X(_0455_));
 sky130_fd_sc_hd__o22a_1 _1685_ (.A1(net172),
    .A2(net815),
    .B1(_0455_),
    .B2(net862),
    .X(net782));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(net106),
    .A1(net39),
    .S(net854),
    .X(_0456_));
 sky130_fd_sc_hd__o22a_1 _1687_ (.A1(net173),
    .A2(net815),
    .B1(_0456_),
    .B2(net862),
    .X(net783));
 sky130_fd_sc_hd__mux2_4 _1688_ (.A0(net107),
    .A1(net40),
    .S(net855),
    .X(_0457_));
 sky130_fd_sc_hd__o22a_1 _1689_ (.A1(net174),
    .A2(net815),
    .B1(_0457_),
    .B2(net862),
    .X(net784));
 sky130_fd_sc_hd__mux2_4 _1690_ (.A0(net109),
    .A1(net42),
    .S(net856),
    .X(_0458_));
 sky130_fd_sc_hd__o22a_1 _1691_ (.A1(net176),
    .A2(net815),
    .B1(_0458_),
    .B2(net864),
    .X(net786));
 sky130_fd_sc_hd__mux2_1 _1692_ (.A0(net110),
    .A1(net43),
    .S(net854),
    .X(_0459_));
 sky130_fd_sc_hd__o22a_1 _1693_ (.A1(net177),
    .A2(net814),
    .B1(_0459_),
    .B2(net864),
    .X(net787));
 sky130_fd_sc_hd__mux2_2 _1694_ (.A0(net111),
    .A1(net44),
    .S(net855),
    .X(_0460_));
 sky130_fd_sc_hd__o22a_1 _1695_ (.A1(net178),
    .A2(net814),
    .B1(_0460_),
    .B2(net864),
    .X(net788));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(net112),
    .A1(net45),
    .S(net855),
    .X(_0461_));
 sky130_fd_sc_hd__o22a_1 _1697_ (.A1(net179),
    .A2(net814),
    .B1(_0461_),
    .B2(net864),
    .X(net789));
 sky130_fd_sc_hd__mux2_1 _1698_ (.A0(net113),
    .A1(net46),
    .S(net855),
    .X(_0462_));
 sky130_fd_sc_hd__o22a_1 _1699_ (.A1(net180),
    .A2(net814),
    .B1(_0462_),
    .B2(net864),
    .X(net790));
 sky130_fd_sc_hd__mux2_1 _1700_ (.A0(net114),
    .A1(net47),
    .S(net855),
    .X(_0463_));
 sky130_fd_sc_hd__o22a_1 _1701_ (.A1(net181),
    .A2(net814),
    .B1(_0463_),
    .B2(net865),
    .X(net791));
 sky130_fd_sc_hd__mux2_1 _1702_ (.A0(net115),
    .A1(net48),
    .S(net855),
    .X(_0464_));
 sky130_fd_sc_hd__o22a_1 _1703_ (.A1(net182),
    .A2(net815),
    .B1(_0464_),
    .B2(net865),
    .X(net792));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(net116),
    .A1(net49),
    .S(net856),
    .X(_0465_));
 sky130_fd_sc_hd__o22a_1 _1705_ (.A1(net183),
    .A2(net814),
    .B1(_0465_),
    .B2(net865),
    .X(net793));
 sky130_fd_sc_hd__mux2_2 _1706_ (.A0(net117),
    .A1(net50),
    .S(net856),
    .X(_0466_));
 sky130_fd_sc_hd__o22a_1 _1707_ (.A1(net184),
    .A2(net814),
    .B1(_0466_),
    .B2(net865),
    .X(net794));
 sky130_fd_sc_hd__mux2_1 _1708_ (.A0(net118),
    .A1(net51),
    .S(net856),
    .X(_0467_));
 sky130_fd_sc_hd__o22a_1 _1709_ (.A1(net185),
    .A2(net814),
    .B1(_0467_),
    .B2(net865),
    .X(net795));
 sky130_fd_sc_hd__mux2_1 _1710_ (.A0(net120),
    .A1(net53),
    .S(net856),
    .X(_0468_));
 sky130_fd_sc_hd__o22a_1 _1711_ (.A1(net187),
    .A2(net814),
    .B1(_0468_),
    .B2(net865),
    .X(net797));
 sky130_fd_sc_hd__mux2_1 _1712_ (.A0(net121),
    .A1(net54),
    .S(net856),
    .X(_0469_));
 sky130_fd_sc_hd__o22a_1 _1713_ (.A1(net188),
    .A2(net814),
    .B1(_0469_),
    .B2(net865),
    .X(net798));
 sky130_fd_sc_hd__mux2_1 _1714_ (.A0(net62),
    .A1(net196),
    .S(net857),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_2 _1715_ (.A1(net129),
    .A2(net816),
    .B1(_0470_),
    .B2(net849),
    .X(net806));
 sky130_fd_sc_hd__mux2_1 _1716_ (.A0(net63),
    .A1(net197),
    .S(net857),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _1717_ (.A1(net130),
    .A2(net816),
    .B1(_0471_),
    .B2(net849),
    .X(net807));
 sky130_fd_sc_hd__mux2_1 _1718_ (.A0(net64),
    .A1(net198),
    .S(net859),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_2 _1719_ (.A1(net131),
    .A2(net816),
    .B1(_0472_),
    .B2(net852),
    .X(net808));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(net65),
    .A1(net199),
    .S(net858),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_2 _1721_ (.A1(net132),
    .A2(net817),
    .B1(_0473_),
    .B2(net849),
    .X(net809));
 sky130_fd_sc_hd__mux2_1 _1722_ (.A0(net67),
    .A1(net201),
    .S(net859),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _1723_ (.A1(net134),
    .A2(net816),
    .B1(_0474_),
    .B2(net849),
    .X(net811));
 sky130_fd_sc_hd__mux2_1 _1724_ (.A0(net66),
    .A1(net200),
    .S(net859),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_2 _1725_ (.A1(net133),
    .A2(net816),
    .B1(_0475_),
    .B2(net849),
    .X(net810));
 sky130_fd_sc_hd__o221ai_4 _1726_ (.A1(_0588_),
    .A2(net948),
    .B1(net939),
    .B2(_0589_),
    .C1(_0401_),
    .Y(net773));
 sky130_fd_sc_hd__a22o_1 _1727_ (.A1(net273),
    .A2(net986),
    .B1(net972),
    .B2(net308),
    .X(_0476_));
 sky130_fd_sc_hd__o22a_1 _1728_ (.A1(net1010),
    .A2(net1012),
    .B1(net343),
    .B2(net942),
    .X(_0477_));
 sky130_fd_sc_hd__a221o_1 _1729_ (.A1(net238),
    .A2(net997),
    .B1(net957),
    .B2(net203),
    .C1(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__or2_4 _1730_ (.A(_0476_),
    .B(_0478_),
    .X(net449));
 sky130_fd_sc_hd__o21a_1 _1731_ (.A1(net354),
    .A2(net940),
    .B1(net992),
    .X(_0479_));
 sky130_fd_sc_hd__a221o_1 _1732_ (.A1(net284),
    .A2(net985),
    .B1(net972),
    .B2(net319),
    .C1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__o211a_1 _1733_ (.A1(net249),
    .A2(net936),
    .B1(net938),
    .C1(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a21o_4 _1734_ (.A1(net214),
    .A2(net956),
    .B1(_0481_),
    .X(net460));
 sky130_fd_sc_hd__o21a_1 _1735_ (.A1(net365),
    .A2(net942),
    .B1(net991),
    .X(_0482_));
 sky130_fd_sc_hd__a221o_1 _1736_ (.A1(net295),
    .A2(net986),
    .B1(net970),
    .B2(net330),
    .C1(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__o211a_1 _1737_ (.A1(net260),
    .A2(net935),
    .B1(net937),
    .C1(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a21o_4 _1738_ (.A1(net225),
    .A2(net958),
    .B1(_0484_),
    .X(net471));
 sky130_fd_sc_hd__o21a_1 _1739_ (.A1(net368),
    .A2(net939),
    .B1(net990),
    .X(_0485_));
 sky130_fd_sc_hd__a221o_1 _1740_ (.A1(net298),
    .A2(net985),
    .B1(net972),
    .B2(net333),
    .C1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__o211a_1 _1741_ (.A1(net263),
    .A2(net935),
    .B1(net937),
    .C1(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a21o_4 _1742_ (.A1(net228),
    .A2(net956),
    .B1(_0487_),
    .X(net474));
 sky130_fd_sc_hd__o21a_1 _1743_ (.A1(net369),
    .A2(net942),
    .B1(net991),
    .X(_0488_));
 sky130_fd_sc_hd__a221o_1 _1744_ (.A1(net299),
    .A2(net988),
    .B1(net970),
    .B2(net334),
    .C1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__o211a_1 _1745_ (.A1(net264),
    .A2(net935),
    .B1(net937),
    .C1(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__a21o_4 _1746_ (.A1(net229),
    .A2(net958),
    .B1(_0490_),
    .X(net475));
 sky130_fd_sc_hd__a22o_1 _1747_ (.A1(net300),
    .A2(net987),
    .B1(net970),
    .B2(net335),
    .X(_0491_));
 sky130_fd_sc_hd__o22a_1 _1748_ (.A1(net1010),
    .A2(net1012),
    .B1(net370),
    .B2(net941),
    .X(_0492_));
 sky130_fd_sc_hd__a221o_1 _1749_ (.A1(net265),
    .A2(net997),
    .B1(net959),
    .B2(net230),
    .C1(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__or2_4 _1750_ (.A(_0491_),
    .B(_0493_),
    .X(net476));
 sky130_fd_sc_hd__o21a_1 _1751_ (.A1(net371),
    .A2(net941),
    .B1(net991),
    .X(_0494_));
 sky130_fd_sc_hd__a221o_2 _1752_ (.A1(net301),
    .A2(net987),
    .B1(net970),
    .B2(net336),
    .C1(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__o211a_1 _1753_ (.A1(net266),
    .A2(net936),
    .B1(net938),
    .C1(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__a21o_4 _1754_ (.A1(net231),
    .A2(net958),
    .B1(_0496_),
    .X(net477));
 sky130_fd_sc_hd__a22o_1 _1755_ (.A1(net302),
    .A2(net988),
    .B1(net971),
    .B2(net337),
    .X(_0497_));
 sky130_fd_sc_hd__o22a_1 _1756_ (.A1(net1011),
    .A2(net1013),
    .B1(net372),
    .B2(net943),
    .X(_0498_));
 sky130_fd_sc_hd__a221o_1 _1757_ (.A1(net267),
    .A2(net997),
    .B1(net959),
    .B2(net232),
    .C1(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__or2_4 _1758_ (.A(_0497_),
    .B(_0499_),
    .X(net478));
 sky130_fd_sc_hd__or2_1 _1759_ (.A(net373),
    .B(net939),
    .X(_0500_));
 sky130_fd_sc_hd__a21o_1 _1760_ (.A1(net1015),
    .A2(net338),
    .B1(net990),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_1 _1761_ (.A1(net303),
    .A2(net989),
    .B1(_0500_),
    .B2(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a21o_1 _1762_ (.A1(net1015),
    .A2(net268),
    .B1(net999),
    .X(_0503_));
 sky130_fd_sc_hd__a22o_4 _1763_ (.A1(net233),
    .A2(net956),
    .B1(_0502_),
    .B2(_0503_),
    .X(net479));
 sky130_fd_sc_hd__or2_1 _1764_ (.A(net374),
    .B(net942),
    .X(_0504_));
 sky130_fd_sc_hd__a21o_1 _1765_ (.A1(net1016),
    .A2(net339),
    .B1(net991),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _1766_ (.A1(net304),
    .A2(net986),
    .B1(_0504_),
    .B2(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__a21o_1 _1767_ (.A1(net1016),
    .A2(net269),
    .B1(net999),
    .X(_0507_));
 sky130_fd_sc_hd__a22o_4 _1768_ (.A1(net234),
    .A2(net958),
    .B1(_0506_),
    .B2(_0507_),
    .X(net480));
 sky130_fd_sc_hd__o21a_1 _1769_ (.A1(net344),
    .A2(net942),
    .B1(net991),
    .X(_0508_));
 sky130_fd_sc_hd__a221o_1 _1770_ (.A1(net274),
    .A2(net986),
    .B1(net970),
    .B2(net309),
    .C1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__o211a_1 _1771_ (.A1(net239),
    .A2(net936),
    .B1(net938),
    .C1(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__a21o_4 _1772_ (.A1(net204),
    .A2(net958),
    .B1(_0510_),
    .X(net450));
 sky130_fd_sc_hd__a22o_1 _1773_ (.A1(net275),
    .A2(net986),
    .B1(net970),
    .B2(net310),
    .X(_0511_));
 sky130_fd_sc_hd__o22a_1 _1774_ (.A1(net1011),
    .A2(net1013),
    .B1(net345),
    .B2(net942),
    .X(_0512_));
 sky130_fd_sc_hd__a221o_1 _1775_ (.A1(net240),
    .A2(net998),
    .B1(net958),
    .B2(net205),
    .C1(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__or2_4 _1776_ (.A(_0511_),
    .B(_0513_),
    .X(net451));
 sky130_fd_sc_hd__o21a_1 _1777_ (.A1(net346),
    .A2(net940),
    .B1(net990),
    .X(_0514_));
 sky130_fd_sc_hd__a221o_1 _1778_ (.A1(net276),
    .A2(net985),
    .B1(net969),
    .B2(net311),
    .C1(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__o211a_1 _1779_ (.A1(net241),
    .A2(net935),
    .B1(net937),
    .C1(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a21o_4 _1780_ (.A1(net206),
    .A2(net956),
    .B1(_0516_),
    .X(net452));
 sky130_fd_sc_hd__or2_1 _1781_ (.A(net347),
    .B(net941),
    .X(_0517_));
 sky130_fd_sc_hd__a21o_1 _1782_ (.A1(net1016),
    .A2(net312),
    .B1(net991),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _1783_ (.A1(net277),
    .A2(net987),
    .B1(_0517_),
    .B2(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__a21o_1 _1784_ (.A1(net1016),
    .A2(net242),
    .B1(_0600_),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_4 _1785_ (.A1(net207),
    .A2(net959),
    .B1(_0519_),
    .B2(_0520_),
    .X(net453));
 sky130_fd_sc_hd__a22o_1 _1786_ (.A1(net278),
    .A2(net988),
    .B1(net971),
    .B2(net313),
    .X(_0521_));
 sky130_fd_sc_hd__o22a_1 _1787_ (.A1(net1011),
    .A2(net1013),
    .B1(net348),
    .B2(net941),
    .X(_0522_));
 sky130_fd_sc_hd__a221o_1 _1788_ (.A1(net243),
    .A2(net998),
    .B1(net959),
    .B2(net208),
    .C1(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__or2_4 _1789_ (.A(_0521_),
    .B(_0523_),
    .X(net454));
 sky130_fd_sc_hd__o221a_1 _1790_ (.A1(net314),
    .A2(_0632_),
    .B1(net939),
    .B2(net349),
    .C1(_0615_),
    .X(_0524_));
 sky130_fd_sc_hd__a21o_1 _1791_ (.A1(net279),
    .A2(net985),
    .B1(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__a21o_1 _1792_ (.A1(net1014),
    .A2(net244),
    .B1(net999),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_4 _1793_ (.A1(net209),
    .A2(net957),
    .B1(_0525_),
    .B2(_0526_),
    .X(net455));
 sky130_fd_sc_hd__o21a_1 _1794_ (.A1(net350),
    .A2(net940),
    .B1(net990),
    .X(_0527_));
 sky130_fd_sc_hd__a221o_1 _1795_ (.A1(net280),
    .A2(net989),
    .B1(net969),
    .B2(net315),
    .C1(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__o211a_1 _1796_ (.A1(net245),
    .A2(net935),
    .B1(net937),
    .C1(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__a21o_4 _1797_ (.A1(net210),
    .A2(net956),
    .B1(_0529_),
    .X(net456));
 sky130_fd_sc_hd__or2_1 _1798_ (.A(net351),
    .B(net939),
    .X(_0530_));
 sky130_fd_sc_hd__a21o_1 _1799_ (.A1(net1015),
    .A2(net316),
    .B1(net990),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _1800_ (.A1(net281),
    .A2(net985),
    .B1(_0530_),
    .B2(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__a21o_1 _1801_ (.A1(net1015),
    .A2(net246),
    .B1(net999),
    .X(_0533_));
 sky130_fd_sc_hd__a22o_4 _1802_ (.A1(net211),
    .A2(net957),
    .B1(_0532_),
    .B2(_0533_),
    .X(net457));
 sky130_fd_sc_hd__o21a_1 _1803_ (.A1(net352),
    .A2(net940),
    .B1(net990),
    .X(_0534_));
 sky130_fd_sc_hd__a221o_2 _1804_ (.A1(net282),
    .A2(net989),
    .B1(net969),
    .B2(net317),
    .C1(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__o211a_1 _1805_ (.A1(net247),
    .A2(net935),
    .B1(net937),
    .C1(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__a21o_4 _1806_ (.A1(net212),
    .A2(net956),
    .B1(_0536_),
    .X(net458));
 sky130_fd_sc_hd__a22o_1 _1807_ (.A1(net283),
    .A2(net987),
    .B1(net971),
    .B2(net318),
    .X(_0537_));
 sky130_fd_sc_hd__o22a_1 _1808_ (.A1(net1011),
    .A2(net1013),
    .B1(net353),
    .B2(net943),
    .X(_0538_));
 sky130_fd_sc_hd__a221o_1 _1809_ (.A1(net248),
    .A2(net998),
    .B1(net959),
    .B2(net213),
    .C1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__or2_4 _1810_ (.A(_0537_),
    .B(_0539_),
    .X(net459));
 sky130_fd_sc_hd__a22o_1 _1811_ (.A1(net285),
    .A2(net986),
    .B1(net970),
    .B2(net320),
    .X(_0540_));
 sky130_fd_sc_hd__o22a_1 _1812_ (.A1(net1011),
    .A2(net1013),
    .B1(net355),
    .B2(net942),
    .X(_0541_));
 sky130_fd_sc_hd__a221o_1 _1813_ (.A1(net250),
    .A2(net997),
    .B1(net958),
    .B2(net215),
    .C1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__or2_4 _1814_ (.A(_0540_),
    .B(_0542_),
    .X(net461));
 sky130_fd_sc_hd__o21a_1 _1815_ (.A1(net356),
    .A2(net940),
    .B1(net990),
    .X(_0543_));
 sky130_fd_sc_hd__a221o_2 _1816_ (.A1(net286),
    .A2(net986),
    .B1(net969),
    .B2(net321),
    .C1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__o211a_1 _1817_ (.A1(net251),
    .A2(net936),
    .B1(net938),
    .C1(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__a21o_4 _1818_ (.A1(net216),
    .A2(net956),
    .B1(_0545_),
    .X(net462));
 sky130_fd_sc_hd__o21a_1 _1819_ (.A1(net357),
    .A2(net942),
    .B1(net990),
    .X(_0546_));
 sky130_fd_sc_hd__a221o_2 _1820_ (.A1(net287),
    .A2(net986),
    .B1(net969),
    .B2(net322),
    .C1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o211a_1 _1821_ (.A1(net252),
    .A2(net936),
    .B1(net938),
    .C1(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__a21o_4 _1822_ (.A1(net217),
    .A2(net956),
    .B1(_0548_),
    .X(net463));
 sky130_fd_sc_hd__o21a_1 _1823_ (.A1(net358),
    .A2(net941),
    .B1(net991),
    .X(_0549_));
 sky130_fd_sc_hd__a221o_2 _1824_ (.A1(net288),
    .A2(net987),
    .B1(net970),
    .B2(net323),
    .C1(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__a22o_1 _1825_ (.A1(net253),
    .A2(net997),
    .B1(net959),
    .B2(net218),
    .X(_0551_));
 sky130_fd_sc_hd__a21o_4 _1826_ (.A1(_0600_),
    .A2(_0550_),
    .B1(_0551_),
    .X(net464));
 sky130_fd_sc_hd__o21a_1 _1827_ (.A1(net359),
    .A2(net940),
    .B1(net990),
    .X(_0552_));
 sky130_fd_sc_hd__a221o_1 _1828_ (.A1(net289),
    .A2(net986),
    .B1(net969),
    .B2(net324),
    .C1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__o211a_1 _1829_ (.A1(net254),
    .A2(net935),
    .B1(net937),
    .C1(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__a21o_4 _1830_ (.A1(net219),
    .A2(net956),
    .B1(_0554_),
    .X(net465));
 sky130_fd_sc_hd__o21a_1 _1831_ (.A1(net360),
    .A2(net941),
    .B1(net991),
    .X(_0555_));
 sky130_fd_sc_hd__a221o_2 _1832_ (.A1(net290),
    .A2(net987),
    .B1(net970),
    .B2(net325),
    .C1(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__o211a_1 _1833_ (.A1(net255),
    .A2(net936),
    .B1(net938),
    .C1(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__a21o_4 _1834_ (.A1(net220),
    .A2(net958),
    .B1(_0557_),
    .X(net466));
 sky130_fd_sc_hd__or2_1 _1835_ (.A(net361),
    .B(net941),
    .X(_0558_));
 sky130_fd_sc_hd__a21o_1 _1836_ (.A1(net1016),
    .A2(net326),
    .B1(net991),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _1837_ (.A1(net291),
    .A2(net987),
    .B1(_0558_),
    .B2(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21o_1 _1838_ (.A1(net1016),
    .A2(net256),
    .B1(net999),
    .X(_0561_));
 sky130_fd_sc_hd__a22o_4 _1839_ (.A1(net221),
    .A2(net958),
    .B1(_0560_),
    .B2(_0561_),
    .X(net467));
 sky130_fd_sc_hd__or2_1 _1840_ (.A(net362),
    .B(net941),
    .X(_0562_));
 sky130_fd_sc_hd__a22o_1 _1841_ (.A1(net292),
    .A2(net987),
    .B1(_0562_),
    .B2(net991),
    .X(_0563_));
 sky130_fd_sc_hd__a211o_1 _1842_ (.A1(net327),
    .A2(net970),
    .B1(_0563_),
    .C1(net997),
    .X(_0564_));
 sky130_fd_sc_hd__a21o_1 _1843_ (.A1(net1016),
    .A2(net257),
    .B1(net999),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_4 _1844_ (.A1(net222),
    .A2(net959),
    .B1(_0564_),
    .B2(_0565_),
    .X(net468));
 sky130_fd_sc_hd__o221a_1 _1845_ (.A1(net328),
    .A2(_0632_),
    .B1(net939),
    .B2(net363),
    .C1(_0615_),
    .X(_0566_));
 sky130_fd_sc_hd__a21o_1 _1846_ (.A1(net293),
    .A2(net989),
    .B1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__a21o_1 _1847_ (.A1(net1015),
    .A2(net258),
    .B1(net999),
    .X(_0568_));
 sky130_fd_sc_hd__a22o_4 _1848_ (.A1(net223),
    .A2(net957),
    .B1(_0567_),
    .B2(_0568_),
    .X(net469));
 sky130_fd_sc_hd__or2_1 _1849_ (.A(net364),
    .B(net942),
    .X(_0569_));
 sky130_fd_sc_hd__a21o_1 _1850_ (.A1(net1016),
    .A2(net329),
    .B1(net992),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _1851_ (.A1(net294),
    .A2(net986),
    .B1(_0569_),
    .B2(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__a21o_1 _1852_ (.A1(net1016),
    .A2(net259),
    .B1(_0600_),
    .X(_0572_));
 sky130_fd_sc_hd__a22o_4 _1853_ (.A1(net224),
    .A2(net956),
    .B1(_0571_),
    .B2(_0572_),
    .X(net470));
 sky130_fd_sc_hd__a22o_4 _1854_ (.A1(net296),
    .A2(net987),
    .B1(net971),
    .B2(net331),
    .X(_0573_));
 sky130_fd_sc_hd__o22a_1 _1855_ (.A1(net1011),
    .A2(net1013),
    .B1(net366),
    .B2(net941),
    .X(_0574_));
 sky130_fd_sc_hd__a221o_1 _1856_ (.A1(net261),
    .A2(net997),
    .B1(net958),
    .B2(net226),
    .C1(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__or2_4 _1857_ (.A(_0573_),
    .B(_0575_),
    .X(net472));
 sky130_fd_sc_hd__or2_1 _1858_ (.A(net367),
    .B(net941),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _1859_ (.A1(net332),
    .A2(net971),
    .B1(_0576_),
    .B2(net992),
    .X(_0577_));
 sky130_fd_sc_hd__a21o_1 _1860_ (.A1(net297),
    .A2(net987),
    .B1(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__a21o_1 _1861_ (.A1(net151),
    .A2(net262),
    .B1(net999),
    .X(_0579_));
 sky130_fd_sc_hd__a22o_4 _1862_ (.A1(net227),
    .A2(net959),
    .B1(_0578_),
    .B2(_0579_),
    .X(net473));
 sky130_fd_sc_hd__a221o_1 _1863_ (.A1(net305),
    .A2(net985),
    .B1(_0405_),
    .B2(net375),
    .C1(_0601_),
    .X(_0580_));
 sky130_fd_sc_hd__a21o_1 _1864_ (.A1(net340),
    .A2(net969),
    .B1(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__o221a_4 _1865_ (.A1(net270),
    .A2(net935),
    .B1(net937),
    .B2(net235),
    .C1(_0581_),
    .X(net481));
 sky130_fd_sc_hd__a221o_1 _1866_ (.A1(net306),
    .A2(net985),
    .B1(_0405_),
    .B2(net376),
    .C1(_0601_),
    .X(_0582_));
 sky130_fd_sc_hd__a21o_1 _1867_ (.A1(net341),
    .A2(net969),
    .B1(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__o221a_4 _1868_ (.A1(net271),
    .A2(net935),
    .B1(net937),
    .B2(net236),
    .C1(_0583_),
    .X(net482));
 sky130_fd_sc_hd__mux2_1 _1869_ (.A0(net342),
    .A1(net163),
    .S(net939),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _1870_ (.A0(net307),
    .A1(_0584_),
    .S(_0632_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_2 _1871_ (.A0(net272),
    .A1(_0585_),
    .S(_0615_),
    .X(_0586_));
 sky130_fd_sc_hd__o22a_1 _1872_ (.A1(net237),
    .A2(net935),
    .B1(net937),
    .B2(net202),
    .X(_0587_));
 sky130_fd_sc_hd__o21a_4 _1873_ (.A1(_0601_),
    .A2(_0586_),
    .B1(_0587_),
    .X(net448));
 sky130_fd_sc_hd__nor2_2 _1874_ (.A(net377),
    .B(net850),
    .Y(_0000_));
 sky130_fd_sc_hd__and2b_1 _1875_ (.A_N(net377),
    .B(net857),
    .X(_0001_));
 sky130_fd_sc_hd__nor2_1 _1876_ (.A(net377),
    .B(_0652_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2b_1 _1877_ (.A_N(net377),
    .B(net490),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_1 _1878_ (.A(net377),
    .B(net934),
    .Y(_0004_));
 sky130_fd_sc_hd__and2b_1 _1879_ (.A_N(net377),
    .B(net912),
    .X(_0005_));
 sky130_fd_sc_hd__nor2_1 _1880_ (.A(net377),
    .B(_0627_),
    .Y(_0006_));
 sky130_fd_sc_hd__and2b_1 _1881_ (.A_N(net377),
    .B(net494),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_1 _1882_ (.A(net377),
    .B(_0640_),
    .Y(_0008_));
 sky130_fd_sc_hd__and2b_1 _1883_ (.A_N(net377),
    .B(net892),
    .X(_0009_));
 sky130_fd_sc_hd__dfxtp_4 _1884_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_0000_),
    .Q(\slave4MultiMaster.arbiter.currentMaster[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1885_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_0001_),
    .Q(\slave4MultiMaster.arbiter.currentMaster[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1886_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_0002_),
    .Q(\slave0MultiMaster.arbiter.currentMaster[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1887_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_0003_),
    .Q(\slave0MultiMaster.arbiter.currentMaster[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1888_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_0004_),
    .Q(\slave1MultiMaster.arbiter.currentMaster[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1889_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_0005_),
    .Q(\slave1MultiMaster.arbiter.currentMaster[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1890_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_0006_),
    .Q(\slave2MultiMaster.arbiter.currentMaster[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1891_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_0007_),
    .Q(\slave2MultiMaster.arbiter.currentMaster[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1892_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_0008_),
    .Q(\slave3MultiMaster.arbiter.currentMaster[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1893_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_0009_),
    .Q(\slave3MultiMaster.arbiter.currentMaster[1] ));
 sky130_fd_sc_hd__clkbuf_2 _1896_ (.A(net17),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_2 _1897_ (.A(net18),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_2 _1898_ (.A(net1008),
    .X(net485));
 sky130_fd_sc_hd__buf_2 _1899_ (.A(net1007),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_2 _1900_ (.A(net1015),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 _1901_ (.A(net152),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__buf_12 fanout1000 (.A(net1004),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_16 fanout1001 (.A(net1003),
    .X(net1001));
 sky130_fd_sc_hd__buf_6 fanout1002 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__buf_6 fanout1003 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_16 fanout1004 (.A(_0598_),
    .X(net1004));
 sky130_fd_sc_hd__buf_12 fanout1005 (.A(_0590_),
    .X(net1005));
 sky130_fd_sc_hd__buf_12 fanout1006 (.A(net96),
    .X(net1006));
 sky130_fd_sc_hd__buf_12 fanout1007 (.A(net85),
    .X(net1007));
 sky130_fd_sc_hd__buf_12 fanout1008 (.A(net84),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_16 fanout1009 (.A(net163),
    .X(net1009));
 sky130_fd_sc_hd__buf_12 fanout1010 (.A(net154),
    .X(net1010));
 sky130_fd_sc_hd__buf_6 fanout1011 (.A(net154),
    .X(net1011));
 sky130_fd_sc_hd__buf_12 fanout1012 (.A(net153),
    .X(net1012));
 sky130_fd_sc_hd__buf_6 fanout1013 (.A(net153),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_16 fanout1014 (.A(net1015),
    .X(net1014));
 sky130_fd_sc_hd__buf_8 fanout1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__buf_12 fanout1016 (.A(net151),
    .X(net1016));
 sky130_fd_sc_hd__buf_6 fanout812 (.A(_0437_),
    .X(net812));
 sky130_fd_sc_hd__buf_2 fanout813 (.A(_0437_),
    .X(net813));
 sky130_fd_sc_hd__buf_4 fanout814 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__buf_6 fanout815 (.A(_0437_),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_8 fanout816 (.A(net817),
    .X(net816));
 sky130_fd_sc_hd__buf_4 fanout817 (.A(_0412_),
    .X(net817));
 sky130_fd_sc_hd__buf_8 fanout818 (.A(_0412_),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 fanout819 (.A(_0412_),
    .X(net819));
 sky130_fd_sc_hd__buf_8 fanout820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__buf_12 fanout821 (.A(net822),
    .X(net821));
 sky130_fd_sc_hd__buf_12 fanout822 (.A(_0362_),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_8 fanout823 (.A(net826),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 fanout824 (.A(net826),
    .X(net824));
 sky130_fd_sc_hd__buf_6 fanout825 (.A(net826),
    .X(net825));
 sky130_fd_sc_hd__buf_8 fanout826 (.A(_0337_),
    .X(net826));
 sky130_fd_sc_hd__buf_6 fanout827 (.A(net829),
    .X(net827));
 sky130_fd_sc_hd__buf_6 fanout828 (.A(net829),
    .X(net828));
 sky130_fd_sc_hd__buf_8 fanout829 (.A(net830),
    .X(net829));
 sky130_fd_sc_hd__buf_12 fanout830 (.A(_0298_),
    .X(net830));
 sky130_fd_sc_hd__buf_6 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__buf_8 fanout832 (.A(_0273_),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_16 fanout833 (.A(_0273_),
    .X(net833));
 sky130_fd_sc_hd__buf_4 fanout834 (.A(net837),
    .X(net834));
 sky130_fd_sc_hd__buf_4 fanout835 (.A(net836),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_8 fanout836 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__buf_4 fanout837 (.A(_0234_),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_8 fanout838 (.A(net841),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_8 fanout839 (.A(net841),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 fanout840 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_8 fanout841 (.A(_0209_),
    .X(net841));
 sky130_fd_sc_hd__buf_4 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_8 fanout843 (.A(_0170_),
    .X(net843));
 sky130_fd_sc_hd__buf_6 fanout844 (.A(_0170_),
    .X(net844));
 sky130_fd_sc_hd__buf_8 fanout845 (.A(net848),
    .X(net845));
 sky130_fd_sc_hd__buf_6 fanout846 (.A(net848),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_4 fanout847 (.A(net848),
    .X(net847));
 sky130_fd_sc_hd__buf_6 fanout848 (.A(_0145_),
    .X(net848));
 sky130_fd_sc_hd__buf_8 fanout849 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__buf_12 fanout850 (.A(net852),
    .X(net850));
 sky130_fd_sc_hd__buf_8 fanout851 (.A(net852),
    .X(net851));
 sky130_fd_sc_hd__buf_6 fanout852 (.A(_0411_),
    .X(net852));
 sky130_fd_sc_hd__buf_6 fanout853 (.A(_0411_),
    .X(net853));
 sky130_fd_sc_hd__buf_4 fanout854 (.A(_0411_),
    .X(net854));
 sky130_fd_sc_hd__buf_6 fanout855 (.A(net856),
    .X(net855));
 sky130_fd_sc_hd__buf_6 fanout856 (.A(_0411_),
    .X(net856));
 sky130_fd_sc_hd__buf_6 fanout857 (.A(net859),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_8 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__buf_12 fanout859 (.A(net861),
    .X(net859));
 sky130_fd_sc_hd__buf_6 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__buf_8 fanout861 (.A(net866),
    .X(net861));
 sky130_fd_sc_hd__buf_6 fanout862 (.A(net863),
    .X(net862));
 sky130_fd_sc_hd__buf_4 fanout863 (.A(net866),
    .X(net863));
 sky130_fd_sc_hd__buf_6 fanout864 (.A(net866),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_4 fanout865 (.A(net866),
    .X(net865));
 sky130_fd_sc_hd__buf_12 fanout866 (.A(_0408_),
    .X(net866));
 sky130_fd_sc_hd__buf_6 fanout867 (.A(net868),
    .X(net867));
 sky130_fd_sc_hd__buf_4 fanout868 (.A(net490),
    .X(net868));
 sky130_fd_sc_hd__buf_6 fanout869 (.A(net875),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_4 fanout870 (.A(net875),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_8 fanout871 (.A(net875),
    .X(net871));
 sky130_fd_sc_hd__buf_6 fanout872 (.A(net874),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 fanout873 (.A(net874),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_4 fanout874 (.A(net875),
    .X(net874));
 sky130_fd_sc_hd__buf_4 fanout875 (.A(net490),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_8 fanout876 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__buf_8 fanout877 (.A(net883),
    .X(net877));
 sky130_fd_sc_hd__buf_6 fanout878 (.A(net882),
    .X(net878));
 sky130_fd_sc_hd__buf_4 fanout879 (.A(net882),
    .X(net879));
 sky130_fd_sc_hd__buf_6 fanout880 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_16 fanout881 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__buf_12 fanout882 (.A(net883),
    .X(net882));
 sky130_fd_sc_hd__buf_8 fanout883 (.A(_0640_),
    .X(net883));
 sky130_fd_sc_hd__buf_6 fanout884 (.A(net886),
    .X(net884));
 sky130_fd_sc_hd__buf_6 fanout885 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__buf_4 fanout886 (.A(net892),
    .X(net886));
 sky130_fd_sc_hd__buf_6 fanout887 (.A(net888),
    .X(net887));
 sky130_fd_sc_hd__buf_6 fanout888 (.A(net892),
    .X(net888));
 sky130_fd_sc_hd__buf_8 fanout889 (.A(net891),
    .X(net889));
 sky130_fd_sc_hd__buf_6 fanout890 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__buf_6 fanout891 (.A(net892),
    .X(net891));
 sky130_fd_sc_hd__buf_12 fanout892 (.A(net496),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_16 fanout893 (.A(net894),
    .X(net893));
 sky130_fd_sc_hd__buf_8 fanout894 (.A(net901),
    .X(net894));
 sky130_fd_sc_hd__buf_8 fanout895 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_8 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_4 fanout897 (.A(net901),
    .X(net897));
 sky130_fd_sc_hd__buf_6 fanout898 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__buf_8 fanout899 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__buf_12 fanout900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_16 fanout901 (.A(_0627_),
    .X(net901));
 sky130_fd_sc_hd__buf_8 fanout902 (.A(net910),
    .X(net902));
 sky130_fd_sc_hd__buf_6 fanout903 (.A(net908),
    .X(net903));
 sky130_fd_sc_hd__buf_8 fanout904 (.A(net908),
    .X(net904));
 sky130_fd_sc_hd__buf_6 fanout905 (.A(net907),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_4 fanout906 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__buf_6 fanout907 (.A(net908),
    .X(net907));
 sky130_fd_sc_hd__buf_6 fanout908 (.A(net909),
    .X(net908));
 sky130_fd_sc_hd__buf_12 fanout909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__buf_12 fanout910 (.A(net494),
    .X(net910));
 sky130_fd_sc_hd__buf_6 fanout911 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_6 fanout912 (.A(net492),
    .X(net912));
 sky130_fd_sc_hd__buf_6 fanout913 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__buf_6 fanout914 (.A(net492),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_8 fanout915 (.A(net918),
    .X(net915));
 sky130_fd_sc_hd__buf_4 fanout916 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_4 fanout917 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_4 fanout918 (.A(net492),
    .X(net918));
 sky130_fd_sc_hd__buf_6 fanout919 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__buf_8 fanout920 (.A(_0652_),
    .X(net920));
 sky130_fd_sc_hd__buf_6 fanout921 (.A(net926),
    .X(net921));
 sky130_fd_sc_hd__buf_4 fanout922 (.A(net926),
    .X(net922));
 sky130_fd_sc_hd__buf_6 fanout923 (.A(net926),
    .X(net923));
 sky130_fd_sc_hd__buf_6 fanout924 (.A(net925),
    .X(net924));
 sky130_fd_sc_hd__buf_8 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__buf_6 fanout926 (.A(_0652_),
    .X(net926));
 sky130_fd_sc_hd__buf_6 fanout927 (.A(net934),
    .X(net927));
 sky130_fd_sc_hd__buf_6 fanout928 (.A(net934),
    .X(net928));
 sky130_fd_sc_hd__buf_6 fanout929 (.A(net931),
    .X(net929));
 sky130_fd_sc_hd__buf_6 fanout930 (.A(net931),
    .X(net930));
 sky130_fd_sc_hd__buf_4 fanout931 (.A(net934),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_8 fanout932 (.A(net933),
    .X(net932));
 sky130_fd_sc_hd__buf_6 fanout933 (.A(net934),
    .X(net933));
 sky130_fd_sc_hd__buf_12 fanout934 (.A(_0610_),
    .X(net934));
 sky130_fd_sc_hd__buf_12 fanout935 (.A(_0603_),
    .X(net935));
 sky130_fd_sc_hd__buf_6 fanout936 (.A(_0603_),
    .X(net936));
 sky130_fd_sc_hd__buf_12 fanout937 (.A(_0645_),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_8 fanout938 (.A(_0645_),
    .X(net938));
 sky130_fd_sc_hd__buf_12 fanout939 (.A(net943),
    .X(net939));
 sky130_fd_sc_hd__buf_4 fanout940 (.A(net943),
    .X(net940));
 sky130_fd_sc_hd__buf_8 fanout941 (.A(net942),
    .X(net941));
 sky130_fd_sc_hd__buf_8 fanout942 (.A(net943),
    .X(net942));
 sky130_fd_sc_hd__buf_12 fanout943 (.A(_0404_),
    .X(net943));
 sky130_fd_sc_hd__buf_12 fanout944 (.A(net947),
    .X(net944));
 sky130_fd_sc_hd__buf_6 fanout945 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__buf_12 fanout946 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__buf_12 fanout947 (.A(_0037_),
    .X(net947));
 sky130_fd_sc_hd__buf_12 fanout948 (.A(net951),
    .X(net948));
 sky130_fd_sc_hd__buf_6 fanout949 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__buf_12 fanout950 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__buf_12 fanout951 (.A(_0656_),
    .X(net951));
 sky130_fd_sc_hd__buf_12 fanout952 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__buf_12 fanout953 (.A(_0650_),
    .X(net953));
 sky130_fd_sc_hd__buf_12 fanout954 (.A(_0650_),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_16 fanout955 (.A(_0650_),
    .X(net955));
 sky130_fd_sc_hd__buf_12 fanout956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_12 fanout957 (.A(_0644_),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_16 fanout958 (.A(net960),
    .X(net958));
 sky130_fd_sc_hd__buf_8 fanout959 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__buf_12 fanout961 (.A(_0642_),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_16 fanout962 (.A(net964),
    .X(net962));
 sky130_fd_sc_hd__buf_8 fanout963 (.A(net964),
    .X(net963));
 sky130_fd_sc_hd__buf_12 fanout964 (.A(_0642_),
    .X(net964));
 sky130_fd_sc_hd__buf_12 fanout965 (.A(_0635_),
    .X(net965));
 sky130_fd_sc_hd__buf_6 fanout966 (.A(_0635_),
    .X(net966));
 sky130_fd_sc_hd__buf_8 fanout967 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_12 fanout968 (.A(_0635_),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_16 fanout969 (.A(net972),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_16 fanout970 (.A(net972),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__buf_12 fanout972 (.A(_0631_),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_16 fanout973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_16 fanout974 (.A(_0629_),
    .X(net974));
 sky130_fd_sc_hd__buf_8 fanout975 (.A(net976),
    .X(net975));
 sky130_fd_sc_hd__buf_12 fanout976 (.A(_0629_),
    .X(net976));
 sky130_fd_sc_hd__buf_12 fanout977 (.A(net980),
    .X(net977));
 sky130_fd_sc_hd__buf_8 fanout978 (.A(net980),
    .X(net978));
 sky130_fd_sc_hd__buf_8 fanout979 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__buf_12 fanout980 (.A(_0623_),
    .X(net980));
 sky130_fd_sc_hd__buf_12 fanout981 (.A(_0619_),
    .X(net981));
 sky130_fd_sc_hd__buf_6 fanout982 (.A(_0619_),
    .X(net982));
 sky130_fd_sc_hd__buf_8 fanout983 (.A(net984),
    .X(net983));
 sky130_fd_sc_hd__buf_6 fanout984 (.A(_0619_),
    .X(net984));
 sky130_fd_sc_hd__buf_12 fanout985 (.A(net989),
    .X(net985));
 sky130_fd_sc_hd__buf_8 fanout986 (.A(net988),
    .X(net986));
 sky130_fd_sc_hd__buf_8 fanout987 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_16 fanout988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_16 fanout989 (.A(_0614_),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_16 fanout990 (.A(net992),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_16 fanout991 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__buf_12 fanout992 (.A(_0613_),
    .X(net992));
 sky130_fd_sc_hd__buf_12 fanout993 (.A(net996),
    .X(net993));
 sky130_fd_sc_hd__buf_6 fanout994 (.A(net996),
    .X(net994));
 sky130_fd_sc_hd__buf_6 fanout995 (.A(net996),
    .X(net995));
 sky130_fd_sc_hd__buf_12 fanout996 (.A(_0606_),
    .X(net996));
 sky130_fd_sc_hd__buf_12 fanout997 (.A(_0602_),
    .X(net997));
 sky130_fd_sc_hd__buf_12 fanout999 (.A(_0600_),
    .X(net999));
 sky130_fd_sc_hd__buf_12 input1 (.A(master0_wb_adr_o[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_12 input10 (.A(master0_wb_adr_o[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_12 input100 (.A(master1_wb_data_o[12]),
    .X(net100));
 sky130_fd_sc_hd__buf_12 input101 (.A(master1_wb_data_o[13]),
    .X(net101));
 sky130_fd_sc_hd__buf_12 input102 (.A(master1_wb_data_o[14]),
    .X(net102));
 sky130_fd_sc_hd__buf_12 input103 (.A(master1_wb_data_o[15]),
    .X(net103));
 sky130_fd_sc_hd__buf_12 input104 (.A(master1_wb_data_o[16]),
    .X(net104));
 sky130_fd_sc_hd__buf_12 input105 (.A(master1_wb_data_o[17]),
    .X(net105));
 sky130_fd_sc_hd__buf_12 input106 (.A(master1_wb_data_o[18]),
    .X(net106));
 sky130_fd_sc_hd__buf_12 input107 (.A(master1_wb_data_o[19]),
    .X(net107));
 sky130_fd_sc_hd__buf_12 input108 (.A(master1_wb_data_o[1]),
    .X(net108));
 sky130_fd_sc_hd__buf_12 input109 (.A(master1_wb_data_o[20]),
    .X(net109));
 sky130_fd_sc_hd__buf_12 input11 (.A(master0_wb_adr_o[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input110 (.A(master1_wb_data_o[21]),
    .X(net110));
 sky130_fd_sc_hd__buf_12 input111 (.A(master1_wb_data_o[22]),
    .X(net111));
 sky130_fd_sc_hd__buf_12 input112 (.A(master1_wb_data_o[23]),
    .X(net112));
 sky130_fd_sc_hd__buf_12 input113 (.A(master1_wb_data_o[24]),
    .X(net113));
 sky130_fd_sc_hd__buf_12 input114 (.A(master1_wb_data_o[25]),
    .X(net114));
 sky130_fd_sc_hd__buf_12 input115 (.A(master1_wb_data_o[26]),
    .X(net115));
 sky130_fd_sc_hd__buf_12 input116 (.A(master1_wb_data_o[27]),
    .X(net116));
 sky130_fd_sc_hd__buf_12 input117 (.A(master1_wb_data_o[28]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_16 input118 (.A(master1_wb_data_o[29]),
    .X(net118));
 sky130_fd_sc_hd__buf_12 input119 (.A(master1_wb_data_o[2]),
    .X(net119));
 sky130_fd_sc_hd__buf_12 input12 (.A(master0_wb_adr_o[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input120 (.A(master1_wb_data_o[30]),
    .X(net120));
 sky130_fd_sc_hd__buf_12 input121 (.A(master1_wb_data_o[31]),
    .X(net121));
 sky130_fd_sc_hd__buf_12 input122 (.A(master1_wb_data_o[3]),
    .X(net122));
 sky130_fd_sc_hd__buf_12 input123 (.A(master1_wb_data_o[4]),
    .X(net123));
 sky130_fd_sc_hd__buf_12 input124 (.A(master1_wb_data_o[5]),
    .X(net124));
 sky130_fd_sc_hd__buf_12 input125 (.A(master1_wb_data_o[6]),
    .X(net125));
 sky130_fd_sc_hd__buf_12 input126 (.A(master1_wb_data_o[7]),
    .X(net126));
 sky130_fd_sc_hd__buf_12 input127 (.A(master1_wb_data_o[8]),
    .X(net127));
 sky130_fd_sc_hd__buf_12 input128 (.A(master1_wb_data_o[9]),
    .X(net128));
 sky130_fd_sc_hd__buf_12 input129 (.A(master1_wb_sel_o[0]),
    .X(net129));
 sky130_fd_sc_hd__buf_12 input13 (.A(master0_wb_adr_o[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_12 input130 (.A(master1_wb_sel_o[1]),
    .X(net130));
 sky130_fd_sc_hd__buf_12 input131 (.A(master1_wb_sel_o[2]),
    .X(net131));
 sky130_fd_sc_hd__buf_12 input132 (.A(master1_wb_sel_o[3]),
    .X(net132));
 sky130_fd_sc_hd__buf_12 input133 (.A(master1_wb_stb_o),
    .X(net133));
 sky130_fd_sc_hd__buf_12 input134 (.A(master1_wb_we_o),
    .X(net134));
 sky130_fd_sc_hd__buf_12 input135 (.A(master2_wb_adr_o[0]),
    .X(net135));
 sky130_fd_sc_hd__buf_12 input136 (.A(master2_wb_adr_o[10]),
    .X(net136));
 sky130_fd_sc_hd__buf_12 input137 (.A(master2_wb_adr_o[11]),
    .X(net137));
 sky130_fd_sc_hd__buf_12 input138 (.A(master2_wb_adr_o[12]),
    .X(net138));
 sky130_fd_sc_hd__buf_12 input139 (.A(master2_wb_adr_o[13]),
    .X(net139));
 sky130_fd_sc_hd__buf_12 input14 (.A(master0_wb_adr_o[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input140 (.A(master2_wb_adr_o[14]),
    .X(net140));
 sky130_fd_sc_hd__buf_12 input141 (.A(master2_wb_adr_o[15]),
    .X(net141));
 sky130_fd_sc_hd__buf_12 input142 (.A(master2_wb_adr_o[16]),
    .X(net142));
 sky130_fd_sc_hd__buf_12 input143 (.A(master2_wb_adr_o[17]),
    .X(net143));
 sky130_fd_sc_hd__buf_12 input144 (.A(master2_wb_adr_o[18]),
    .X(net144));
 sky130_fd_sc_hd__buf_12 input145 (.A(master2_wb_adr_o[19]),
    .X(net145));
 sky130_fd_sc_hd__buf_12 input146 (.A(master2_wb_adr_o[1]),
    .X(net146));
 sky130_fd_sc_hd__buf_12 input147 (.A(master2_wb_adr_o[20]),
    .X(net147));
 sky130_fd_sc_hd__buf_12 input148 (.A(master2_wb_adr_o[21]),
    .X(net148));
 sky130_fd_sc_hd__buf_12 input149 (.A(master2_wb_adr_o[22]),
    .X(net149));
 sky130_fd_sc_hd__buf_12 input15 (.A(master0_wb_adr_o[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_12 input150 (.A(master2_wb_adr_o[23]),
    .X(net150));
 sky130_fd_sc_hd__buf_12 input151 (.A(master2_wb_adr_o[24]),
    .X(net151));
 sky130_fd_sc_hd__buf_8 input152 (.A(master2_wb_adr_o[25]),
    .X(net152));
 sky130_fd_sc_hd__buf_6 input153 (.A(master2_wb_adr_o[26]),
    .X(net153));
 sky130_fd_sc_hd__buf_6 input154 (.A(master2_wb_adr_o[27]),
    .X(net154));
 sky130_fd_sc_hd__buf_12 input155 (.A(master2_wb_adr_o[2]),
    .X(net155));
 sky130_fd_sc_hd__buf_12 input156 (.A(master2_wb_adr_o[3]),
    .X(net156));
 sky130_fd_sc_hd__buf_12 input157 (.A(master2_wb_adr_o[4]),
    .X(net157));
 sky130_fd_sc_hd__buf_12 input158 (.A(master2_wb_adr_o[5]),
    .X(net158));
 sky130_fd_sc_hd__buf_12 input159 (.A(master2_wb_adr_o[6]),
    .X(net159));
 sky130_fd_sc_hd__buf_12 input16 (.A(master0_wb_adr_o[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input160 (.A(master2_wb_adr_o[7]),
    .X(net160));
 sky130_fd_sc_hd__buf_12 input161 (.A(master2_wb_adr_o[8]),
    .X(net161));
 sky130_fd_sc_hd__buf_12 input162 (.A(master2_wb_adr_o[9]),
    .X(net162));
 sky130_fd_sc_hd__buf_8 input163 (.A(master2_wb_cyc_o),
    .X(net163));
 sky130_fd_sc_hd__buf_12 input164 (.A(master2_wb_data_o[0]),
    .X(net164));
 sky130_fd_sc_hd__buf_12 input165 (.A(master2_wb_data_o[10]),
    .X(net165));
 sky130_fd_sc_hd__buf_12 input166 (.A(master2_wb_data_o[11]),
    .X(net166));
 sky130_fd_sc_hd__buf_12 input167 (.A(master2_wb_data_o[12]),
    .X(net167));
 sky130_fd_sc_hd__buf_12 input168 (.A(master2_wb_data_o[13]),
    .X(net168));
 sky130_fd_sc_hd__buf_12 input169 (.A(master2_wb_data_o[14]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_16 input17 (.A(master0_wb_adr_o[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_12 input170 (.A(master2_wb_data_o[15]),
    .X(net170));
 sky130_fd_sc_hd__buf_12 input171 (.A(master2_wb_data_o[16]),
    .X(net171));
 sky130_fd_sc_hd__buf_12 input172 (.A(master2_wb_data_o[17]),
    .X(net172));
 sky130_fd_sc_hd__buf_12 input173 (.A(master2_wb_data_o[18]),
    .X(net173));
 sky130_fd_sc_hd__buf_12 input174 (.A(master2_wb_data_o[19]),
    .X(net174));
 sky130_fd_sc_hd__buf_12 input175 (.A(master2_wb_data_o[1]),
    .X(net175));
 sky130_fd_sc_hd__buf_12 input176 (.A(master2_wb_data_o[20]),
    .X(net176));
 sky130_fd_sc_hd__buf_12 input177 (.A(master2_wb_data_o[21]),
    .X(net177));
 sky130_fd_sc_hd__buf_12 input178 (.A(master2_wb_data_o[22]),
    .X(net178));
 sky130_fd_sc_hd__buf_12 input179 (.A(master2_wb_data_o[23]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_16 input18 (.A(master0_wb_adr_o[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_12 input180 (.A(master2_wb_data_o[24]),
    .X(net180));
 sky130_fd_sc_hd__buf_12 input181 (.A(master2_wb_data_o[25]),
    .X(net181));
 sky130_fd_sc_hd__buf_12 input182 (.A(master2_wb_data_o[26]),
    .X(net182));
 sky130_fd_sc_hd__buf_12 input183 (.A(master2_wb_data_o[27]),
    .X(net183));
 sky130_fd_sc_hd__buf_12 input184 (.A(master2_wb_data_o[28]),
    .X(net184));
 sky130_fd_sc_hd__buf_12 input185 (.A(master2_wb_data_o[29]),
    .X(net185));
 sky130_fd_sc_hd__buf_12 input186 (.A(master2_wb_data_o[2]),
    .X(net186));
 sky130_fd_sc_hd__buf_12 input187 (.A(master2_wb_data_o[30]),
    .X(net187));
 sky130_fd_sc_hd__buf_12 input188 (.A(master2_wb_data_o[31]),
    .X(net188));
 sky130_fd_sc_hd__buf_12 input189 (.A(master2_wb_data_o[3]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_16 input19 (.A(master0_wb_adr_o[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_12 input190 (.A(master2_wb_data_o[4]),
    .X(net190));
 sky130_fd_sc_hd__buf_12 input191 (.A(master2_wb_data_o[5]),
    .X(net191));
 sky130_fd_sc_hd__buf_12 input192 (.A(master2_wb_data_o[6]),
    .X(net192));
 sky130_fd_sc_hd__buf_12 input193 (.A(master2_wb_data_o[7]),
    .X(net193));
 sky130_fd_sc_hd__buf_12 input194 (.A(master2_wb_data_o[8]),
    .X(net194));
 sky130_fd_sc_hd__buf_12 input195 (.A(master2_wb_data_o[9]),
    .X(net195));
 sky130_fd_sc_hd__buf_12 input196 (.A(master2_wb_sel_o[0]),
    .X(net196));
 sky130_fd_sc_hd__buf_12 input197 (.A(master2_wb_sel_o[1]),
    .X(net197));
 sky130_fd_sc_hd__buf_12 input198 (.A(master2_wb_sel_o[2]),
    .X(net198));
 sky130_fd_sc_hd__buf_12 input199 (.A(master2_wb_sel_o[3]),
    .X(net199));
 sky130_fd_sc_hd__buf_12 input2 (.A(master0_wb_adr_o[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input20 (.A(master0_wb_adr_o[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_12 input200 (.A(master2_wb_stb_o),
    .X(net200));
 sky130_fd_sc_hd__buf_12 input201 (.A(master2_wb_we_o),
    .X(net201));
 sky130_fd_sc_hd__buf_12 input202 (.A(slave0_wb_ack_o),
    .X(net202));
 sky130_fd_sc_hd__buf_6 input203 (.A(slave0_wb_data_o[0]),
    .X(net203));
 sky130_fd_sc_hd__buf_6 input204 (.A(slave0_wb_data_o[10]),
    .X(net204));
 sky130_fd_sc_hd__buf_8 input205 (.A(slave0_wb_data_o[11]),
    .X(net205));
 sky130_fd_sc_hd__buf_12 input206 (.A(slave0_wb_data_o[12]),
    .X(net206));
 sky130_fd_sc_hd__buf_6 input207 (.A(slave0_wb_data_o[13]),
    .X(net207));
 sky130_fd_sc_hd__buf_4 input208 (.A(slave0_wb_data_o[14]),
    .X(net208));
 sky130_fd_sc_hd__buf_12 input209 (.A(slave0_wb_data_o[15]),
    .X(net209));
 sky130_fd_sc_hd__buf_12 input21 (.A(master0_wb_adr_o[2]),
    .X(net21));
 sky130_fd_sc_hd__buf_12 input210 (.A(slave0_wb_data_o[16]),
    .X(net210));
 sky130_fd_sc_hd__buf_12 input211 (.A(slave0_wb_data_o[17]),
    .X(net211));
 sky130_fd_sc_hd__buf_12 input212 (.A(slave0_wb_data_o[18]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_8 input213 (.A(slave0_wb_data_o[19]),
    .X(net213));
 sky130_fd_sc_hd__buf_8 input214 (.A(slave0_wb_data_o[1]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_16 input215 (.A(slave0_wb_data_o[20]),
    .X(net215));
 sky130_fd_sc_hd__buf_12 input216 (.A(slave0_wb_data_o[21]),
    .X(net216));
 sky130_fd_sc_hd__buf_12 input217 (.A(slave0_wb_data_o[22]),
    .X(net217));
 sky130_fd_sc_hd__buf_6 input218 (.A(slave0_wb_data_o[23]),
    .X(net218));
 sky130_fd_sc_hd__buf_12 input219 (.A(slave0_wb_data_o[24]),
    .X(net219));
 sky130_fd_sc_hd__buf_12 input22 (.A(master0_wb_adr_o[3]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 input220 (.A(slave0_wb_data_o[25]),
    .X(net220));
 sky130_fd_sc_hd__buf_8 input221 (.A(slave0_wb_data_o[26]),
    .X(net221));
 sky130_fd_sc_hd__buf_6 input222 (.A(slave0_wb_data_o[27]),
    .X(net222));
 sky130_fd_sc_hd__buf_12 input223 (.A(slave0_wb_data_o[28]),
    .X(net223));
 sky130_fd_sc_hd__buf_12 input224 (.A(slave0_wb_data_o[29]),
    .X(net224));
 sky130_fd_sc_hd__buf_6 input225 (.A(slave0_wb_data_o[2]),
    .X(net225));
 sky130_fd_sc_hd__buf_8 input226 (.A(slave0_wb_data_o[30]),
    .X(net226));
 sky130_fd_sc_hd__buf_6 input227 (.A(slave0_wb_data_o[31]),
    .X(net227));
 sky130_fd_sc_hd__buf_8 input228 (.A(slave0_wb_data_o[3]),
    .X(net228));
 sky130_fd_sc_hd__buf_6 input229 (.A(slave0_wb_data_o[4]),
    .X(net229));
 sky130_fd_sc_hd__buf_12 input23 (.A(master0_wb_adr_o[4]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input230 (.A(slave0_wb_data_o[5]),
    .X(net230));
 sky130_fd_sc_hd__buf_6 input231 (.A(slave0_wb_data_o[6]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 input232 (.A(slave0_wb_data_o[7]),
    .X(net232));
 sky130_fd_sc_hd__buf_12 input233 (.A(slave0_wb_data_o[8]),
    .X(net233));
 sky130_fd_sc_hd__buf_8 input234 (.A(slave0_wb_data_o[9]),
    .X(net234));
 sky130_fd_sc_hd__buf_12 input235 (.A(slave0_wb_error_o),
    .X(net235));
 sky130_fd_sc_hd__buf_12 input236 (.A(slave0_wb_stall_o),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 input237 (.A(slave1_wb_ack_o),
    .X(net237));
 sky130_fd_sc_hd__buf_4 input238 (.A(slave1_wb_data_o[0]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_8 input239 (.A(slave1_wb_data_o[10]),
    .X(net239));
 sky130_fd_sc_hd__buf_12 input24 (.A(master0_wb_adr_o[5]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input240 (.A(slave1_wb_data_o[11]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 input241 (.A(slave1_wb_data_o[12]),
    .X(net241));
 sky130_fd_sc_hd__buf_6 input242 (.A(slave1_wb_data_o[13]),
    .X(net242));
 sky130_fd_sc_hd__buf_8 input243 (.A(slave1_wb_data_o[14]),
    .X(net243));
 sky130_fd_sc_hd__buf_4 input244 (.A(slave1_wb_data_o[15]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 input245 (.A(slave1_wb_data_o[16]),
    .X(net245));
 sky130_fd_sc_hd__buf_4 input246 (.A(slave1_wb_data_o[17]),
    .X(net246));
 sky130_fd_sc_hd__buf_4 input247 (.A(slave1_wb_data_o[18]),
    .X(net247));
 sky130_fd_sc_hd__buf_8 input248 (.A(slave1_wb_data_o[19]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 input249 (.A(slave1_wb_data_o[1]),
    .X(net249));
 sky130_fd_sc_hd__buf_12 input25 (.A(master0_wb_adr_o[6]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input250 (.A(slave1_wb_data_o[20]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 input251 (.A(slave1_wb_data_o[21]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_4 input252 (.A(slave1_wb_data_o[22]),
    .X(net252));
 sky130_fd_sc_hd__buf_6 input253 (.A(slave1_wb_data_o[23]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 input254 (.A(slave1_wb_data_o[24]),
    .X(net254));
 sky130_fd_sc_hd__buf_6 input255 (.A(slave1_wb_data_o[25]),
    .X(net255));
 sky130_fd_sc_hd__buf_6 input256 (.A(slave1_wb_data_o[26]),
    .X(net256));
 sky130_fd_sc_hd__buf_6 input257 (.A(slave1_wb_data_o[27]),
    .X(net257));
 sky130_fd_sc_hd__buf_4 input258 (.A(slave1_wb_data_o[28]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 input259 (.A(slave1_wb_data_o[29]),
    .X(net259));
 sky130_fd_sc_hd__buf_12 input26 (.A(master0_wb_adr_o[7]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input260 (.A(slave1_wb_data_o[2]),
    .X(net260));
 sky130_fd_sc_hd__buf_6 input261 (.A(slave1_wb_data_o[30]),
    .X(net261));
 sky130_fd_sc_hd__buf_6 input262 (.A(slave1_wb_data_o[31]),
    .X(net262));
 sky130_fd_sc_hd__buf_2 input263 (.A(slave1_wb_data_o[3]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_8 input264 (.A(slave1_wb_data_o[4]),
    .X(net264));
 sky130_fd_sc_hd__buf_6 input265 (.A(slave1_wb_data_o[5]),
    .X(net265));
 sky130_fd_sc_hd__buf_6 input266 (.A(slave1_wb_data_o[6]),
    .X(net266));
 sky130_fd_sc_hd__buf_8 input267 (.A(slave1_wb_data_o[7]),
    .X(net267));
 sky130_fd_sc_hd__buf_2 input268 (.A(slave1_wb_data_o[8]),
    .X(net268));
 sky130_fd_sc_hd__buf_4 input269 (.A(slave1_wb_data_o[9]),
    .X(net269));
 sky130_fd_sc_hd__buf_12 input27 (.A(master0_wb_adr_o[8]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input270 (.A(slave1_wb_error_o),
    .X(net270));
 sky130_fd_sc_hd__buf_4 input271 (.A(slave1_wb_stall_o),
    .X(net271));
 sky130_fd_sc_hd__buf_12 input272 (.A(slave2_wb_ack_o),
    .X(net272));
 sky130_fd_sc_hd__buf_8 input273 (.A(slave2_wb_data_o[0]),
    .X(net273));
 sky130_fd_sc_hd__buf_6 input274 (.A(slave2_wb_data_o[10]),
    .X(net274));
 sky130_fd_sc_hd__buf_6 input275 (.A(slave2_wb_data_o[11]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_16 input276 (.A(slave2_wb_data_o[12]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_8 input277 (.A(slave2_wb_data_o[13]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 input278 (.A(slave2_wb_data_o[14]),
    .X(net278));
 sky130_fd_sc_hd__buf_12 input279 (.A(slave2_wb_data_o[15]),
    .X(net279));
 sky130_fd_sc_hd__buf_12 input28 (.A(master0_wb_adr_o[9]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_16 input280 (.A(slave2_wb_data_o[16]),
    .X(net280));
 sky130_fd_sc_hd__buf_12 input281 (.A(slave2_wb_data_o[17]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_16 input282 (.A(slave2_wb_data_o[18]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 input283 (.A(slave2_wb_data_o[19]),
    .X(net283));
 sky130_fd_sc_hd__buf_8 input284 (.A(slave2_wb_data_o[1]),
    .X(net284));
 sky130_fd_sc_hd__buf_8 input285 (.A(slave2_wb_data_o[20]),
    .X(net285));
 sky130_fd_sc_hd__buf_8 input286 (.A(slave2_wb_data_o[21]),
    .X(net286));
 sky130_fd_sc_hd__buf_8 input287 (.A(slave2_wb_data_o[22]),
    .X(net287));
 sky130_fd_sc_hd__buf_6 input288 (.A(slave2_wb_data_o[23]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_16 input289 (.A(slave2_wb_data_o[24]),
    .X(net289));
 sky130_fd_sc_hd__buf_6 input29 (.A(master0_wb_cyc_o),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input290 (.A(slave2_wb_data_o[25]),
    .X(net290));
 sky130_fd_sc_hd__buf_6 input291 (.A(slave2_wb_data_o[26]),
    .X(net291));
 sky130_fd_sc_hd__buf_6 input292 (.A(slave2_wb_data_o[27]),
    .X(net292));
 sky130_fd_sc_hd__buf_12 input293 (.A(slave2_wb_data_o[28]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_16 input294 (.A(slave2_wb_data_o[29]),
    .X(net294));
 sky130_fd_sc_hd__buf_6 input295 (.A(slave2_wb_data_o[2]),
    .X(net295));
 sky130_fd_sc_hd__buf_6 input296 (.A(slave2_wb_data_o[30]),
    .X(net296));
 sky130_fd_sc_hd__buf_6 input297 (.A(slave2_wb_data_o[31]),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_16 input298 (.A(slave2_wb_data_o[3]),
    .X(net298));
 sky130_fd_sc_hd__buf_6 input299 (.A(slave2_wb_data_o[4]),
    .X(net299));
 sky130_fd_sc_hd__buf_12 input3 (.A(master0_wb_adr_o[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_12 input30 (.A(master0_wb_data_o[0]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input300 (.A(slave2_wb_data_o[5]),
    .X(net300));
 sky130_fd_sc_hd__buf_4 input301 (.A(slave2_wb_data_o[6]),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 input302 (.A(slave2_wb_data_o[7]),
    .X(net302));
 sky130_fd_sc_hd__buf_8 input303 (.A(slave2_wb_data_o[8]),
    .X(net303));
 sky130_fd_sc_hd__buf_6 input304 (.A(slave2_wb_data_o[9]),
    .X(net304));
 sky130_fd_sc_hd__buf_12 input305 (.A(slave2_wb_error_o),
    .X(net305));
 sky130_fd_sc_hd__buf_12 input306 (.A(slave2_wb_stall_o),
    .X(net306));
 sky130_fd_sc_hd__buf_8 input307 (.A(slave3_wb_ack_o),
    .X(net307));
 sky130_fd_sc_hd__buf_4 input308 (.A(slave3_wb_data_o[0]),
    .X(net308));
 sky130_fd_sc_hd__buf_4 input309 (.A(slave3_wb_data_o[10]),
    .X(net309));
 sky130_fd_sc_hd__buf_12 input31 (.A(master0_wb_data_o[10]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 input310 (.A(slave3_wb_data_o[11]),
    .X(net310));
 sky130_fd_sc_hd__buf_8 input311 (.A(slave3_wb_data_o[12]),
    .X(net311));
 sky130_fd_sc_hd__buf_4 input312 (.A(slave3_wb_data_o[13]),
    .X(net312));
 sky130_fd_sc_hd__buf_4 input313 (.A(slave3_wb_data_o[14]),
    .X(net313));
 sky130_fd_sc_hd__buf_12 input314 (.A(slave3_wb_data_o[15]),
    .X(net314));
 sky130_fd_sc_hd__buf_8 input315 (.A(slave3_wb_data_o[16]),
    .X(net315));
 sky130_fd_sc_hd__buf_12 input316 (.A(slave3_wb_data_o[17]),
    .X(net316));
 sky130_fd_sc_hd__buf_8 input317 (.A(slave3_wb_data_o[18]),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 input318 (.A(slave3_wb_data_o[19]),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_8 input319 (.A(slave3_wb_data_o[1]),
    .X(net319));
 sky130_fd_sc_hd__buf_12 input32 (.A(master0_wb_data_o[11]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input320 (.A(slave3_wb_data_o[20]),
    .X(net320));
 sky130_fd_sc_hd__buf_8 input321 (.A(slave3_wb_data_o[21]),
    .X(net321));
 sky130_fd_sc_hd__buf_8 input322 (.A(slave3_wb_data_o[22]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_8 input323 (.A(slave3_wb_data_o[23]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_16 input324 (.A(slave3_wb_data_o[24]),
    .X(net324));
 sky130_fd_sc_hd__buf_6 input325 (.A(slave3_wb_data_o[25]),
    .X(net325));
 sky130_fd_sc_hd__buf_6 input326 (.A(slave3_wb_data_o[26]),
    .X(net326));
 sky130_fd_sc_hd__buf_6 input327 (.A(slave3_wb_data_o[27]),
    .X(net327));
 sky130_fd_sc_hd__buf_12 input328 (.A(slave3_wb_data_o[28]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_16 input329 (.A(slave3_wb_data_o[29]),
    .X(net329));
 sky130_fd_sc_hd__buf_12 input33 (.A(master0_wb_data_o[12]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input330 (.A(slave3_wb_data_o[2]),
    .X(net330));
 sky130_fd_sc_hd__buf_6 input331 (.A(slave3_wb_data_o[30]),
    .X(net331));
 sky130_fd_sc_hd__buf_6 input332 (.A(slave3_wb_data_o[31]),
    .X(net332));
 sky130_fd_sc_hd__buf_6 input333 (.A(slave3_wb_data_o[3]),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 input334 (.A(slave3_wb_data_o[4]),
    .X(net334));
 sky130_fd_sc_hd__buf_4 input335 (.A(slave3_wb_data_o[5]),
    .X(net335));
 sky130_fd_sc_hd__buf_4 input336 (.A(slave3_wb_data_o[6]),
    .X(net336));
 sky130_fd_sc_hd__buf_6 input337 (.A(slave3_wb_data_o[7]),
    .X(net337));
 sky130_fd_sc_hd__buf_6 input338 (.A(slave3_wb_data_o[8]),
    .X(net338));
 sky130_fd_sc_hd__buf_6 input339 (.A(slave3_wb_data_o[9]),
    .X(net339));
 sky130_fd_sc_hd__buf_12 input34 (.A(master0_wb_data_o[13]),
    .X(net34));
 sky130_fd_sc_hd__buf_8 input340 (.A(slave3_wb_error_o),
    .X(net340));
 sky130_fd_sc_hd__buf_8 input341 (.A(slave3_wb_stall_o),
    .X(net341));
 sky130_fd_sc_hd__buf_6 input342 (.A(slave4_wb_ack_o),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_16 input343 (.A(slave4_wb_data_o[0]),
    .X(net343));
 sky130_fd_sc_hd__buf_8 input344 (.A(slave4_wb_data_o[10]),
    .X(net344));
 sky130_fd_sc_hd__buf_6 input345 (.A(slave4_wb_data_o[11]),
    .X(net345));
 sky130_fd_sc_hd__buf_4 input346 (.A(slave4_wb_data_o[12]),
    .X(net346));
 sky130_fd_sc_hd__buf_8 input347 (.A(slave4_wb_data_o[13]),
    .X(net347));
 sky130_fd_sc_hd__buf_12 input348 (.A(slave4_wb_data_o[14]),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_4 input349 (.A(slave4_wb_data_o[15]),
    .X(net349));
 sky130_fd_sc_hd__buf_12 input35 (.A(master0_wb_data_o[14]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input350 (.A(slave4_wb_data_o[16]),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_4 input351 (.A(slave4_wb_data_o[17]),
    .X(net351));
 sky130_fd_sc_hd__buf_2 input352 (.A(slave4_wb_data_o[18]),
    .X(net352));
 sky130_fd_sc_hd__buf_8 input353 (.A(slave4_wb_data_o[19]),
    .X(net353));
 sky130_fd_sc_hd__buf_8 input354 (.A(slave4_wb_data_o[1]),
    .X(net354));
 sky130_fd_sc_hd__buf_4 input355 (.A(slave4_wb_data_o[20]),
    .X(net355));
 sky130_fd_sc_hd__buf_2 input356 (.A(slave4_wb_data_o[21]),
    .X(net356));
 sky130_fd_sc_hd__buf_4 input357 (.A(slave4_wb_data_o[22]),
    .X(net357));
 sky130_fd_sc_hd__buf_6 input358 (.A(slave4_wb_data_o[23]),
    .X(net358));
 sky130_fd_sc_hd__buf_2 input359 (.A(slave4_wb_data_o[24]),
    .X(net359));
 sky130_fd_sc_hd__buf_12 input36 (.A(master0_wb_data_o[15]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input360 (.A(slave4_wb_data_o[25]),
    .X(net360));
 sky130_fd_sc_hd__buf_6 input361 (.A(slave4_wb_data_o[26]),
    .X(net361));
 sky130_fd_sc_hd__buf_6 input362 (.A(slave4_wb_data_o[27]),
    .X(net362));
 sky130_fd_sc_hd__buf_6 input363 (.A(slave4_wb_data_o[28]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 input364 (.A(slave4_wb_data_o[29]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_16 input365 (.A(slave4_wb_data_o[2]),
    .X(net365));
 sky130_fd_sc_hd__buf_6 input366 (.A(slave4_wb_data_o[30]),
    .X(net366));
 sky130_fd_sc_hd__buf_4 input367 (.A(slave4_wb_data_o[31]),
    .X(net367));
 sky130_fd_sc_hd__buf_6 input368 (.A(slave4_wb_data_o[3]),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_16 input369 (.A(slave4_wb_data_o[4]),
    .X(net369));
 sky130_fd_sc_hd__buf_12 input37 (.A(master0_wb_data_o[16]),
    .X(net37));
 sky130_fd_sc_hd__buf_12 input370 (.A(slave4_wb_data_o[5]),
    .X(net370));
 sky130_fd_sc_hd__buf_12 input371 (.A(slave4_wb_data_o[6]),
    .X(net371));
 sky130_fd_sc_hd__buf_12 input372 (.A(slave4_wb_data_o[7]),
    .X(net372));
 sky130_fd_sc_hd__buf_6 input373 (.A(slave4_wb_data_o[8]),
    .X(net373));
 sky130_fd_sc_hd__buf_6 input374 (.A(slave4_wb_data_o[9]),
    .X(net374));
 sky130_fd_sc_hd__buf_6 input375 (.A(slave4_wb_error_o),
    .X(net375));
 sky130_fd_sc_hd__buf_6 input376 (.A(slave4_wb_stall_o),
    .X(net376));
 sky130_fd_sc_hd__buf_6 input377 (.A(wb_rst_i),
    .X(net377));
 sky130_fd_sc_hd__buf_12 input38 (.A(master0_wb_data_o[17]),
    .X(net38));
 sky130_fd_sc_hd__buf_12 input39 (.A(master0_wb_data_o[18]),
    .X(net39));
 sky130_fd_sc_hd__buf_12 input4 (.A(master0_wb_adr_o[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input40 (.A(master0_wb_data_o[19]),
    .X(net40));
 sky130_fd_sc_hd__buf_12 input41 (.A(master0_wb_data_o[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_12 input42 (.A(master0_wb_data_o[20]),
    .X(net42));
 sky130_fd_sc_hd__buf_12 input43 (.A(master0_wb_data_o[21]),
    .X(net43));
 sky130_fd_sc_hd__buf_12 input44 (.A(master0_wb_data_o[22]),
    .X(net44));
 sky130_fd_sc_hd__buf_12 input45 (.A(master0_wb_data_o[23]),
    .X(net45));
 sky130_fd_sc_hd__buf_12 input46 (.A(master0_wb_data_o[24]),
    .X(net46));
 sky130_fd_sc_hd__buf_12 input47 (.A(master0_wb_data_o[25]),
    .X(net47));
 sky130_fd_sc_hd__buf_12 input48 (.A(master0_wb_data_o[26]),
    .X(net48));
 sky130_fd_sc_hd__buf_12 input49 (.A(master0_wb_data_o[27]),
    .X(net49));
 sky130_fd_sc_hd__buf_12 input5 (.A(master0_wb_adr_o[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input50 (.A(master0_wb_data_o[28]),
    .X(net50));
 sky130_fd_sc_hd__buf_12 input51 (.A(master0_wb_data_o[29]),
    .X(net51));
 sky130_fd_sc_hd__buf_12 input52 (.A(master0_wb_data_o[2]),
    .X(net52));
 sky130_fd_sc_hd__buf_12 input53 (.A(master0_wb_data_o[30]),
    .X(net53));
 sky130_fd_sc_hd__buf_12 input54 (.A(master0_wb_data_o[31]),
    .X(net54));
 sky130_fd_sc_hd__buf_12 input55 (.A(master0_wb_data_o[3]),
    .X(net55));
 sky130_fd_sc_hd__buf_12 input56 (.A(master0_wb_data_o[4]),
    .X(net56));
 sky130_fd_sc_hd__buf_12 input57 (.A(master0_wb_data_o[5]),
    .X(net57));
 sky130_fd_sc_hd__buf_12 input58 (.A(master0_wb_data_o[6]),
    .X(net58));
 sky130_fd_sc_hd__buf_12 input59 (.A(master0_wb_data_o[7]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input6 (.A(master0_wb_adr_o[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input60 (.A(master0_wb_data_o[8]),
    .X(net60));
 sky130_fd_sc_hd__buf_12 input61 (.A(master0_wb_data_o[9]),
    .X(net61));
 sky130_fd_sc_hd__buf_12 input62 (.A(master0_wb_sel_o[0]),
    .X(net62));
 sky130_fd_sc_hd__buf_12 input63 (.A(master0_wb_sel_o[1]),
    .X(net63));
 sky130_fd_sc_hd__buf_12 input64 (.A(master0_wb_sel_o[2]),
    .X(net64));
 sky130_fd_sc_hd__buf_12 input65 (.A(master0_wb_sel_o[3]),
    .X(net65));
 sky130_fd_sc_hd__buf_12 input66 (.A(master0_wb_stb_o),
    .X(net66));
 sky130_fd_sc_hd__buf_12 input67 (.A(master0_wb_we_o),
    .X(net67));
 sky130_fd_sc_hd__buf_12 input68 (.A(master1_wb_adr_o[0]),
    .X(net68));
 sky130_fd_sc_hd__buf_12 input69 (.A(master1_wb_adr_o[10]),
    .X(net69));
 sky130_fd_sc_hd__buf_12 input7 (.A(master0_wb_adr_o[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_12 input70 (.A(master1_wb_adr_o[11]),
    .X(net70));
 sky130_fd_sc_hd__buf_12 input71 (.A(master1_wb_adr_o[12]),
    .X(net71));
 sky130_fd_sc_hd__buf_12 input72 (.A(master1_wb_adr_o[13]),
    .X(net72));
 sky130_fd_sc_hd__buf_12 input73 (.A(master1_wb_adr_o[14]),
    .X(net73));
 sky130_fd_sc_hd__buf_12 input74 (.A(master1_wb_adr_o[15]),
    .X(net74));
 sky130_fd_sc_hd__buf_12 input75 (.A(master1_wb_adr_o[16]),
    .X(net75));
 sky130_fd_sc_hd__buf_12 input76 (.A(master1_wb_adr_o[17]),
    .X(net76));
 sky130_fd_sc_hd__buf_12 input77 (.A(master1_wb_adr_o[18]),
    .X(net77));
 sky130_fd_sc_hd__buf_12 input78 (.A(master1_wb_adr_o[19]),
    .X(net78));
 sky130_fd_sc_hd__buf_12 input79 (.A(master1_wb_adr_o[1]),
    .X(net79));
 sky130_fd_sc_hd__buf_12 input8 (.A(master0_wb_adr_o[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input80 (.A(master1_wb_adr_o[20]),
    .X(net80));
 sky130_fd_sc_hd__buf_12 input81 (.A(master1_wb_adr_o[21]),
    .X(net81));
 sky130_fd_sc_hd__buf_12 input82 (.A(master1_wb_adr_o[22]),
    .X(net82));
 sky130_fd_sc_hd__buf_12 input83 (.A(master1_wb_adr_o[23]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(master1_wb_adr_o[24]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(master1_wb_adr_o[25]),
    .X(net85));
 sky130_fd_sc_hd__buf_12 input86 (.A(master1_wb_adr_o[26]),
    .X(net86));
 sky130_fd_sc_hd__buf_12 input87 (.A(master1_wb_adr_o[27]),
    .X(net87));
 sky130_fd_sc_hd__buf_12 input88 (.A(master1_wb_adr_o[2]),
    .X(net88));
 sky130_fd_sc_hd__buf_12 input89 (.A(master1_wb_adr_o[3]),
    .X(net89));
 sky130_fd_sc_hd__buf_12 input9 (.A(master0_wb_adr_o[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input90 (.A(master1_wb_adr_o[4]),
    .X(net90));
 sky130_fd_sc_hd__buf_12 input91 (.A(master1_wb_adr_o[5]),
    .X(net91));
 sky130_fd_sc_hd__buf_12 input92 (.A(master1_wb_adr_o[6]),
    .X(net92));
 sky130_fd_sc_hd__buf_12 input93 (.A(master1_wb_adr_o[7]),
    .X(net93));
 sky130_fd_sc_hd__buf_12 input94 (.A(master1_wb_adr_o[8]),
    .X(net94));
 sky130_fd_sc_hd__buf_12 input95 (.A(master1_wb_adr_o[9]),
    .X(net95));
 sky130_fd_sc_hd__buf_8 input96 (.A(master1_wb_cyc_o),
    .X(net96));
 sky130_fd_sc_hd__buf_12 input97 (.A(master1_wb_data_o[0]),
    .X(net97));
 sky130_fd_sc_hd__buf_12 input98 (.A(master1_wb_data_o[10]),
    .X(net98));
 sky130_fd_sc_hd__buf_12 input99 (.A(master1_wb_data_o[11]),
    .X(net99));
 sky130_fd_sc_hd__buf_4 output378 (.A(net378),
    .X(master0_wb_ack_i));
 sky130_fd_sc_hd__buf_4 output379 (.A(net379),
    .X(master0_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output380 (.A(net380),
    .X(master0_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output381 (.A(net381),
    .X(master0_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output382 (.A(net382),
    .X(master0_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output383 (.A(net383),
    .X(master0_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output384 (.A(net384),
    .X(master0_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output385 (.A(net385),
    .X(master0_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output386 (.A(net386),
    .X(master0_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output387 (.A(net387),
    .X(master0_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output388 (.A(net388),
    .X(master0_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output389 (.A(net389),
    .X(master0_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output390 (.A(net390),
    .X(master0_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output391 (.A(net391),
    .X(master0_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output392 (.A(net392),
    .X(master0_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output393 (.A(net393),
    .X(master0_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output394 (.A(net394),
    .X(master0_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output395 (.A(net395),
    .X(master0_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output396 (.A(net396),
    .X(master0_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output397 (.A(net397),
    .X(master0_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output398 (.A(net398),
    .X(master0_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output399 (.A(net399),
    .X(master0_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output400 (.A(net400),
    .X(master0_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output401 (.A(net401),
    .X(master0_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output402 (.A(net402),
    .X(master0_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output403 (.A(net403),
    .X(master0_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output404 (.A(net404),
    .X(master0_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output405 (.A(net405),
    .X(master0_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output406 (.A(net406),
    .X(master0_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output407 (.A(net407),
    .X(master0_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output408 (.A(net408),
    .X(master0_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output409 (.A(net409),
    .X(master0_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output410 (.A(net410),
    .X(master0_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output411 (.A(net411),
    .X(master0_wb_error_i));
 sky130_fd_sc_hd__buf_4 output412 (.A(net412),
    .X(master0_wb_stall_i));
 sky130_fd_sc_hd__buf_4 output413 (.A(net413),
    .X(master1_wb_ack_i));
 sky130_fd_sc_hd__buf_4 output414 (.A(net414),
    .X(master1_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output415 (.A(net415),
    .X(master1_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output416 (.A(net416),
    .X(master1_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output417 (.A(net417),
    .X(master1_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output418 (.A(net418),
    .X(master1_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output419 (.A(net419),
    .X(master1_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output420 (.A(net420),
    .X(master1_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output421 (.A(net421),
    .X(master1_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output422 (.A(net422),
    .X(master1_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output423 (.A(net423),
    .X(master1_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output424 (.A(net424),
    .X(master1_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output425 (.A(net425),
    .X(master1_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output426 (.A(net426),
    .X(master1_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output427 (.A(net427),
    .X(master1_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output428 (.A(net428),
    .X(master1_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output429 (.A(net429),
    .X(master1_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output430 (.A(net430),
    .X(master1_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output431 (.A(net431),
    .X(master1_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output432 (.A(net432),
    .X(master1_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output433 (.A(net433),
    .X(master1_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output434 (.A(net434),
    .X(master1_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output435 (.A(net435),
    .X(master1_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output436 (.A(net436),
    .X(master1_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output437 (.A(net437),
    .X(master1_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output438 (.A(net438),
    .X(master1_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output439 (.A(net439),
    .X(master1_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output440 (.A(net440),
    .X(master1_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output441 (.A(net441),
    .X(master1_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output442 (.A(net442),
    .X(master1_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output443 (.A(net443),
    .X(master1_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output444 (.A(net444),
    .X(master1_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output445 (.A(net445),
    .X(master1_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output446 (.A(net446),
    .X(master1_wb_error_i));
 sky130_fd_sc_hd__buf_4 output447 (.A(net447),
    .X(master1_wb_stall_i));
 sky130_fd_sc_hd__buf_4 output448 (.A(net448),
    .X(master2_wb_ack_i));
 sky130_fd_sc_hd__buf_4 output449 (.A(net449),
    .X(master2_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output450 (.A(net450),
    .X(master2_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output451 (.A(net451),
    .X(master2_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output452 (.A(net452),
    .X(master2_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output453 (.A(net453),
    .X(master2_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output454 (.A(net454),
    .X(master2_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output455 (.A(net455),
    .X(master2_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output456 (.A(net456),
    .X(master2_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output457 (.A(net457),
    .X(master2_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output458 (.A(net458),
    .X(master2_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output459 (.A(net459),
    .X(master2_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output460 (.A(net460),
    .X(master2_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output461 (.A(net461),
    .X(master2_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output462 (.A(net462),
    .X(master2_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output463 (.A(net463),
    .X(master2_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output464 (.A(net464),
    .X(master2_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output465 (.A(net465),
    .X(master2_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output466 (.A(net466),
    .X(master2_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output467 (.A(net467),
    .X(master2_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output468 (.A(net468),
    .X(master2_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output469 (.A(net469),
    .X(master2_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output470 (.A(net470),
    .X(master2_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output471 (.A(net471),
    .X(master2_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output472 (.A(net472),
    .X(master2_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output473 (.A(net473),
    .X(master2_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output474 (.A(net474),
    .X(master2_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output475 (.A(net475),
    .X(master2_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output476 (.A(net476),
    .X(master2_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output477 (.A(net477),
    .X(master2_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output478 (.A(net478),
    .X(master2_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output479 (.A(net479),
    .X(master2_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output480 (.A(net480),
    .X(master2_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output481 (.A(net481),
    .X(master2_wb_error_i));
 sky130_fd_sc_hd__buf_4 output482 (.A(net482),
    .X(master2_wb_stall_i));
 sky130_fd_sc_hd__buf_4 output483 (.A(net483),
    .X(probe_master0_currentSlave[0]));
 sky130_fd_sc_hd__buf_4 output484 (.A(net484),
    .X(probe_master0_currentSlave[1]));
 sky130_fd_sc_hd__buf_4 output485 (.A(net485),
    .X(probe_master1_currentSlave[0]));
 sky130_fd_sc_hd__buf_4 output486 (.A(net486),
    .X(probe_master1_currentSlave[1]));
 sky130_fd_sc_hd__buf_4 output487 (.A(net487),
    .X(probe_master2_currentSlave[0]));
 sky130_fd_sc_hd__buf_4 output488 (.A(net488),
    .X(probe_master2_currentSlave[1]));
 sky130_fd_sc_hd__buf_4 output489 (.A(net489),
    .X(probe_slave0_currentMaster[0]));
 sky130_fd_sc_hd__buf_4 output490 (.A(net490),
    .X(probe_slave0_currentMaster[1]));
 sky130_fd_sc_hd__buf_4 output491 (.A(net491),
    .X(probe_slave1_currentMaster[0]));
 sky130_fd_sc_hd__buf_4 output492 (.A(net912),
    .X(probe_slave1_currentMaster[1]));
 sky130_fd_sc_hd__buf_4 output493 (.A(net493),
    .X(probe_slave2_currentMaster[0]));
 sky130_fd_sc_hd__buf_4 output494 (.A(net494),
    .X(probe_slave2_currentMaster[1]));
 sky130_fd_sc_hd__buf_4 output495 (.A(net495),
    .X(probe_slave3_currentMaster[0]));
 sky130_fd_sc_hd__buf_4 output496 (.A(net892),
    .X(probe_slave3_currentMaster[1]));
 sky130_fd_sc_hd__buf_4 output497 (.A(net497),
    .X(slave0_wb_adr_i[0]));
 sky130_fd_sc_hd__buf_4 output498 (.A(net498),
    .X(slave0_wb_adr_i[10]));
 sky130_fd_sc_hd__buf_4 output499 (.A(net499),
    .X(slave0_wb_adr_i[11]));
 sky130_fd_sc_hd__buf_4 output500 (.A(net500),
    .X(slave0_wb_adr_i[12]));
 sky130_fd_sc_hd__buf_4 output501 (.A(net501),
    .X(slave0_wb_adr_i[13]));
 sky130_fd_sc_hd__buf_4 output502 (.A(net502),
    .X(slave0_wb_adr_i[14]));
 sky130_fd_sc_hd__buf_4 output503 (.A(net503),
    .X(slave0_wb_adr_i[15]));
 sky130_fd_sc_hd__buf_4 output504 (.A(net504),
    .X(slave0_wb_adr_i[16]));
 sky130_fd_sc_hd__buf_4 output505 (.A(net505),
    .X(slave0_wb_adr_i[17]));
 sky130_fd_sc_hd__buf_4 output506 (.A(net506),
    .X(slave0_wb_adr_i[18]));
 sky130_fd_sc_hd__buf_4 output507 (.A(net507),
    .X(slave0_wb_adr_i[19]));
 sky130_fd_sc_hd__buf_4 output508 (.A(net508),
    .X(slave0_wb_adr_i[1]));
 sky130_fd_sc_hd__buf_4 output509 (.A(net509),
    .X(slave0_wb_adr_i[20]));
 sky130_fd_sc_hd__buf_4 output510 (.A(net510),
    .X(slave0_wb_adr_i[21]));
 sky130_fd_sc_hd__buf_4 output511 (.A(net511),
    .X(slave0_wb_adr_i[22]));
 sky130_fd_sc_hd__buf_4 output512 (.A(net512),
    .X(slave0_wb_adr_i[23]));
 sky130_fd_sc_hd__buf_4 output513 (.A(net513),
    .X(slave0_wb_adr_i[2]));
 sky130_fd_sc_hd__buf_4 output514 (.A(net514),
    .X(slave0_wb_adr_i[3]));
 sky130_fd_sc_hd__buf_4 output515 (.A(net515),
    .X(slave0_wb_adr_i[4]));
 sky130_fd_sc_hd__buf_4 output516 (.A(net516),
    .X(slave0_wb_adr_i[5]));
 sky130_fd_sc_hd__buf_4 output517 (.A(net517),
    .X(slave0_wb_adr_i[6]));
 sky130_fd_sc_hd__buf_4 output518 (.A(net518),
    .X(slave0_wb_adr_i[7]));
 sky130_fd_sc_hd__buf_4 output519 (.A(net519),
    .X(slave0_wb_adr_i[8]));
 sky130_fd_sc_hd__buf_4 output520 (.A(net520),
    .X(slave0_wb_adr_i[9]));
 sky130_fd_sc_hd__buf_4 output521 (.A(net521),
    .X(slave0_wb_cyc_i));
 sky130_fd_sc_hd__buf_4 output522 (.A(net522),
    .X(slave0_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output523 (.A(net523),
    .X(slave0_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output524 (.A(net524),
    .X(slave0_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output525 (.A(net525),
    .X(slave0_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output526 (.A(net526),
    .X(slave0_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output527 (.A(net527),
    .X(slave0_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output528 (.A(net528),
    .X(slave0_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output529 (.A(net529),
    .X(slave0_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output530 (.A(net530),
    .X(slave0_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output531 (.A(net531),
    .X(slave0_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output532 (.A(net532),
    .X(slave0_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output533 (.A(net533),
    .X(slave0_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output534 (.A(net534),
    .X(slave0_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output535 (.A(net535),
    .X(slave0_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output536 (.A(net536),
    .X(slave0_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output537 (.A(net537),
    .X(slave0_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output538 (.A(net538),
    .X(slave0_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output539 (.A(net539),
    .X(slave0_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output540 (.A(net540),
    .X(slave0_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output541 (.A(net541),
    .X(slave0_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output542 (.A(net542),
    .X(slave0_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output543 (.A(net543),
    .X(slave0_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output544 (.A(net544),
    .X(slave0_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output545 (.A(net545),
    .X(slave0_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output546 (.A(net546),
    .X(slave0_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output547 (.A(net547),
    .X(slave0_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output548 (.A(net548),
    .X(slave0_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output549 (.A(net549),
    .X(slave0_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output550 (.A(net550),
    .X(slave0_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output551 (.A(net551),
    .X(slave0_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output552 (.A(net552),
    .X(slave0_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output553 (.A(net553),
    .X(slave0_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output554 (.A(net554),
    .X(slave0_wb_sel_i[0]));
 sky130_fd_sc_hd__buf_4 output555 (.A(net555),
    .X(slave0_wb_sel_i[1]));
 sky130_fd_sc_hd__buf_4 output556 (.A(net556),
    .X(slave0_wb_sel_i[2]));
 sky130_fd_sc_hd__buf_4 output557 (.A(net557),
    .X(slave0_wb_sel_i[3]));
 sky130_fd_sc_hd__buf_4 output558 (.A(net558),
    .X(slave0_wb_stb_i));
 sky130_fd_sc_hd__buf_4 output559 (.A(net559),
    .X(slave0_wb_we_i));
 sky130_fd_sc_hd__buf_4 output560 (.A(net560),
    .X(slave1_wb_adr_i[0]));
 sky130_fd_sc_hd__buf_4 output561 (.A(net561),
    .X(slave1_wb_adr_i[10]));
 sky130_fd_sc_hd__buf_4 output562 (.A(net562),
    .X(slave1_wb_adr_i[11]));
 sky130_fd_sc_hd__buf_4 output563 (.A(net563),
    .X(slave1_wb_adr_i[12]));
 sky130_fd_sc_hd__buf_4 output564 (.A(net564),
    .X(slave1_wb_adr_i[13]));
 sky130_fd_sc_hd__buf_4 output565 (.A(net565),
    .X(slave1_wb_adr_i[14]));
 sky130_fd_sc_hd__buf_4 output566 (.A(net566),
    .X(slave1_wb_adr_i[15]));
 sky130_fd_sc_hd__buf_4 output567 (.A(net567),
    .X(slave1_wb_adr_i[16]));
 sky130_fd_sc_hd__buf_4 output568 (.A(net568),
    .X(slave1_wb_adr_i[17]));
 sky130_fd_sc_hd__buf_4 output569 (.A(net569),
    .X(slave1_wb_adr_i[18]));
 sky130_fd_sc_hd__buf_4 output570 (.A(net570),
    .X(slave1_wb_adr_i[19]));
 sky130_fd_sc_hd__buf_4 output571 (.A(net571),
    .X(slave1_wb_adr_i[1]));
 sky130_fd_sc_hd__buf_4 output572 (.A(net572),
    .X(slave1_wb_adr_i[20]));
 sky130_fd_sc_hd__buf_4 output573 (.A(net573),
    .X(slave1_wb_adr_i[21]));
 sky130_fd_sc_hd__buf_4 output574 (.A(net574),
    .X(slave1_wb_adr_i[22]));
 sky130_fd_sc_hd__buf_4 output575 (.A(net575),
    .X(slave1_wb_adr_i[23]));
 sky130_fd_sc_hd__buf_4 output576 (.A(net576),
    .X(slave1_wb_adr_i[2]));
 sky130_fd_sc_hd__buf_4 output577 (.A(net577),
    .X(slave1_wb_adr_i[3]));
 sky130_fd_sc_hd__buf_4 output578 (.A(net578),
    .X(slave1_wb_adr_i[4]));
 sky130_fd_sc_hd__buf_4 output579 (.A(net579),
    .X(slave1_wb_adr_i[5]));
 sky130_fd_sc_hd__buf_4 output580 (.A(net580),
    .X(slave1_wb_adr_i[6]));
 sky130_fd_sc_hd__buf_4 output581 (.A(net581),
    .X(slave1_wb_adr_i[7]));
 sky130_fd_sc_hd__buf_4 output582 (.A(net582),
    .X(slave1_wb_adr_i[8]));
 sky130_fd_sc_hd__buf_4 output583 (.A(net583),
    .X(slave1_wb_adr_i[9]));
 sky130_fd_sc_hd__buf_4 output584 (.A(net584),
    .X(slave1_wb_cyc_i));
 sky130_fd_sc_hd__buf_4 output585 (.A(net585),
    .X(slave1_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output586 (.A(net586),
    .X(slave1_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output587 (.A(net587),
    .X(slave1_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output588 (.A(net588),
    .X(slave1_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output589 (.A(net589),
    .X(slave1_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output590 (.A(net590),
    .X(slave1_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output591 (.A(net591),
    .X(slave1_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output592 (.A(net592),
    .X(slave1_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output593 (.A(net593),
    .X(slave1_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output594 (.A(net594),
    .X(slave1_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output595 (.A(net595),
    .X(slave1_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output596 (.A(net596),
    .X(slave1_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output597 (.A(net597),
    .X(slave1_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output598 (.A(net598),
    .X(slave1_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output599 (.A(net599),
    .X(slave1_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output600 (.A(net600),
    .X(slave1_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output601 (.A(net601),
    .X(slave1_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output602 (.A(net602),
    .X(slave1_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output603 (.A(net603),
    .X(slave1_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output604 (.A(net604),
    .X(slave1_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output605 (.A(net605),
    .X(slave1_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output606 (.A(net606),
    .X(slave1_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output607 (.A(net607),
    .X(slave1_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output608 (.A(net608),
    .X(slave1_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output609 (.A(net609),
    .X(slave1_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output610 (.A(net610),
    .X(slave1_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output611 (.A(net611),
    .X(slave1_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output612 (.A(net612),
    .X(slave1_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output613 (.A(net613),
    .X(slave1_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output614 (.A(net614),
    .X(slave1_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output615 (.A(net615),
    .X(slave1_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output616 (.A(net616),
    .X(slave1_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output617 (.A(net617),
    .X(slave1_wb_sel_i[0]));
 sky130_fd_sc_hd__buf_4 output618 (.A(net618),
    .X(slave1_wb_sel_i[1]));
 sky130_fd_sc_hd__buf_4 output619 (.A(net619),
    .X(slave1_wb_sel_i[2]));
 sky130_fd_sc_hd__buf_4 output620 (.A(net620),
    .X(slave1_wb_sel_i[3]));
 sky130_fd_sc_hd__buf_4 output621 (.A(net621),
    .X(slave1_wb_stb_i));
 sky130_fd_sc_hd__buf_4 output622 (.A(net622),
    .X(slave1_wb_we_i));
 sky130_fd_sc_hd__buf_4 output623 (.A(net623),
    .X(slave2_wb_adr_i[0]));
 sky130_fd_sc_hd__buf_4 output624 (.A(net624),
    .X(slave2_wb_adr_i[10]));
 sky130_fd_sc_hd__buf_4 output625 (.A(net625),
    .X(slave2_wb_adr_i[11]));
 sky130_fd_sc_hd__buf_4 output626 (.A(net626),
    .X(slave2_wb_adr_i[12]));
 sky130_fd_sc_hd__buf_4 output627 (.A(net627),
    .X(slave2_wb_adr_i[13]));
 sky130_fd_sc_hd__buf_4 output628 (.A(net628),
    .X(slave2_wb_adr_i[14]));
 sky130_fd_sc_hd__buf_4 output629 (.A(net629),
    .X(slave2_wb_adr_i[15]));
 sky130_fd_sc_hd__buf_4 output630 (.A(net630),
    .X(slave2_wb_adr_i[16]));
 sky130_fd_sc_hd__buf_4 output631 (.A(net631),
    .X(slave2_wb_adr_i[17]));
 sky130_fd_sc_hd__buf_4 output632 (.A(net632),
    .X(slave2_wb_adr_i[18]));
 sky130_fd_sc_hd__buf_4 output633 (.A(net633),
    .X(slave2_wb_adr_i[19]));
 sky130_fd_sc_hd__buf_4 output634 (.A(net634),
    .X(slave2_wb_adr_i[1]));
 sky130_fd_sc_hd__buf_4 output635 (.A(net635),
    .X(slave2_wb_adr_i[20]));
 sky130_fd_sc_hd__buf_4 output636 (.A(net636),
    .X(slave2_wb_adr_i[21]));
 sky130_fd_sc_hd__buf_4 output637 (.A(net637),
    .X(slave2_wb_adr_i[22]));
 sky130_fd_sc_hd__buf_4 output638 (.A(net638),
    .X(slave2_wb_adr_i[23]));
 sky130_fd_sc_hd__buf_4 output639 (.A(net639),
    .X(slave2_wb_adr_i[2]));
 sky130_fd_sc_hd__buf_4 output640 (.A(net640),
    .X(slave2_wb_adr_i[3]));
 sky130_fd_sc_hd__buf_4 output641 (.A(net641),
    .X(slave2_wb_adr_i[4]));
 sky130_fd_sc_hd__buf_4 output642 (.A(net642),
    .X(slave2_wb_adr_i[5]));
 sky130_fd_sc_hd__buf_4 output643 (.A(net643),
    .X(slave2_wb_adr_i[6]));
 sky130_fd_sc_hd__buf_4 output644 (.A(net644),
    .X(slave2_wb_adr_i[7]));
 sky130_fd_sc_hd__buf_4 output645 (.A(net645),
    .X(slave2_wb_adr_i[8]));
 sky130_fd_sc_hd__buf_4 output646 (.A(net646),
    .X(slave2_wb_adr_i[9]));
 sky130_fd_sc_hd__buf_4 output647 (.A(net647),
    .X(slave2_wb_cyc_i));
 sky130_fd_sc_hd__buf_4 output648 (.A(net648),
    .X(slave2_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output649 (.A(net649),
    .X(slave2_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output650 (.A(net650),
    .X(slave2_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output651 (.A(net651),
    .X(slave2_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output652 (.A(net652),
    .X(slave2_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output653 (.A(net653),
    .X(slave2_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output654 (.A(net654),
    .X(slave2_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output655 (.A(net655),
    .X(slave2_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output656 (.A(net656),
    .X(slave2_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output657 (.A(net657),
    .X(slave2_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output658 (.A(net658),
    .X(slave2_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output659 (.A(net659),
    .X(slave2_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output660 (.A(net660),
    .X(slave2_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output661 (.A(net661),
    .X(slave2_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output662 (.A(net662),
    .X(slave2_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output663 (.A(net663),
    .X(slave2_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output664 (.A(net664),
    .X(slave2_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output665 (.A(net665),
    .X(slave2_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output666 (.A(net666),
    .X(slave2_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output667 (.A(net667),
    .X(slave2_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output668 (.A(net668),
    .X(slave2_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output669 (.A(net669),
    .X(slave2_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output670 (.A(net670),
    .X(slave2_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output671 (.A(net671),
    .X(slave2_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output672 (.A(net672),
    .X(slave2_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output673 (.A(net673),
    .X(slave2_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output674 (.A(net674),
    .X(slave2_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output675 (.A(net675),
    .X(slave2_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output676 (.A(net676),
    .X(slave2_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output677 (.A(net677),
    .X(slave2_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output678 (.A(net678),
    .X(slave2_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output679 (.A(net679),
    .X(slave2_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output680 (.A(net680),
    .X(slave2_wb_sel_i[0]));
 sky130_fd_sc_hd__buf_4 output681 (.A(net681),
    .X(slave2_wb_sel_i[1]));
 sky130_fd_sc_hd__buf_4 output682 (.A(net682),
    .X(slave2_wb_sel_i[2]));
 sky130_fd_sc_hd__buf_4 output683 (.A(net683),
    .X(slave2_wb_sel_i[3]));
 sky130_fd_sc_hd__buf_4 output684 (.A(net684),
    .X(slave2_wb_stb_i));
 sky130_fd_sc_hd__buf_4 output685 (.A(net685),
    .X(slave2_wb_we_i));
 sky130_fd_sc_hd__buf_4 output686 (.A(net686),
    .X(slave3_wb_adr_i[0]));
 sky130_fd_sc_hd__buf_4 output687 (.A(net687),
    .X(slave3_wb_adr_i[10]));
 sky130_fd_sc_hd__buf_4 output688 (.A(net688),
    .X(slave3_wb_adr_i[11]));
 sky130_fd_sc_hd__buf_4 output689 (.A(net689),
    .X(slave3_wb_adr_i[12]));
 sky130_fd_sc_hd__buf_4 output690 (.A(net690),
    .X(slave3_wb_adr_i[13]));
 sky130_fd_sc_hd__buf_4 output691 (.A(net691),
    .X(slave3_wb_adr_i[14]));
 sky130_fd_sc_hd__buf_4 output692 (.A(net692),
    .X(slave3_wb_adr_i[15]));
 sky130_fd_sc_hd__buf_4 output693 (.A(net693),
    .X(slave3_wb_adr_i[16]));
 sky130_fd_sc_hd__buf_4 output694 (.A(net694),
    .X(slave3_wb_adr_i[17]));
 sky130_fd_sc_hd__buf_4 output695 (.A(net695),
    .X(slave3_wb_adr_i[18]));
 sky130_fd_sc_hd__buf_4 output696 (.A(net696),
    .X(slave3_wb_adr_i[19]));
 sky130_fd_sc_hd__buf_4 output697 (.A(net697),
    .X(slave3_wb_adr_i[1]));
 sky130_fd_sc_hd__buf_4 output698 (.A(net698),
    .X(slave3_wb_adr_i[20]));
 sky130_fd_sc_hd__buf_4 output699 (.A(net699),
    .X(slave3_wb_adr_i[21]));
 sky130_fd_sc_hd__buf_4 output700 (.A(net700),
    .X(slave3_wb_adr_i[22]));
 sky130_fd_sc_hd__buf_4 output701 (.A(net701),
    .X(slave3_wb_adr_i[23]));
 sky130_fd_sc_hd__buf_4 output702 (.A(net702),
    .X(slave3_wb_adr_i[2]));
 sky130_fd_sc_hd__buf_4 output703 (.A(net703),
    .X(slave3_wb_adr_i[3]));
 sky130_fd_sc_hd__buf_4 output704 (.A(net704),
    .X(slave3_wb_adr_i[4]));
 sky130_fd_sc_hd__buf_4 output705 (.A(net705),
    .X(slave3_wb_adr_i[5]));
 sky130_fd_sc_hd__buf_4 output706 (.A(net706),
    .X(slave3_wb_adr_i[6]));
 sky130_fd_sc_hd__buf_4 output707 (.A(net707),
    .X(slave3_wb_adr_i[7]));
 sky130_fd_sc_hd__buf_4 output708 (.A(net708),
    .X(slave3_wb_adr_i[8]));
 sky130_fd_sc_hd__buf_4 output709 (.A(net709),
    .X(slave3_wb_adr_i[9]));
 sky130_fd_sc_hd__buf_4 output710 (.A(net710),
    .X(slave3_wb_cyc_i));
 sky130_fd_sc_hd__buf_4 output711 (.A(net711),
    .X(slave3_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output712 (.A(net712),
    .X(slave3_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output713 (.A(net713),
    .X(slave3_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output714 (.A(net714),
    .X(slave3_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output715 (.A(net715),
    .X(slave3_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output716 (.A(net716),
    .X(slave3_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output717 (.A(net717),
    .X(slave3_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output718 (.A(net718),
    .X(slave3_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output719 (.A(net719),
    .X(slave3_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output720 (.A(net720),
    .X(slave3_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output721 (.A(net721),
    .X(slave3_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output722 (.A(net722),
    .X(slave3_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output723 (.A(net723),
    .X(slave3_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output724 (.A(net724),
    .X(slave3_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output725 (.A(net725),
    .X(slave3_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output726 (.A(net726),
    .X(slave3_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output727 (.A(net727),
    .X(slave3_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output728 (.A(net728),
    .X(slave3_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output729 (.A(net729),
    .X(slave3_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output730 (.A(net730),
    .X(slave3_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output731 (.A(net731),
    .X(slave3_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output732 (.A(net732),
    .X(slave3_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output733 (.A(net733),
    .X(slave3_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output734 (.A(net734),
    .X(slave3_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output735 (.A(net735),
    .X(slave3_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output736 (.A(net736),
    .X(slave3_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output737 (.A(net737),
    .X(slave3_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output738 (.A(net738),
    .X(slave3_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output739 (.A(net739),
    .X(slave3_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output740 (.A(net740),
    .X(slave3_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output741 (.A(net741),
    .X(slave3_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output742 (.A(net742),
    .X(slave3_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output743 (.A(net743),
    .X(slave3_wb_sel_i[0]));
 sky130_fd_sc_hd__buf_4 output744 (.A(net744),
    .X(slave3_wb_sel_i[1]));
 sky130_fd_sc_hd__buf_4 output745 (.A(net745),
    .X(slave3_wb_sel_i[2]));
 sky130_fd_sc_hd__buf_4 output746 (.A(net746),
    .X(slave3_wb_sel_i[3]));
 sky130_fd_sc_hd__buf_4 output747 (.A(net747),
    .X(slave3_wb_stb_i));
 sky130_fd_sc_hd__buf_4 output748 (.A(net748),
    .X(slave3_wb_we_i));
 sky130_fd_sc_hd__buf_4 output749 (.A(net749),
    .X(slave4_wb_adr_i[0]));
 sky130_fd_sc_hd__buf_4 output750 (.A(net750),
    .X(slave4_wb_adr_i[10]));
 sky130_fd_sc_hd__buf_4 output751 (.A(net751),
    .X(slave4_wb_adr_i[11]));
 sky130_fd_sc_hd__buf_4 output752 (.A(net752),
    .X(slave4_wb_adr_i[12]));
 sky130_fd_sc_hd__buf_4 output753 (.A(net753),
    .X(slave4_wb_adr_i[13]));
 sky130_fd_sc_hd__buf_4 output754 (.A(net754),
    .X(slave4_wb_adr_i[14]));
 sky130_fd_sc_hd__buf_4 output755 (.A(net755),
    .X(slave4_wb_adr_i[15]));
 sky130_fd_sc_hd__buf_4 output756 (.A(net756),
    .X(slave4_wb_adr_i[16]));
 sky130_fd_sc_hd__buf_4 output757 (.A(net757),
    .X(slave4_wb_adr_i[17]));
 sky130_fd_sc_hd__buf_4 output758 (.A(net758),
    .X(slave4_wb_adr_i[18]));
 sky130_fd_sc_hd__buf_4 output759 (.A(net759),
    .X(slave4_wb_adr_i[19]));
 sky130_fd_sc_hd__buf_4 output760 (.A(net760),
    .X(slave4_wb_adr_i[1]));
 sky130_fd_sc_hd__buf_4 output761 (.A(net761),
    .X(slave4_wb_adr_i[20]));
 sky130_fd_sc_hd__buf_4 output762 (.A(net762),
    .X(slave4_wb_adr_i[21]));
 sky130_fd_sc_hd__buf_4 output763 (.A(net763),
    .X(slave4_wb_adr_i[22]));
 sky130_fd_sc_hd__buf_4 output764 (.A(net764),
    .X(slave4_wb_adr_i[23]));
 sky130_fd_sc_hd__buf_4 output765 (.A(net765),
    .X(slave4_wb_adr_i[2]));
 sky130_fd_sc_hd__buf_4 output766 (.A(net766),
    .X(slave4_wb_adr_i[3]));
 sky130_fd_sc_hd__buf_4 output767 (.A(net767),
    .X(slave4_wb_adr_i[4]));
 sky130_fd_sc_hd__buf_4 output768 (.A(net768),
    .X(slave4_wb_adr_i[5]));
 sky130_fd_sc_hd__buf_4 output769 (.A(net769),
    .X(slave4_wb_adr_i[6]));
 sky130_fd_sc_hd__buf_4 output770 (.A(net770),
    .X(slave4_wb_adr_i[7]));
 sky130_fd_sc_hd__buf_4 output771 (.A(net771),
    .X(slave4_wb_adr_i[8]));
 sky130_fd_sc_hd__buf_4 output772 (.A(net772),
    .X(slave4_wb_adr_i[9]));
 sky130_fd_sc_hd__buf_4 output773 (.A(net773),
    .X(slave4_wb_cyc_i));
 sky130_fd_sc_hd__buf_4 output774 (.A(net774),
    .X(slave4_wb_data_i[0]));
 sky130_fd_sc_hd__buf_4 output775 (.A(net775),
    .X(slave4_wb_data_i[10]));
 sky130_fd_sc_hd__buf_4 output776 (.A(net776),
    .X(slave4_wb_data_i[11]));
 sky130_fd_sc_hd__buf_4 output777 (.A(net777),
    .X(slave4_wb_data_i[12]));
 sky130_fd_sc_hd__buf_4 output778 (.A(net778),
    .X(slave4_wb_data_i[13]));
 sky130_fd_sc_hd__buf_4 output779 (.A(net779),
    .X(slave4_wb_data_i[14]));
 sky130_fd_sc_hd__buf_4 output780 (.A(net780),
    .X(slave4_wb_data_i[15]));
 sky130_fd_sc_hd__buf_4 output781 (.A(net781),
    .X(slave4_wb_data_i[16]));
 sky130_fd_sc_hd__buf_4 output782 (.A(net782),
    .X(slave4_wb_data_i[17]));
 sky130_fd_sc_hd__buf_4 output783 (.A(net783),
    .X(slave4_wb_data_i[18]));
 sky130_fd_sc_hd__buf_4 output784 (.A(net784),
    .X(slave4_wb_data_i[19]));
 sky130_fd_sc_hd__buf_4 output785 (.A(net785),
    .X(slave4_wb_data_i[1]));
 sky130_fd_sc_hd__buf_4 output786 (.A(net786),
    .X(slave4_wb_data_i[20]));
 sky130_fd_sc_hd__buf_4 output787 (.A(net787),
    .X(slave4_wb_data_i[21]));
 sky130_fd_sc_hd__buf_4 output788 (.A(net788),
    .X(slave4_wb_data_i[22]));
 sky130_fd_sc_hd__buf_4 output789 (.A(net789),
    .X(slave4_wb_data_i[23]));
 sky130_fd_sc_hd__buf_4 output790 (.A(net790),
    .X(slave4_wb_data_i[24]));
 sky130_fd_sc_hd__buf_4 output791 (.A(net791),
    .X(slave4_wb_data_i[25]));
 sky130_fd_sc_hd__buf_4 output792 (.A(net792),
    .X(slave4_wb_data_i[26]));
 sky130_fd_sc_hd__buf_4 output793 (.A(net793),
    .X(slave4_wb_data_i[27]));
 sky130_fd_sc_hd__buf_4 output794 (.A(net794),
    .X(slave4_wb_data_i[28]));
 sky130_fd_sc_hd__buf_4 output795 (.A(net795),
    .X(slave4_wb_data_i[29]));
 sky130_fd_sc_hd__buf_4 output796 (.A(net796),
    .X(slave4_wb_data_i[2]));
 sky130_fd_sc_hd__buf_4 output797 (.A(net797),
    .X(slave4_wb_data_i[30]));
 sky130_fd_sc_hd__buf_4 output798 (.A(net798),
    .X(slave4_wb_data_i[31]));
 sky130_fd_sc_hd__buf_4 output799 (.A(net799),
    .X(slave4_wb_data_i[3]));
 sky130_fd_sc_hd__buf_4 output800 (.A(net800),
    .X(slave4_wb_data_i[4]));
 sky130_fd_sc_hd__buf_4 output801 (.A(net801),
    .X(slave4_wb_data_i[5]));
 sky130_fd_sc_hd__buf_4 output802 (.A(net802),
    .X(slave4_wb_data_i[6]));
 sky130_fd_sc_hd__buf_4 output803 (.A(net803),
    .X(slave4_wb_data_i[7]));
 sky130_fd_sc_hd__buf_4 output804 (.A(net804),
    .X(slave4_wb_data_i[8]));
 sky130_fd_sc_hd__buf_4 output805 (.A(net805),
    .X(slave4_wb_data_i[9]));
 sky130_fd_sc_hd__buf_4 output806 (.A(net806),
    .X(slave4_wb_sel_i[0]));
 sky130_fd_sc_hd__buf_4 output807 (.A(net807),
    .X(slave4_wb_sel_i[1]));
 sky130_fd_sc_hd__buf_4 output808 (.A(net808),
    .X(slave4_wb_sel_i[2]));
 sky130_fd_sc_hd__buf_4 output809 (.A(net809),
    .X(slave4_wb_sel_i[3]));
 sky130_fd_sc_hd__buf_4 output810 (.A(net810),
    .X(slave4_wb_stb_i));
 sky130_fd_sc_hd__buf_4 output811 (.A(net811),
    .X(slave4_wb_we_i));
 sky130_fd_sc_hd__buf_6 wire960 (.A(_0644_),
    .X(net960));
 sky130_fd_sc_hd__buf_6 wire998 (.A(_0602_),
    .X(net998));
 assign probe_master3_currentSlave[0] = net1017;
 assign probe_master3_currentSlave[1] = net1018;
endmodule

