magic
tech sky130A
magscale 1 2
timestamp 1658164597
<< obsli1 >>
rect 1104 2159 98808 157777
<< obsm1 >>
rect 14 1300 99990 158908
<< metal2 >>
rect 1214 159200 1270 160000
rect 3698 159200 3754 160000
rect 6274 159200 6330 160000
rect 8850 159200 8906 160000
rect 11426 159200 11482 160000
rect 14002 159200 14058 160000
rect 16578 159200 16634 160000
rect 19154 159200 19210 160000
rect 21638 159200 21694 160000
rect 24214 159200 24270 160000
rect 26790 159200 26846 160000
rect 29366 159200 29422 160000
rect 31942 159200 31998 160000
rect 34518 159200 34574 160000
rect 37094 159200 37150 160000
rect 39670 159200 39726 160000
rect 42154 159200 42210 160000
rect 44730 159200 44786 160000
rect 47306 159200 47362 160000
rect 49882 159200 49938 160000
rect 52458 159200 52514 160000
rect 55034 159200 55090 160000
rect 57610 159200 57666 160000
rect 60186 159200 60242 160000
rect 62670 159200 62726 160000
rect 65246 159200 65302 160000
rect 67822 159200 67878 160000
rect 70398 159200 70454 160000
rect 72974 159200 73030 160000
rect 75550 159200 75606 160000
rect 78126 159200 78182 160000
rect 80702 159200 80758 160000
rect 83186 159200 83242 160000
rect 85762 159200 85818 160000
rect 88338 159200 88394 160000
rect 90914 159200 90970 160000
rect 93490 159200 93546 160000
rect 96066 159200 96122 160000
rect 98642 159200 98698 160000
rect 846 0 902 800
rect 2594 0 2650 800
rect 4342 0 4398 800
rect 6182 0 6238 800
rect 7930 0 7986 800
rect 9770 0 9826 800
rect 11518 0 11574 800
rect 13266 0 13322 800
rect 15106 0 15162 800
rect 16854 0 16910 800
rect 18694 0 18750 800
rect 20442 0 20498 800
rect 22190 0 22246 800
rect 24030 0 24086 800
rect 25778 0 25834 800
rect 27618 0 27674 800
rect 29366 0 29422 800
rect 31114 0 31170 800
rect 32954 0 33010 800
rect 34702 0 34758 800
rect 36542 0 36598 800
rect 38290 0 38346 800
rect 40130 0 40186 800
rect 41878 0 41934 800
rect 43626 0 43682 800
rect 45466 0 45522 800
rect 47214 0 47270 800
rect 49054 0 49110 800
rect 50802 0 50858 800
rect 52550 0 52606 800
rect 54390 0 54446 800
rect 56138 0 56194 800
rect 57978 0 58034 800
rect 59726 0 59782 800
rect 61474 0 61530 800
rect 63314 0 63370 800
rect 65062 0 65118 800
rect 66902 0 66958 800
rect 68650 0 68706 800
rect 70490 0 70546 800
rect 72238 0 72294 800
rect 73986 0 74042 800
rect 75826 0 75882 800
rect 77574 0 77630 800
rect 79414 0 79470 800
rect 81162 0 81218 800
rect 82910 0 82966 800
rect 84750 0 84806 800
rect 86498 0 86554 800
rect 88338 0 88394 800
rect 90086 0 90142 800
rect 91834 0 91890 800
rect 93674 0 93730 800
rect 95422 0 95478 800
rect 97262 0 97318 800
rect 99010 0 99066 800
<< obsm2 >>
rect 18 159144 1158 159497
rect 1326 159144 3642 159497
rect 3810 159144 6218 159497
rect 6386 159144 8794 159497
rect 8962 159144 11370 159497
rect 11538 159144 13946 159497
rect 14114 159144 16522 159497
rect 16690 159144 19098 159497
rect 19266 159144 21582 159497
rect 21750 159144 24158 159497
rect 24326 159144 26734 159497
rect 26902 159144 29310 159497
rect 29478 159144 31886 159497
rect 32054 159144 34462 159497
rect 34630 159144 37038 159497
rect 37206 159144 39614 159497
rect 39782 159144 42098 159497
rect 42266 159144 44674 159497
rect 44842 159144 47250 159497
rect 47418 159144 49826 159497
rect 49994 159144 52402 159497
rect 52570 159144 54978 159497
rect 55146 159144 57554 159497
rect 57722 159144 60130 159497
rect 60298 159144 62614 159497
rect 62782 159144 65190 159497
rect 65358 159144 67766 159497
rect 67934 159144 70342 159497
rect 70510 159144 72918 159497
rect 73086 159144 75494 159497
rect 75662 159144 78070 159497
rect 78238 159144 80646 159497
rect 80814 159144 83130 159497
rect 83298 159144 85706 159497
rect 85874 159144 88282 159497
rect 88450 159144 90858 159497
rect 91026 159144 93434 159497
rect 93602 159144 96010 159497
rect 96178 159144 98586 159497
rect 98754 159144 99984 159497
rect 18 856 99984 159144
rect 18 303 790 856
rect 958 303 2538 856
rect 2706 303 4286 856
rect 4454 303 6126 856
rect 6294 303 7874 856
rect 8042 303 9714 856
rect 9882 303 11462 856
rect 11630 303 13210 856
rect 13378 303 15050 856
rect 15218 303 16798 856
rect 16966 303 18638 856
rect 18806 303 20386 856
rect 20554 303 22134 856
rect 22302 303 23974 856
rect 24142 303 25722 856
rect 25890 303 27562 856
rect 27730 303 29310 856
rect 29478 303 31058 856
rect 31226 303 32898 856
rect 33066 303 34646 856
rect 34814 303 36486 856
rect 36654 303 38234 856
rect 38402 303 40074 856
rect 40242 303 41822 856
rect 41990 303 43570 856
rect 43738 303 45410 856
rect 45578 303 47158 856
rect 47326 303 48998 856
rect 49166 303 50746 856
rect 50914 303 52494 856
rect 52662 303 54334 856
rect 54502 303 56082 856
rect 56250 303 57922 856
rect 58090 303 59670 856
rect 59838 303 61418 856
rect 61586 303 63258 856
rect 63426 303 65006 856
rect 65174 303 66846 856
rect 67014 303 68594 856
rect 68762 303 70434 856
rect 70602 303 72182 856
rect 72350 303 73930 856
rect 74098 303 75770 856
rect 75938 303 77518 856
rect 77686 303 79358 856
rect 79526 303 81106 856
rect 81274 303 82854 856
rect 83022 303 84694 856
rect 84862 303 86442 856
rect 86610 303 88282 856
rect 88450 303 90030 856
rect 90198 303 91778 856
rect 91946 303 93618 856
rect 93786 303 95366 856
rect 95534 303 97206 856
rect 97374 303 98954 856
rect 99122 303 99984 856
<< metal3 >>
rect 0 159400 800 159520
rect 99200 159400 100000 159520
rect 0 158584 800 158704
rect 99200 158584 100000 158704
rect 0 157768 800 157888
rect 99200 157768 100000 157888
rect 0 156952 800 157072
rect 99200 156952 100000 157072
rect 0 156136 800 156256
rect 99200 156136 100000 156256
rect 0 155320 800 155440
rect 99200 155456 100000 155576
rect 0 154504 800 154624
rect 99200 154640 100000 154760
rect 0 153688 800 153808
rect 99200 153824 100000 153944
rect 0 152872 800 152992
rect 99200 153008 100000 153128
rect 0 152056 800 152176
rect 99200 152192 100000 152312
rect 99200 151376 100000 151496
rect 0 151104 800 151224
rect 99200 150696 100000 150816
rect 0 150288 800 150408
rect 99200 149880 100000 150000
rect 0 149472 800 149592
rect 99200 149064 100000 149184
rect 0 148656 800 148776
rect 99200 148248 100000 148368
rect 0 147840 800 147960
rect 99200 147432 100000 147552
rect 0 147024 800 147144
rect 99200 146752 100000 146872
rect 0 146208 800 146328
rect 99200 145936 100000 146056
rect 0 145392 800 145512
rect 99200 145120 100000 145240
rect 0 144576 800 144696
rect 99200 144304 100000 144424
rect 0 143760 800 143880
rect 99200 143488 100000 143608
rect 0 142944 800 143064
rect 99200 142672 100000 142792
rect 0 141992 800 142112
rect 99200 141992 100000 142112
rect 0 141176 800 141296
rect 99200 141176 100000 141296
rect 0 140360 800 140480
rect 99200 140360 100000 140480
rect 0 139544 800 139664
rect 99200 139544 100000 139664
rect 0 138728 800 138848
rect 99200 138728 100000 138848
rect 0 137912 800 138032
rect 99200 137912 100000 138032
rect 0 137096 800 137216
rect 99200 137232 100000 137352
rect 0 136280 800 136400
rect 99200 136416 100000 136536
rect 0 135464 800 135584
rect 99200 135600 100000 135720
rect 0 134648 800 134768
rect 99200 134784 100000 134904
rect 0 133832 800 133952
rect 99200 133968 100000 134088
rect 99200 133288 100000 133408
rect 0 132880 800 133000
rect 99200 132472 100000 132592
rect 0 132064 800 132184
rect 99200 131656 100000 131776
rect 0 131248 800 131368
rect 99200 130840 100000 130960
rect 0 130432 800 130552
rect 99200 130024 100000 130144
rect 0 129616 800 129736
rect 99200 129208 100000 129328
rect 0 128800 800 128920
rect 99200 128528 100000 128648
rect 0 127984 800 128104
rect 99200 127712 100000 127832
rect 0 127168 800 127288
rect 99200 126896 100000 127016
rect 0 126352 800 126472
rect 99200 126080 100000 126200
rect 0 125536 800 125656
rect 99200 125264 100000 125384
rect 0 124584 800 124704
rect 99200 124584 100000 124704
rect 0 123768 800 123888
rect 99200 123768 100000 123888
rect 0 122952 800 123072
rect 99200 122952 100000 123072
rect 0 122136 800 122256
rect 99200 122136 100000 122256
rect 0 121320 800 121440
rect 99200 121320 100000 121440
rect 0 120504 800 120624
rect 99200 120504 100000 120624
rect 0 119688 800 119808
rect 99200 119824 100000 119944
rect 0 118872 800 118992
rect 99200 119008 100000 119128
rect 0 118056 800 118176
rect 99200 118192 100000 118312
rect 0 117240 800 117360
rect 99200 117376 100000 117496
rect 0 116424 800 116544
rect 99200 116560 100000 116680
rect 99200 115744 100000 115864
rect 0 115472 800 115592
rect 99200 115064 100000 115184
rect 0 114656 800 114776
rect 99200 114248 100000 114368
rect 0 113840 800 113960
rect 99200 113432 100000 113552
rect 0 113024 800 113144
rect 99200 112616 100000 112736
rect 0 112208 800 112328
rect 99200 111800 100000 111920
rect 0 111392 800 111512
rect 99200 111120 100000 111240
rect 0 110576 800 110696
rect 99200 110304 100000 110424
rect 0 109760 800 109880
rect 99200 109488 100000 109608
rect 0 108944 800 109064
rect 99200 108672 100000 108792
rect 0 108128 800 108248
rect 99200 107856 100000 107976
rect 0 107312 800 107432
rect 99200 107040 100000 107160
rect 0 106360 800 106480
rect 99200 106360 100000 106480
rect 0 105544 800 105664
rect 99200 105544 100000 105664
rect 0 104728 800 104848
rect 99200 104728 100000 104848
rect 0 103912 800 104032
rect 99200 103912 100000 104032
rect 0 103096 800 103216
rect 99200 103096 100000 103216
rect 0 102280 800 102400
rect 99200 102416 100000 102536
rect 0 101464 800 101584
rect 99200 101600 100000 101720
rect 0 100648 800 100768
rect 99200 100784 100000 100904
rect 0 99832 800 99952
rect 99200 99968 100000 100088
rect 0 99016 800 99136
rect 99200 99152 100000 99272
rect 0 98200 800 98320
rect 99200 98336 100000 98456
rect 99200 97656 100000 97776
rect 0 97248 800 97368
rect 99200 96840 100000 96960
rect 0 96432 800 96552
rect 99200 96024 100000 96144
rect 0 95616 800 95736
rect 99200 95208 100000 95328
rect 0 94800 800 94920
rect 99200 94392 100000 94512
rect 0 93984 800 94104
rect 99200 93576 100000 93696
rect 0 93168 800 93288
rect 99200 92896 100000 93016
rect 0 92352 800 92472
rect 99200 92080 100000 92200
rect 0 91536 800 91656
rect 99200 91264 100000 91384
rect 0 90720 800 90840
rect 99200 90448 100000 90568
rect 0 89904 800 90024
rect 99200 89632 100000 89752
rect 0 88952 800 89072
rect 99200 88952 100000 89072
rect 0 88136 800 88256
rect 99200 88136 100000 88256
rect 0 87320 800 87440
rect 99200 87320 100000 87440
rect 0 86504 800 86624
rect 99200 86504 100000 86624
rect 0 85688 800 85808
rect 99200 85688 100000 85808
rect 0 84872 800 84992
rect 99200 84872 100000 84992
rect 0 84056 800 84176
rect 99200 84192 100000 84312
rect 0 83240 800 83360
rect 99200 83376 100000 83496
rect 0 82424 800 82544
rect 99200 82560 100000 82680
rect 0 81608 800 81728
rect 99200 81744 100000 81864
rect 0 80792 800 80912
rect 99200 80928 100000 81048
rect 99200 80248 100000 80368
rect 0 79840 800 79960
rect 99200 79432 100000 79552
rect 0 79024 800 79144
rect 99200 78616 100000 78736
rect 0 78208 800 78328
rect 99200 77800 100000 77920
rect 0 77392 800 77512
rect 99200 76984 100000 77104
rect 0 76576 800 76696
rect 99200 76168 100000 76288
rect 0 75760 800 75880
rect 99200 75488 100000 75608
rect 0 74944 800 75064
rect 99200 74672 100000 74792
rect 0 74128 800 74248
rect 99200 73856 100000 73976
rect 0 73312 800 73432
rect 99200 73040 100000 73160
rect 0 72496 800 72616
rect 99200 72224 100000 72344
rect 0 71680 800 71800
rect 99200 71408 100000 71528
rect 0 70728 800 70848
rect 99200 70728 100000 70848
rect 0 69912 800 70032
rect 99200 69912 100000 70032
rect 0 69096 800 69216
rect 99200 69096 100000 69216
rect 0 68280 800 68400
rect 99200 68280 100000 68400
rect 0 67464 800 67584
rect 99200 67464 100000 67584
rect 0 66648 800 66768
rect 99200 66784 100000 66904
rect 0 65832 800 65952
rect 99200 65968 100000 66088
rect 0 65016 800 65136
rect 99200 65152 100000 65272
rect 0 64200 800 64320
rect 99200 64336 100000 64456
rect 0 63384 800 63504
rect 99200 63520 100000 63640
rect 99200 62704 100000 62824
rect 0 62432 800 62552
rect 99200 62024 100000 62144
rect 0 61616 800 61736
rect 99200 61208 100000 61328
rect 0 60800 800 60920
rect 99200 60392 100000 60512
rect 0 59984 800 60104
rect 99200 59576 100000 59696
rect 0 59168 800 59288
rect 99200 58760 100000 58880
rect 0 58352 800 58472
rect 99200 57944 100000 58064
rect 0 57536 800 57656
rect 99200 57264 100000 57384
rect 0 56720 800 56840
rect 99200 56448 100000 56568
rect 0 55904 800 56024
rect 99200 55632 100000 55752
rect 0 55088 800 55208
rect 99200 54816 100000 54936
rect 0 54272 800 54392
rect 99200 54000 100000 54120
rect 0 53320 800 53440
rect 99200 53320 100000 53440
rect 0 52504 800 52624
rect 99200 52504 100000 52624
rect 0 51688 800 51808
rect 99200 51688 100000 51808
rect 0 50872 800 50992
rect 99200 50872 100000 50992
rect 0 50056 800 50176
rect 99200 50056 100000 50176
rect 0 49240 800 49360
rect 99200 49240 100000 49360
rect 0 48424 800 48544
rect 99200 48560 100000 48680
rect 0 47608 800 47728
rect 99200 47744 100000 47864
rect 0 46792 800 46912
rect 99200 46928 100000 47048
rect 0 45976 800 46096
rect 99200 46112 100000 46232
rect 0 45160 800 45280
rect 99200 45296 100000 45416
rect 99200 44616 100000 44736
rect 0 44208 800 44328
rect 99200 43800 100000 43920
rect 0 43392 800 43512
rect 99200 42984 100000 43104
rect 0 42576 800 42696
rect 99200 42168 100000 42288
rect 0 41760 800 41880
rect 99200 41352 100000 41472
rect 0 40944 800 41064
rect 99200 40536 100000 40656
rect 0 40128 800 40248
rect 99200 39856 100000 39976
rect 0 39312 800 39432
rect 99200 39040 100000 39160
rect 0 38496 800 38616
rect 99200 38224 100000 38344
rect 0 37680 800 37800
rect 99200 37408 100000 37528
rect 0 36864 800 36984
rect 99200 36592 100000 36712
rect 0 36048 800 36168
rect 99200 35776 100000 35896
rect 0 35096 800 35216
rect 99200 35096 100000 35216
rect 0 34280 800 34400
rect 99200 34280 100000 34400
rect 0 33464 800 33584
rect 99200 33464 100000 33584
rect 0 32648 800 32768
rect 99200 32648 100000 32768
rect 0 31832 800 31952
rect 99200 31832 100000 31952
rect 0 31016 800 31136
rect 99200 31152 100000 31272
rect 0 30200 800 30320
rect 99200 30336 100000 30456
rect 0 29384 800 29504
rect 99200 29520 100000 29640
rect 0 28568 800 28688
rect 99200 28704 100000 28824
rect 0 27752 800 27872
rect 99200 27888 100000 28008
rect 99200 27072 100000 27192
rect 0 26800 800 26920
rect 99200 26392 100000 26512
rect 0 25984 800 26104
rect 99200 25576 100000 25696
rect 0 25168 800 25288
rect 99200 24760 100000 24880
rect 0 24352 800 24472
rect 99200 23944 100000 24064
rect 0 23536 800 23656
rect 99200 23128 100000 23248
rect 0 22720 800 22840
rect 99200 22448 100000 22568
rect 0 21904 800 22024
rect 99200 21632 100000 21752
rect 0 21088 800 21208
rect 99200 20816 100000 20936
rect 0 20272 800 20392
rect 99200 20000 100000 20120
rect 0 19456 800 19576
rect 99200 19184 100000 19304
rect 0 18640 800 18760
rect 99200 18368 100000 18488
rect 0 17688 800 17808
rect 99200 17688 100000 17808
rect 0 16872 800 16992
rect 99200 16872 100000 16992
rect 0 16056 800 16176
rect 99200 16056 100000 16176
rect 0 15240 800 15360
rect 99200 15240 100000 15360
rect 0 14424 800 14544
rect 99200 14424 100000 14544
rect 0 13608 800 13728
rect 99200 13608 100000 13728
rect 0 12792 800 12912
rect 99200 12928 100000 13048
rect 0 11976 800 12096
rect 99200 12112 100000 12232
rect 0 11160 800 11280
rect 99200 11296 100000 11416
rect 0 10344 800 10464
rect 99200 10480 100000 10600
rect 0 9528 800 9648
rect 99200 9664 100000 9784
rect 99200 8984 100000 9104
rect 0 8576 800 8696
rect 99200 8168 100000 8288
rect 0 7760 800 7880
rect 99200 7352 100000 7472
rect 0 6944 800 7064
rect 99200 6536 100000 6656
rect 0 6128 800 6248
rect 99200 5720 100000 5840
rect 0 5312 800 5432
rect 99200 4904 100000 5024
rect 0 4496 800 4616
rect 99200 4224 100000 4344
rect 0 3680 800 3800
rect 99200 3408 100000 3528
rect 0 2864 800 2984
rect 99200 2592 100000 2712
rect 0 2048 800 2168
rect 99200 1776 100000 1896
rect 0 1232 800 1352
rect 99200 960 100000 1080
rect 0 416 800 536
rect 99200 280 100000 400
<< obsm3 >>
rect 880 159320 99120 159493
rect 13 158784 99899 159320
rect 880 158504 99120 158784
rect 13 157968 99899 158504
rect 880 157688 99120 157968
rect 13 157152 99899 157688
rect 880 156872 99120 157152
rect 13 156336 99899 156872
rect 880 156056 99120 156336
rect 13 155656 99899 156056
rect 13 155520 99120 155656
rect 880 155376 99120 155520
rect 880 155240 99899 155376
rect 13 154840 99899 155240
rect 13 154704 99120 154840
rect 880 154560 99120 154704
rect 880 154424 99899 154560
rect 13 154024 99899 154424
rect 13 153888 99120 154024
rect 880 153744 99120 153888
rect 880 153608 99899 153744
rect 13 153208 99899 153608
rect 13 153072 99120 153208
rect 880 152928 99120 153072
rect 880 152792 99899 152928
rect 13 152392 99899 152792
rect 13 152256 99120 152392
rect 880 152112 99120 152256
rect 880 151976 99899 152112
rect 13 151576 99899 151976
rect 13 151304 99120 151576
rect 880 151296 99120 151304
rect 880 151024 99899 151296
rect 13 150896 99899 151024
rect 13 150616 99120 150896
rect 13 150488 99899 150616
rect 880 150208 99899 150488
rect 13 150080 99899 150208
rect 13 149800 99120 150080
rect 13 149672 99899 149800
rect 880 149392 99899 149672
rect 13 149264 99899 149392
rect 13 148984 99120 149264
rect 13 148856 99899 148984
rect 880 148576 99899 148856
rect 13 148448 99899 148576
rect 13 148168 99120 148448
rect 13 148040 99899 148168
rect 880 147760 99899 148040
rect 13 147632 99899 147760
rect 13 147352 99120 147632
rect 13 147224 99899 147352
rect 880 146952 99899 147224
rect 880 146944 99120 146952
rect 13 146672 99120 146944
rect 13 146408 99899 146672
rect 880 146136 99899 146408
rect 880 146128 99120 146136
rect 13 145856 99120 146128
rect 13 145592 99899 145856
rect 880 145320 99899 145592
rect 880 145312 99120 145320
rect 13 145040 99120 145312
rect 13 144776 99899 145040
rect 880 144504 99899 144776
rect 880 144496 99120 144504
rect 13 144224 99120 144496
rect 13 143960 99899 144224
rect 880 143688 99899 143960
rect 880 143680 99120 143688
rect 13 143408 99120 143680
rect 13 143144 99899 143408
rect 880 142872 99899 143144
rect 880 142864 99120 142872
rect 13 142592 99120 142864
rect 13 142192 99899 142592
rect 880 141912 99120 142192
rect 13 141376 99899 141912
rect 880 141096 99120 141376
rect 13 140560 99899 141096
rect 880 140280 99120 140560
rect 13 139744 99899 140280
rect 880 139464 99120 139744
rect 13 138928 99899 139464
rect 880 138648 99120 138928
rect 13 138112 99899 138648
rect 880 137832 99120 138112
rect 13 137432 99899 137832
rect 13 137296 99120 137432
rect 880 137152 99120 137296
rect 880 137016 99899 137152
rect 13 136616 99899 137016
rect 13 136480 99120 136616
rect 880 136336 99120 136480
rect 880 136200 99899 136336
rect 13 135800 99899 136200
rect 13 135664 99120 135800
rect 880 135520 99120 135664
rect 880 135384 99899 135520
rect 13 134984 99899 135384
rect 13 134848 99120 134984
rect 880 134704 99120 134848
rect 880 134568 99899 134704
rect 13 134168 99899 134568
rect 13 134032 99120 134168
rect 880 133888 99120 134032
rect 880 133752 99899 133888
rect 13 133488 99899 133752
rect 13 133208 99120 133488
rect 13 133080 99899 133208
rect 880 132800 99899 133080
rect 13 132672 99899 132800
rect 13 132392 99120 132672
rect 13 132264 99899 132392
rect 880 131984 99899 132264
rect 13 131856 99899 131984
rect 13 131576 99120 131856
rect 13 131448 99899 131576
rect 880 131168 99899 131448
rect 13 131040 99899 131168
rect 13 130760 99120 131040
rect 13 130632 99899 130760
rect 880 130352 99899 130632
rect 13 130224 99899 130352
rect 13 129944 99120 130224
rect 13 129816 99899 129944
rect 880 129536 99899 129816
rect 13 129408 99899 129536
rect 13 129128 99120 129408
rect 13 129000 99899 129128
rect 880 128728 99899 129000
rect 880 128720 99120 128728
rect 13 128448 99120 128720
rect 13 128184 99899 128448
rect 880 127912 99899 128184
rect 880 127904 99120 127912
rect 13 127632 99120 127904
rect 13 127368 99899 127632
rect 880 127096 99899 127368
rect 880 127088 99120 127096
rect 13 126816 99120 127088
rect 13 126552 99899 126816
rect 880 126280 99899 126552
rect 880 126272 99120 126280
rect 13 126000 99120 126272
rect 13 125736 99899 126000
rect 880 125464 99899 125736
rect 880 125456 99120 125464
rect 13 125184 99120 125456
rect 13 124784 99899 125184
rect 880 124504 99120 124784
rect 13 123968 99899 124504
rect 880 123688 99120 123968
rect 13 123152 99899 123688
rect 880 122872 99120 123152
rect 13 122336 99899 122872
rect 880 122056 99120 122336
rect 13 121520 99899 122056
rect 880 121240 99120 121520
rect 13 120704 99899 121240
rect 880 120424 99120 120704
rect 13 120024 99899 120424
rect 13 119888 99120 120024
rect 880 119744 99120 119888
rect 880 119608 99899 119744
rect 13 119208 99899 119608
rect 13 119072 99120 119208
rect 880 118928 99120 119072
rect 880 118792 99899 118928
rect 13 118392 99899 118792
rect 13 118256 99120 118392
rect 880 118112 99120 118256
rect 880 117976 99899 118112
rect 13 117576 99899 117976
rect 13 117440 99120 117576
rect 880 117296 99120 117440
rect 880 117160 99899 117296
rect 13 116760 99899 117160
rect 13 116624 99120 116760
rect 880 116480 99120 116624
rect 880 116344 99899 116480
rect 13 115944 99899 116344
rect 13 115672 99120 115944
rect 880 115664 99120 115672
rect 880 115392 99899 115664
rect 13 115264 99899 115392
rect 13 114984 99120 115264
rect 13 114856 99899 114984
rect 880 114576 99899 114856
rect 13 114448 99899 114576
rect 13 114168 99120 114448
rect 13 114040 99899 114168
rect 880 113760 99899 114040
rect 13 113632 99899 113760
rect 13 113352 99120 113632
rect 13 113224 99899 113352
rect 880 112944 99899 113224
rect 13 112816 99899 112944
rect 13 112536 99120 112816
rect 13 112408 99899 112536
rect 880 112128 99899 112408
rect 13 112000 99899 112128
rect 13 111720 99120 112000
rect 13 111592 99899 111720
rect 880 111320 99899 111592
rect 880 111312 99120 111320
rect 13 111040 99120 111312
rect 13 110776 99899 111040
rect 880 110504 99899 110776
rect 880 110496 99120 110504
rect 13 110224 99120 110496
rect 13 109960 99899 110224
rect 880 109688 99899 109960
rect 880 109680 99120 109688
rect 13 109408 99120 109680
rect 13 109144 99899 109408
rect 880 108872 99899 109144
rect 880 108864 99120 108872
rect 13 108592 99120 108864
rect 13 108328 99899 108592
rect 880 108056 99899 108328
rect 880 108048 99120 108056
rect 13 107776 99120 108048
rect 13 107512 99899 107776
rect 880 107240 99899 107512
rect 880 107232 99120 107240
rect 13 106960 99120 107232
rect 13 106560 99899 106960
rect 880 106280 99120 106560
rect 13 105744 99899 106280
rect 880 105464 99120 105744
rect 13 104928 99899 105464
rect 880 104648 99120 104928
rect 13 104112 99899 104648
rect 880 103832 99120 104112
rect 13 103296 99899 103832
rect 880 103016 99120 103296
rect 13 102616 99899 103016
rect 13 102480 99120 102616
rect 880 102336 99120 102480
rect 880 102200 99899 102336
rect 13 101800 99899 102200
rect 13 101664 99120 101800
rect 880 101520 99120 101664
rect 880 101384 99899 101520
rect 13 100984 99899 101384
rect 13 100848 99120 100984
rect 880 100704 99120 100848
rect 880 100568 99899 100704
rect 13 100168 99899 100568
rect 13 100032 99120 100168
rect 880 99888 99120 100032
rect 880 99752 99899 99888
rect 13 99352 99899 99752
rect 13 99216 99120 99352
rect 880 99072 99120 99216
rect 880 98936 99899 99072
rect 13 98536 99899 98936
rect 13 98400 99120 98536
rect 880 98256 99120 98400
rect 880 98120 99899 98256
rect 13 97856 99899 98120
rect 13 97576 99120 97856
rect 13 97448 99899 97576
rect 880 97168 99899 97448
rect 13 97040 99899 97168
rect 13 96760 99120 97040
rect 13 96632 99899 96760
rect 880 96352 99899 96632
rect 13 96224 99899 96352
rect 13 95944 99120 96224
rect 13 95816 99899 95944
rect 880 95536 99899 95816
rect 13 95408 99899 95536
rect 13 95128 99120 95408
rect 13 95000 99899 95128
rect 880 94720 99899 95000
rect 13 94592 99899 94720
rect 13 94312 99120 94592
rect 13 94184 99899 94312
rect 880 93904 99899 94184
rect 13 93776 99899 93904
rect 13 93496 99120 93776
rect 13 93368 99899 93496
rect 880 93096 99899 93368
rect 880 93088 99120 93096
rect 13 92816 99120 93088
rect 13 92552 99899 92816
rect 880 92280 99899 92552
rect 880 92272 99120 92280
rect 13 92000 99120 92272
rect 13 91736 99899 92000
rect 880 91464 99899 91736
rect 880 91456 99120 91464
rect 13 91184 99120 91456
rect 13 90920 99899 91184
rect 880 90648 99899 90920
rect 880 90640 99120 90648
rect 13 90368 99120 90640
rect 13 90104 99899 90368
rect 880 89832 99899 90104
rect 880 89824 99120 89832
rect 13 89552 99120 89824
rect 13 89152 99899 89552
rect 880 88872 99120 89152
rect 13 88336 99899 88872
rect 880 88056 99120 88336
rect 13 87520 99899 88056
rect 880 87240 99120 87520
rect 13 86704 99899 87240
rect 880 86424 99120 86704
rect 13 85888 99899 86424
rect 880 85608 99120 85888
rect 13 85072 99899 85608
rect 880 84792 99120 85072
rect 13 84392 99899 84792
rect 13 84256 99120 84392
rect 880 84112 99120 84256
rect 880 83976 99899 84112
rect 13 83576 99899 83976
rect 13 83440 99120 83576
rect 880 83296 99120 83440
rect 880 83160 99899 83296
rect 13 82760 99899 83160
rect 13 82624 99120 82760
rect 880 82480 99120 82624
rect 880 82344 99899 82480
rect 13 81944 99899 82344
rect 13 81808 99120 81944
rect 880 81664 99120 81808
rect 880 81528 99899 81664
rect 13 81128 99899 81528
rect 13 80992 99120 81128
rect 880 80848 99120 80992
rect 880 80712 99899 80848
rect 13 80448 99899 80712
rect 13 80168 99120 80448
rect 13 80040 99899 80168
rect 880 79760 99899 80040
rect 13 79632 99899 79760
rect 13 79352 99120 79632
rect 13 79224 99899 79352
rect 880 78944 99899 79224
rect 13 78816 99899 78944
rect 13 78536 99120 78816
rect 13 78408 99899 78536
rect 880 78128 99899 78408
rect 13 78000 99899 78128
rect 13 77720 99120 78000
rect 13 77592 99899 77720
rect 880 77312 99899 77592
rect 13 77184 99899 77312
rect 13 76904 99120 77184
rect 13 76776 99899 76904
rect 880 76496 99899 76776
rect 13 76368 99899 76496
rect 13 76088 99120 76368
rect 13 75960 99899 76088
rect 880 75688 99899 75960
rect 880 75680 99120 75688
rect 13 75408 99120 75680
rect 13 75144 99899 75408
rect 880 74872 99899 75144
rect 880 74864 99120 74872
rect 13 74592 99120 74864
rect 13 74328 99899 74592
rect 880 74056 99899 74328
rect 880 74048 99120 74056
rect 13 73776 99120 74048
rect 13 73512 99899 73776
rect 880 73240 99899 73512
rect 880 73232 99120 73240
rect 13 72960 99120 73232
rect 13 72696 99899 72960
rect 880 72424 99899 72696
rect 880 72416 99120 72424
rect 13 72144 99120 72416
rect 13 71880 99899 72144
rect 880 71608 99899 71880
rect 880 71600 99120 71608
rect 13 71328 99120 71600
rect 13 70928 99899 71328
rect 880 70648 99120 70928
rect 13 70112 99899 70648
rect 880 69832 99120 70112
rect 13 69296 99899 69832
rect 880 69016 99120 69296
rect 13 68480 99899 69016
rect 880 68200 99120 68480
rect 13 67664 99899 68200
rect 880 67384 99120 67664
rect 13 66984 99899 67384
rect 13 66848 99120 66984
rect 880 66704 99120 66848
rect 880 66568 99899 66704
rect 13 66168 99899 66568
rect 13 66032 99120 66168
rect 880 65888 99120 66032
rect 880 65752 99899 65888
rect 13 65352 99899 65752
rect 13 65216 99120 65352
rect 880 65072 99120 65216
rect 880 64936 99899 65072
rect 13 64536 99899 64936
rect 13 64400 99120 64536
rect 880 64256 99120 64400
rect 880 64120 99899 64256
rect 13 63720 99899 64120
rect 13 63584 99120 63720
rect 880 63440 99120 63584
rect 880 63304 99899 63440
rect 13 62904 99899 63304
rect 13 62632 99120 62904
rect 880 62624 99120 62632
rect 880 62352 99899 62624
rect 13 62224 99899 62352
rect 13 61944 99120 62224
rect 13 61816 99899 61944
rect 880 61536 99899 61816
rect 13 61408 99899 61536
rect 13 61128 99120 61408
rect 13 61000 99899 61128
rect 880 60720 99899 61000
rect 13 60592 99899 60720
rect 13 60312 99120 60592
rect 13 60184 99899 60312
rect 880 59904 99899 60184
rect 13 59776 99899 59904
rect 13 59496 99120 59776
rect 13 59368 99899 59496
rect 880 59088 99899 59368
rect 13 58960 99899 59088
rect 13 58680 99120 58960
rect 13 58552 99899 58680
rect 880 58272 99899 58552
rect 13 58144 99899 58272
rect 13 57864 99120 58144
rect 13 57736 99899 57864
rect 880 57464 99899 57736
rect 880 57456 99120 57464
rect 13 57184 99120 57456
rect 13 56920 99899 57184
rect 880 56648 99899 56920
rect 880 56640 99120 56648
rect 13 56368 99120 56640
rect 13 56104 99899 56368
rect 880 55832 99899 56104
rect 880 55824 99120 55832
rect 13 55552 99120 55824
rect 13 55288 99899 55552
rect 880 55016 99899 55288
rect 880 55008 99120 55016
rect 13 54736 99120 55008
rect 13 54472 99899 54736
rect 880 54200 99899 54472
rect 880 54192 99120 54200
rect 13 53920 99120 54192
rect 13 53520 99899 53920
rect 880 53240 99120 53520
rect 13 52704 99899 53240
rect 880 52424 99120 52704
rect 13 51888 99899 52424
rect 880 51608 99120 51888
rect 13 51072 99899 51608
rect 880 50792 99120 51072
rect 13 50256 99899 50792
rect 880 49976 99120 50256
rect 13 49440 99899 49976
rect 880 49160 99120 49440
rect 13 48760 99899 49160
rect 13 48624 99120 48760
rect 880 48480 99120 48624
rect 880 48344 99899 48480
rect 13 47944 99899 48344
rect 13 47808 99120 47944
rect 880 47664 99120 47808
rect 880 47528 99899 47664
rect 13 47128 99899 47528
rect 13 46992 99120 47128
rect 880 46848 99120 46992
rect 880 46712 99899 46848
rect 13 46312 99899 46712
rect 13 46176 99120 46312
rect 880 46032 99120 46176
rect 880 45896 99899 46032
rect 13 45496 99899 45896
rect 13 45360 99120 45496
rect 880 45216 99120 45360
rect 880 45080 99899 45216
rect 13 44816 99899 45080
rect 13 44536 99120 44816
rect 13 44408 99899 44536
rect 880 44128 99899 44408
rect 13 44000 99899 44128
rect 13 43720 99120 44000
rect 13 43592 99899 43720
rect 880 43312 99899 43592
rect 13 43184 99899 43312
rect 13 42904 99120 43184
rect 13 42776 99899 42904
rect 880 42496 99899 42776
rect 13 42368 99899 42496
rect 13 42088 99120 42368
rect 13 41960 99899 42088
rect 880 41680 99899 41960
rect 13 41552 99899 41680
rect 13 41272 99120 41552
rect 13 41144 99899 41272
rect 880 40864 99899 41144
rect 13 40736 99899 40864
rect 13 40456 99120 40736
rect 13 40328 99899 40456
rect 880 40056 99899 40328
rect 880 40048 99120 40056
rect 13 39776 99120 40048
rect 13 39512 99899 39776
rect 880 39240 99899 39512
rect 880 39232 99120 39240
rect 13 38960 99120 39232
rect 13 38696 99899 38960
rect 880 38424 99899 38696
rect 880 38416 99120 38424
rect 13 38144 99120 38416
rect 13 37880 99899 38144
rect 880 37608 99899 37880
rect 880 37600 99120 37608
rect 13 37328 99120 37600
rect 13 37064 99899 37328
rect 880 36792 99899 37064
rect 880 36784 99120 36792
rect 13 36512 99120 36784
rect 13 36248 99899 36512
rect 880 35976 99899 36248
rect 880 35968 99120 35976
rect 13 35696 99120 35968
rect 13 35296 99899 35696
rect 880 35016 99120 35296
rect 13 34480 99899 35016
rect 880 34200 99120 34480
rect 13 33664 99899 34200
rect 880 33384 99120 33664
rect 13 32848 99899 33384
rect 880 32568 99120 32848
rect 13 32032 99899 32568
rect 880 31752 99120 32032
rect 13 31352 99899 31752
rect 13 31216 99120 31352
rect 880 31072 99120 31216
rect 880 30936 99899 31072
rect 13 30536 99899 30936
rect 13 30400 99120 30536
rect 880 30256 99120 30400
rect 880 30120 99899 30256
rect 13 29720 99899 30120
rect 13 29584 99120 29720
rect 880 29440 99120 29584
rect 880 29304 99899 29440
rect 13 28904 99899 29304
rect 13 28768 99120 28904
rect 880 28624 99120 28768
rect 880 28488 99899 28624
rect 13 28088 99899 28488
rect 13 27952 99120 28088
rect 880 27808 99120 27952
rect 880 27672 99899 27808
rect 13 27272 99899 27672
rect 13 27000 99120 27272
rect 880 26992 99120 27000
rect 880 26720 99899 26992
rect 13 26592 99899 26720
rect 13 26312 99120 26592
rect 13 26184 99899 26312
rect 880 25904 99899 26184
rect 13 25776 99899 25904
rect 13 25496 99120 25776
rect 13 25368 99899 25496
rect 880 25088 99899 25368
rect 13 24960 99899 25088
rect 13 24680 99120 24960
rect 13 24552 99899 24680
rect 880 24272 99899 24552
rect 13 24144 99899 24272
rect 13 23864 99120 24144
rect 13 23736 99899 23864
rect 880 23456 99899 23736
rect 13 23328 99899 23456
rect 13 23048 99120 23328
rect 13 22920 99899 23048
rect 880 22648 99899 22920
rect 880 22640 99120 22648
rect 13 22368 99120 22640
rect 13 22104 99899 22368
rect 880 21832 99899 22104
rect 880 21824 99120 21832
rect 13 21552 99120 21824
rect 13 21288 99899 21552
rect 880 21016 99899 21288
rect 880 21008 99120 21016
rect 13 20736 99120 21008
rect 13 20472 99899 20736
rect 880 20200 99899 20472
rect 880 20192 99120 20200
rect 13 19920 99120 20192
rect 13 19656 99899 19920
rect 880 19384 99899 19656
rect 880 19376 99120 19384
rect 13 19104 99120 19376
rect 13 18840 99899 19104
rect 880 18568 99899 18840
rect 880 18560 99120 18568
rect 13 18288 99120 18560
rect 13 17888 99899 18288
rect 880 17608 99120 17888
rect 13 17072 99899 17608
rect 880 16792 99120 17072
rect 13 16256 99899 16792
rect 880 15976 99120 16256
rect 13 15440 99899 15976
rect 880 15160 99120 15440
rect 13 14624 99899 15160
rect 880 14344 99120 14624
rect 13 13808 99899 14344
rect 880 13528 99120 13808
rect 13 13128 99899 13528
rect 13 12992 99120 13128
rect 880 12848 99120 12992
rect 880 12712 99899 12848
rect 13 12312 99899 12712
rect 13 12176 99120 12312
rect 880 12032 99120 12176
rect 880 11896 99899 12032
rect 13 11496 99899 11896
rect 13 11360 99120 11496
rect 880 11216 99120 11360
rect 880 11080 99899 11216
rect 13 10680 99899 11080
rect 13 10544 99120 10680
rect 880 10400 99120 10544
rect 880 10264 99899 10400
rect 13 9864 99899 10264
rect 13 9728 99120 9864
rect 880 9584 99120 9728
rect 880 9448 99899 9584
rect 13 9184 99899 9448
rect 13 8904 99120 9184
rect 13 8776 99899 8904
rect 880 8496 99899 8776
rect 13 8368 99899 8496
rect 13 8088 99120 8368
rect 13 7960 99899 8088
rect 880 7680 99899 7960
rect 13 7552 99899 7680
rect 13 7272 99120 7552
rect 13 7144 99899 7272
rect 880 6864 99899 7144
rect 13 6736 99899 6864
rect 13 6456 99120 6736
rect 13 6328 99899 6456
rect 880 6048 99899 6328
rect 13 5920 99899 6048
rect 13 5640 99120 5920
rect 13 5512 99899 5640
rect 880 5232 99899 5512
rect 13 5104 99899 5232
rect 13 4824 99120 5104
rect 13 4696 99899 4824
rect 880 4424 99899 4696
rect 880 4416 99120 4424
rect 13 4144 99120 4416
rect 13 3880 99899 4144
rect 880 3608 99899 3880
rect 880 3600 99120 3608
rect 13 3328 99120 3600
rect 13 3064 99899 3328
rect 880 2792 99899 3064
rect 880 2784 99120 2792
rect 13 2512 99120 2784
rect 13 2248 99899 2512
rect 880 1976 99899 2248
rect 880 1968 99120 1976
rect 13 1696 99120 1968
rect 13 1432 99899 1696
rect 880 1160 99899 1432
rect 880 1152 99120 1160
rect 13 880 99120 1152
rect 13 616 99899 880
rect 880 480 99899 616
rect 880 336 99120 480
rect 13 307 99120 336
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
<< obsm4 >>
rect 2083 4795 4128 155141
rect 4608 4795 19488 155141
rect 19968 4795 34848 155141
rect 35328 4795 50208 155141
rect 50688 4795 65568 155141
rect 66048 4795 80928 155141
rect 81408 4795 96288 155141
rect 96768 4795 99117 155141
<< labels >>
rlabel metal3 s 0 10344 800 10464 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 103912 800 104032 6 addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 clk0
port 19 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 clk1
port 20 nsew signal output
rlabel metal2 s 1214 159200 1270 160000 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 3698 159200 3754 160000 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 6274 159200 6330 160000 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 8850 159200 8906 160000 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 11426 159200 11482 160000 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 14002 159200 14058 160000 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 16578 159200 16634 160000 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 19154 159200 19210 160000 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 99200 1776 100000 1896 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 99200 6536 100000 6656 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 99200 33464 100000 33584 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 99200 35776 100000 35896 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 99200 38224 100000 38344 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 99200 40536 100000 40656 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 99200 42984 100000 43104 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 99200 45296 100000 45416 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 99200 47744 100000 47864 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 99200 50056 100000 50176 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 99200 52504 100000 52624 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 99200 54816 100000 54936 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 99200 9664 100000 9784 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 99200 57264 100000 57384 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 99200 59576 100000 59696 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 99200 62024 100000 62144 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 99200 64336 100000 64456 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 99200 66784 100000 66904 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 99200 69096 100000 69216 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 99200 71408 100000 71528 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 99200 73856 100000 73976 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 99200 12928 100000 13048 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 99200 16056 100000 16176 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 99200 19184 100000 19304 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 99200 21632 100000 21752 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 99200 23944 100000 24064 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 99200 26392 100000 26512 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 99200 28704 100000 28824 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 99200 31152 100000 31272 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 99200 2592 100000 2712 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 99200 7352 100000 7472 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 99200 34280 100000 34400 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 99200 36592 100000 36712 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 99200 39040 100000 39160 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 99200 41352 100000 41472 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 99200 43800 100000 43920 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 99200 46112 100000 46232 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 99200 48560 100000 48680 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 99200 50872 100000 50992 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 99200 53320 100000 53440 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 99200 55632 100000 55752 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 99200 10480 100000 10600 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 99200 57944 100000 58064 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 99200 60392 100000 60512 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 99200 62704 100000 62824 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 99200 65152 100000 65272 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 99200 67464 100000 67584 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 99200 69912 100000 70032 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 99200 72224 100000 72344 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 99200 74672 100000 74792 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 99200 76168 100000 76288 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 99200 77800 100000 77920 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 99200 13608 100000 13728 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 99200 79432 100000 79552 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 99200 80928 100000 81048 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 99200 16872 100000 16992 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 99200 20000 100000 20120 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 99200 22448 100000 22568 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 99200 24760 100000 24880 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 99200 27072 100000 27192 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 99200 29520 100000 29640 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 99200 31832 100000 31952 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 99200 8168 100000 8288 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 99200 35096 100000 35216 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 99200 37408 100000 37528 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 99200 39856 100000 39976 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 99200 42168 100000 42288 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 99200 44616 100000 44736 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 99200 46928 100000 47048 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 99200 49240 100000 49360 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 99200 51688 100000 51808 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 99200 54000 100000 54120 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 99200 56448 100000 56568 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 99200 11296 100000 11416 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 99200 58760 100000 58880 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 99200 61208 100000 61328 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 99200 63520 100000 63640 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 99200 65968 100000 66088 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 99200 68280 100000 68400 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 99200 70728 100000 70848 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 99200 73040 100000 73160 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 99200 75488 100000 75608 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 99200 76984 100000 77104 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 99200 78616 100000 78736 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 99200 14424 100000 14544 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 99200 80248 100000 80368 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 99200 81744 100000 81864 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 99200 17688 100000 17808 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 99200 20816 100000 20936 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 99200 23128 100000 23248 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 99200 25576 100000 25696 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 99200 27888 100000 28008 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 99200 30336 100000 30456 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 99200 32648 100000 32768 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 99200 3408 100000 3528 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 99200 8984 100000 9104 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 99200 12112 100000 12232 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 99200 15240 100000 15360 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 99200 18368 100000 18488 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 99200 4224 100000 4344 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 99200 4904 100000 5024 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 99200 5720 100000 5840 6 core_wb_we_o
port 130 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 csb0[0]
port 131 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 csb0[1]
port 132 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 csb1[1]
port 134 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 din0[0]
port 135 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 din0[10]
port 136 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 din0[11]
port 137 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 din0[12]
port 138 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 din0[13]
port 139 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 din0[14]
port 140 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 din0[15]
port 141 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 din0[16]
port 142 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 din0[17]
port 143 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 din0[18]
port 144 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 din0[19]
port 145 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 din0[1]
port 146 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 din0[20]
port 147 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 din0[21]
port 148 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 din0[22]
port 149 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 din0[23]
port 150 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 din0[24]
port 151 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 din0[25]
port 152 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 din0[26]
port 153 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 din0[27]
port 154 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 din0[28]
port 155 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 din0[29]
port 156 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 din0[2]
port 157 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 din0[30]
port 158 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 din0[31]
port 159 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 din0[3]
port 160 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 din0[4]
port 161 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 din0[5]
port 162 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 din0[6]
port 163 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 din0[7]
port 164 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 din0[8]
port 165 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 din0[9]
port 166 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 dout0[0]
port 167 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 dout0[10]
port 168 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 dout0[11]
port 169 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 dout0[12]
port 170 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 dout0[13]
port 171 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 dout0[14]
port 172 nsew signal input
rlabel metal3 s 0 56720 800 56840 6 dout0[15]
port 173 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 dout0[16]
port 174 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 dout0[17]
port 175 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 dout0[18]
port 176 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 dout0[19]
port 177 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 dout0[1]
port 178 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 dout0[20]
port 179 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 dout0[21]
port 180 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 dout0[22]
port 181 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 dout0[23]
port 182 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 dout0[24]
port 183 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 dout0[25]
port 184 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 dout0[26]
port 185 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 dout0[27]
port 186 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 dout0[28]
port 187 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 dout0[29]
port 188 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 dout0[2]
port 189 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 dout0[30]
port 190 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 dout0[31]
port 191 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 dout0[32]
port 192 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 dout0[33]
port 193 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 dout0[34]
port 194 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 dout0[35]
port 195 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 dout0[36]
port 196 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 dout0[37]
port 197 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 dout0[38]
port 198 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 dout0[39]
port 199 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 dout0[3]
port 200 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 dout0[40]
port 201 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 dout0[41]
port 202 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 dout0[42]
port 203 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 dout0[43]
port 204 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 dout0[44]
port 205 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 dout0[45]
port 206 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 dout0[46]
port 207 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 dout0[47]
port 208 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 dout0[48]
port 209 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 dout0[49]
port 210 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 dout0[4]
port 211 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 dout0[50]
port 212 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 dout0[51]
port 213 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 dout0[52]
port 214 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 dout0[53]
port 215 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 dout0[54]
port 216 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 dout0[55]
port 217 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 dout0[56]
port 218 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 dout0[57]
port 219 nsew signal input
rlabel metal3 s 0 92352 800 92472 6 dout0[58]
port 220 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 dout0[59]
port 221 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 dout0[5]
port 222 nsew signal input
rlabel metal3 s 0 93984 800 94104 6 dout0[60]
port 223 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 dout0[61]
port 224 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 dout0[62]
port 225 nsew signal input
rlabel metal3 s 0 96432 800 96552 6 dout0[63]
port 226 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 dout0[6]
port 227 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 dout0[7]
port 228 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 dout0[8]
port 229 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 dout0[9]
port 230 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 dout1[0]
port 231 nsew signal input
rlabel metal3 s 0 115472 800 115592 6 dout1[10]
port 232 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 dout1[11]
port 233 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 dout1[12]
port 234 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 dout1[13]
port 235 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 dout1[14]
port 236 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 dout1[15]
port 237 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 dout1[16]
port 238 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 dout1[17]
port 239 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 dout1[18]
port 240 nsew signal input
rlabel metal3 s 0 122952 800 123072 6 dout1[19]
port 241 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 dout1[1]
port 242 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 dout1[20]
port 243 nsew signal input
rlabel metal3 s 0 124584 800 124704 6 dout1[21]
port 244 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 dout1[22]
port 245 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 dout1[23]
port 246 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 dout1[24]
port 247 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 dout1[25]
port 248 nsew signal input
rlabel metal3 s 0 128800 800 128920 6 dout1[26]
port 249 nsew signal input
rlabel metal3 s 0 129616 800 129736 6 dout1[27]
port 250 nsew signal input
rlabel metal3 s 0 130432 800 130552 6 dout1[28]
port 251 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 dout1[29]
port 252 nsew signal input
rlabel metal3 s 0 108944 800 109064 6 dout1[2]
port 253 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 dout1[30]
port 254 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 dout1[31]
port 255 nsew signal input
rlabel metal3 s 0 133832 800 133952 6 dout1[32]
port 256 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 dout1[33]
port 257 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 dout1[34]
port 258 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 dout1[35]
port 259 nsew signal input
rlabel metal3 s 0 137096 800 137216 6 dout1[36]
port 260 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 dout1[37]
port 261 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 dout1[38]
port 262 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 dout1[39]
port 263 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 dout1[3]
port 264 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 dout1[40]
port 265 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 dout1[41]
port 266 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 dout1[42]
port 267 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 dout1[43]
port 268 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 dout1[44]
port 269 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 dout1[45]
port 270 nsew signal input
rlabel metal3 s 0 145392 800 145512 6 dout1[46]
port 271 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 dout1[47]
port 272 nsew signal input
rlabel metal3 s 0 147024 800 147144 6 dout1[48]
port 273 nsew signal input
rlabel metal3 s 0 147840 800 147960 6 dout1[49]
port 274 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 dout1[4]
port 275 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 dout1[50]
port 276 nsew signal input
rlabel metal3 s 0 149472 800 149592 6 dout1[51]
port 277 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 dout1[52]
port 278 nsew signal input
rlabel metal3 s 0 151104 800 151224 6 dout1[53]
port 279 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 dout1[54]
port 280 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 dout1[55]
port 281 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 dout1[56]
port 282 nsew signal input
rlabel metal3 s 0 154504 800 154624 6 dout1[57]
port 283 nsew signal input
rlabel metal3 s 0 155320 800 155440 6 dout1[58]
port 284 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 dout1[59]
port 285 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 dout1[5]
port 286 nsew signal input
rlabel metal3 s 0 156952 800 157072 6 dout1[60]
port 287 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 dout1[61]
port 288 nsew signal input
rlabel metal3 s 0 158584 800 158704 6 dout1[62]
port 289 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 dout1[63]
port 290 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 dout1[6]
port 291 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 dout1[7]
port 292 nsew signal input
rlabel metal3 s 0 113840 800 113960 6 dout1[8]
port 293 nsew signal input
rlabel metal3 s 0 114656 800 114776 6 dout1[9]
port 294 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 irq[0]
port 295 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 irq[10]
port 296 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 irq[11]
port 297 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 irq[12]
port 298 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 irq[13]
port 299 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 irq[14]
port 300 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 irq[15]
port 301 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 irq[1]
port 302 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 irq[2]
port 303 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 irq[3]
port 304 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 irq[4]
port 305 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 irq[5]
port 306 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 irq[6]
port 307 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 irq[7]
port 308 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 irq[8]
port 309 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 irq[9]
port 310 nsew signal input
rlabel metal3 s 0 416 800 536 6 jtag_tck
port 311 nsew signal input
rlabel metal3 s 0 1232 800 1352 6 jtag_tdi
port 312 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 jtag_tdo
port 313 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 jtag_tms
port 314 nsew signal input
rlabel metal3 s 99200 82560 100000 82680 6 localMemory_wb_ack_o
port 315 nsew signal output
rlabel metal3 s 99200 87320 100000 87440 6 localMemory_wb_adr_i[0]
port 316 nsew signal input
rlabel metal3 s 99200 114248 100000 114368 6 localMemory_wb_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 99200 116560 100000 116680 6 localMemory_wb_adr_i[11]
port 318 nsew signal input
rlabel metal3 s 99200 119008 100000 119128 6 localMemory_wb_adr_i[12]
port 319 nsew signal input
rlabel metal3 s 99200 121320 100000 121440 6 localMemory_wb_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 99200 123768 100000 123888 6 localMemory_wb_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 99200 126080 100000 126200 6 localMemory_wb_adr_i[15]
port 322 nsew signal input
rlabel metal3 s 99200 128528 100000 128648 6 localMemory_wb_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 99200 130840 100000 130960 6 localMemory_wb_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 99200 133288 100000 133408 6 localMemory_wb_adr_i[18]
port 325 nsew signal input
rlabel metal3 s 99200 135600 100000 135720 6 localMemory_wb_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 99200 90448 100000 90568 6 localMemory_wb_adr_i[1]
port 327 nsew signal input
rlabel metal3 s 99200 137912 100000 138032 6 localMemory_wb_adr_i[20]
port 328 nsew signal input
rlabel metal3 s 99200 140360 100000 140480 6 localMemory_wb_adr_i[21]
port 329 nsew signal input
rlabel metal3 s 99200 142672 100000 142792 6 localMemory_wb_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 99200 145120 100000 145240 6 localMemory_wb_adr_i[23]
port 331 nsew signal input
rlabel metal3 s 99200 93576 100000 93696 6 localMemory_wb_adr_i[2]
port 332 nsew signal input
rlabel metal3 s 99200 96840 100000 96960 6 localMemory_wb_adr_i[3]
port 333 nsew signal input
rlabel metal3 s 99200 99968 100000 100088 6 localMemory_wb_adr_i[4]
port 334 nsew signal input
rlabel metal3 s 99200 102416 100000 102536 6 localMemory_wb_adr_i[5]
port 335 nsew signal input
rlabel metal3 s 99200 104728 100000 104848 6 localMemory_wb_adr_i[6]
port 336 nsew signal input
rlabel metal3 s 99200 107040 100000 107160 6 localMemory_wb_adr_i[7]
port 337 nsew signal input
rlabel metal3 s 99200 109488 100000 109608 6 localMemory_wb_adr_i[8]
port 338 nsew signal input
rlabel metal3 s 99200 111800 100000 111920 6 localMemory_wb_adr_i[9]
port 339 nsew signal input
rlabel metal3 s 99200 83376 100000 83496 6 localMemory_wb_cyc_i
port 340 nsew signal input
rlabel metal3 s 99200 88136 100000 88256 6 localMemory_wb_data_i[0]
port 341 nsew signal input
rlabel metal3 s 99200 115064 100000 115184 6 localMemory_wb_data_i[10]
port 342 nsew signal input
rlabel metal3 s 99200 117376 100000 117496 6 localMemory_wb_data_i[11]
port 343 nsew signal input
rlabel metal3 s 99200 119824 100000 119944 6 localMemory_wb_data_i[12]
port 344 nsew signal input
rlabel metal3 s 99200 122136 100000 122256 6 localMemory_wb_data_i[13]
port 345 nsew signal input
rlabel metal3 s 99200 124584 100000 124704 6 localMemory_wb_data_i[14]
port 346 nsew signal input
rlabel metal3 s 99200 126896 100000 127016 6 localMemory_wb_data_i[15]
port 347 nsew signal input
rlabel metal3 s 99200 129208 100000 129328 6 localMemory_wb_data_i[16]
port 348 nsew signal input
rlabel metal3 s 99200 131656 100000 131776 6 localMemory_wb_data_i[17]
port 349 nsew signal input
rlabel metal3 s 99200 133968 100000 134088 6 localMemory_wb_data_i[18]
port 350 nsew signal input
rlabel metal3 s 99200 136416 100000 136536 6 localMemory_wb_data_i[19]
port 351 nsew signal input
rlabel metal3 s 99200 91264 100000 91384 6 localMemory_wb_data_i[1]
port 352 nsew signal input
rlabel metal3 s 99200 138728 100000 138848 6 localMemory_wb_data_i[20]
port 353 nsew signal input
rlabel metal3 s 99200 141176 100000 141296 6 localMemory_wb_data_i[21]
port 354 nsew signal input
rlabel metal3 s 99200 143488 100000 143608 6 localMemory_wb_data_i[22]
port 355 nsew signal input
rlabel metal3 s 99200 145936 100000 146056 6 localMemory_wb_data_i[23]
port 356 nsew signal input
rlabel metal3 s 99200 147432 100000 147552 6 localMemory_wb_data_i[24]
port 357 nsew signal input
rlabel metal3 s 99200 149064 100000 149184 6 localMemory_wb_data_i[25]
port 358 nsew signal input
rlabel metal3 s 99200 150696 100000 150816 6 localMemory_wb_data_i[26]
port 359 nsew signal input
rlabel metal3 s 99200 152192 100000 152312 6 localMemory_wb_data_i[27]
port 360 nsew signal input
rlabel metal3 s 99200 153824 100000 153944 6 localMemory_wb_data_i[28]
port 361 nsew signal input
rlabel metal3 s 99200 155456 100000 155576 6 localMemory_wb_data_i[29]
port 362 nsew signal input
rlabel metal3 s 99200 94392 100000 94512 6 localMemory_wb_data_i[2]
port 363 nsew signal input
rlabel metal3 s 99200 156952 100000 157072 6 localMemory_wb_data_i[30]
port 364 nsew signal input
rlabel metal3 s 99200 158584 100000 158704 6 localMemory_wb_data_i[31]
port 365 nsew signal input
rlabel metal3 s 99200 97656 100000 97776 6 localMemory_wb_data_i[3]
port 366 nsew signal input
rlabel metal3 s 99200 100784 100000 100904 6 localMemory_wb_data_i[4]
port 367 nsew signal input
rlabel metal3 s 99200 103096 100000 103216 6 localMemory_wb_data_i[5]
port 368 nsew signal input
rlabel metal3 s 99200 105544 100000 105664 6 localMemory_wb_data_i[6]
port 369 nsew signal input
rlabel metal3 s 99200 107856 100000 107976 6 localMemory_wb_data_i[7]
port 370 nsew signal input
rlabel metal3 s 99200 110304 100000 110424 6 localMemory_wb_data_i[8]
port 371 nsew signal input
rlabel metal3 s 99200 112616 100000 112736 6 localMemory_wb_data_i[9]
port 372 nsew signal input
rlabel metal3 s 99200 88952 100000 89072 6 localMemory_wb_data_o[0]
port 373 nsew signal output
rlabel metal3 s 99200 115744 100000 115864 6 localMemory_wb_data_o[10]
port 374 nsew signal output
rlabel metal3 s 99200 118192 100000 118312 6 localMemory_wb_data_o[11]
port 375 nsew signal output
rlabel metal3 s 99200 120504 100000 120624 6 localMemory_wb_data_o[12]
port 376 nsew signal output
rlabel metal3 s 99200 122952 100000 123072 6 localMemory_wb_data_o[13]
port 377 nsew signal output
rlabel metal3 s 99200 125264 100000 125384 6 localMemory_wb_data_o[14]
port 378 nsew signal output
rlabel metal3 s 99200 127712 100000 127832 6 localMemory_wb_data_o[15]
port 379 nsew signal output
rlabel metal3 s 99200 130024 100000 130144 6 localMemory_wb_data_o[16]
port 380 nsew signal output
rlabel metal3 s 99200 132472 100000 132592 6 localMemory_wb_data_o[17]
port 381 nsew signal output
rlabel metal3 s 99200 134784 100000 134904 6 localMemory_wb_data_o[18]
port 382 nsew signal output
rlabel metal3 s 99200 137232 100000 137352 6 localMemory_wb_data_o[19]
port 383 nsew signal output
rlabel metal3 s 99200 92080 100000 92200 6 localMemory_wb_data_o[1]
port 384 nsew signal output
rlabel metal3 s 99200 139544 100000 139664 6 localMemory_wb_data_o[20]
port 385 nsew signal output
rlabel metal3 s 99200 141992 100000 142112 6 localMemory_wb_data_o[21]
port 386 nsew signal output
rlabel metal3 s 99200 144304 100000 144424 6 localMemory_wb_data_o[22]
port 387 nsew signal output
rlabel metal3 s 99200 146752 100000 146872 6 localMemory_wb_data_o[23]
port 388 nsew signal output
rlabel metal3 s 99200 148248 100000 148368 6 localMemory_wb_data_o[24]
port 389 nsew signal output
rlabel metal3 s 99200 149880 100000 150000 6 localMemory_wb_data_o[25]
port 390 nsew signal output
rlabel metal3 s 99200 151376 100000 151496 6 localMemory_wb_data_o[26]
port 391 nsew signal output
rlabel metal3 s 99200 153008 100000 153128 6 localMemory_wb_data_o[27]
port 392 nsew signal output
rlabel metal3 s 99200 154640 100000 154760 6 localMemory_wb_data_o[28]
port 393 nsew signal output
rlabel metal3 s 99200 156136 100000 156256 6 localMemory_wb_data_o[29]
port 394 nsew signal output
rlabel metal3 s 99200 95208 100000 95328 6 localMemory_wb_data_o[2]
port 395 nsew signal output
rlabel metal3 s 99200 157768 100000 157888 6 localMemory_wb_data_o[30]
port 396 nsew signal output
rlabel metal3 s 99200 159400 100000 159520 6 localMemory_wb_data_o[31]
port 397 nsew signal output
rlabel metal3 s 99200 98336 100000 98456 6 localMemory_wb_data_o[3]
port 398 nsew signal output
rlabel metal3 s 99200 101600 100000 101720 6 localMemory_wb_data_o[4]
port 399 nsew signal output
rlabel metal3 s 99200 103912 100000 104032 6 localMemory_wb_data_o[5]
port 400 nsew signal output
rlabel metal3 s 99200 106360 100000 106480 6 localMemory_wb_data_o[6]
port 401 nsew signal output
rlabel metal3 s 99200 108672 100000 108792 6 localMemory_wb_data_o[7]
port 402 nsew signal output
rlabel metal3 s 99200 111120 100000 111240 6 localMemory_wb_data_o[8]
port 403 nsew signal output
rlabel metal3 s 99200 113432 100000 113552 6 localMemory_wb_data_o[9]
port 404 nsew signal output
rlabel metal3 s 99200 84192 100000 84312 6 localMemory_wb_error_o
port 405 nsew signal output
rlabel metal3 s 99200 89632 100000 89752 6 localMemory_wb_sel_i[0]
port 406 nsew signal input
rlabel metal3 s 99200 92896 100000 93016 6 localMemory_wb_sel_i[1]
port 407 nsew signal input
rlabel metal3 s 99200 96024 100000 96144 6 localMemory_wb_sel_i[2]
port 408 nsew signal input
rlabel metal3 s 99200 99152 100000 99272 6 localMemory_wb_sel_i[3]
port 409 nsew signal input
rlabel metal3 s 99200 84872 100000 84992 6 localMemory_wb_stall_o
port 410 nsew signal output
rlabel metal3 s 99200 85688 100000 85808 6 localMemory_wb_stb_i
port 411 nsew signal input
rlabel metal3 s 99200 86504 100000 86624 6 localMemory_wb_we_i
port 412 nsew signal input
rlabel metal2 s 21638 159200 21694 160000 6 manufacturerID[0]
port 413 nsew signal input
rlabel metal2 s 47306 159200 47362 160000 6 manufacturerID[10]
port 414 nsew signal input
rlabel metal2 s 24214 159200 24270 160000 6 manufacturerID[1]
port 415 nsew signal input
rlabel metal2 s 26790 159200 26846 160000 6 manufacturerID[2]
port 416 nsew signal input
rlabel metal2 s 29366 159200 29422 160000 6 manufacturerID[3]
port 417 nsew signal input
rlabel metal2 s 31942 159200 31998 160000 6 manufacturerID[4]
port 418 nsew signal input
rlabel metal2 s 34518 159200 34574 160000 6 manufacturerID[5]
port 419 nsew signal input
rlabel metal2 s 37094 159200 37150 160000 6 manufacturerID[6]
port 420 nsew signal input
rlabel metal2 s 39670 159200 39726 160000 6 manufacturerID[7]
port 421 nsew signal input
rlabel metal2 s 42154 159200 42210 160000 6 manufacturerID[8]
port 422 nsew signal input
rlabel metal2 s 44730 159200 44786 160000 6 manufacturerID[9]
port 423 nsew signal input
rlabel metal2 s 49882 159200 49938 160000 6 partID[0]
port 424 nsew signal input
rlabel metal2 s 75550 159200 75606 160000 6 partID[10]
port 425 nsew signal input
rlabel metal2 s 78126 159200 78182 160000 6 partID[11]
port 426 nsew signal input
rlabel metal2 s 80702 159200 80758 160000 6 partID[12]
port 427 nsew signal input
rlabel metal2 s 83186 159200 83242 160000 6 partID[13]
port 428 nsew signal input
rlabel metal2 s 85762 159200 85818 160000 6 partID[14]
port 429 nsew signal input
rlabel metal2 s 88338 159200 88394 160000 6 partID[15]
port 430 nsew signal input
rlabel metal2 s 52458 159200 52514 160000 6 partID[1]
port 431 nsew signal input
rlabel metal2 s 55034 159200 55090 160000 6 partID[2]
port 432 nsew signal input
rlabel metal2 s 57610 159200 57666 160000 6 partID[3]
port 433 nsew signal input
rlabel metal2 s 60186 159200 60242 160000 6 partID[4]
port 434 nsew signal input
rlabel metal2 s 62670 159200 62726 160000 6 partID[5]
port 435 nsew signal input
rlabel metal2 s 65246 159200 65302 160000 6 partID[6]
port 436 nsew signal input
rlabel metal2 s 67822 159200 67878 160000 6 partID[7]
port 437 nsew signal input
rlabel metal2 s 70398 159200 70454 160000 6 partID[8]
port 438 nsew signal input
rlabel metal2 s 72974 159200 73030 160000 6 partID[9]
port 439 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 probe_env[0]
port 440 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 probe_env[1]
port 441 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 probe_jtagInstruction[0]
port 442 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 probe_jtagInstruction[1]
port 443 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 probe_jtagInstruction[2]
port 444 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 probe_jtagInstruction[3]
port 445 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 probe_jtagInstruction[4]
port 446 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 probe_programCounter[0]
port 447 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 probe_programCounter[10]
port 448 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 probe_programCounter[11]
port 449 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 probe_programCounter[12]
port 450 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 probe_programCounter[13]
port 451 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 probe_programCounter[14]
port 452 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 probe_programCounter[15]
port 453 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 probe_programCounter[16]
port 454 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 probe_programCounter[17]
port 455 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 probe_programCounter[18]
port 456 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 probe_programCounter[19]
port 457 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 probe_programCounter[1]
port 458 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 probe_programCounter[20]
port 459 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 probe_programCounter[21]
port 460 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 probe_programCounter[22]
port 461 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 probe_programCounter[23]
port 462 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 probe_programCounter[24]
port 463 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 probe_programCounter[25]
port 464 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 probe_programCounter[26]
port 465 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 probe_programCounter[27]
port 466 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 probe_programCounter[28]
port 467 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 probe_programCounter[29]
port 468 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 probe_programCounter[2]
port 469 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 probe_programCounter[30]
port 470 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 probe_programCounter[31]
port 471 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 probe_programCounter[3]
port 472 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 probe_programCounter[4]
port 473 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 probe_programCounter[5]
port 474 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 probe_programCounter[6]
port 475 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 probe_programCounter[7]
port 476 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 probe_programCounter[8]
port 477 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 probe_programCounter[9]
port 478 nsew signal output
rlabel metal2 s 846 0 902 800 6 probe_state
port 479 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 480 nsew power input
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 480 nsew power input
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 480 nsew power input
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 480 nsew power input
rlabel metal2 s 90914 159200 90970 160000 6 versionID[0]
port 481 nsew signal input
rlabel metal2 s 93490 159200 93546 160000 6 versionID[1]
port 482 nsew signal input
rlabel metal2 s 96066 159200 96122 160000 6 versionID[2]
port 483 nsew signal input
rlabel metal2 s 98642 159200 98698 160000 6 versionID[3]
port 484 nsew signal input
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 485 nsew ground input
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 485 nsew ground input
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 485 nsew ground input
rlabel metal3 s 99200 280 100000 400 6 wb_clk_i
port 486 nsew signal input
rlabel metal3 s 99200 960 100000 1080 6 wb_rst_i
port 487 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 web0
port 488 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 wmask0[0]
port 489 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 wmask0[1]
port 490 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 wmask0[2]
port 491 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 wmask0[3]
port 492 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 52348876
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/finishing/ExperiarCore.magic.gds
string GDS_START 1513918
<< end >>

