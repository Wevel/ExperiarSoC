VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Video
  CLASS BLOCK ;
  FOREIGN Video ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN sram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 496.000 5.430 500.000 ;
    END
  END sram_addr0[0]
  PIN sram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 496.000 17.850 500.000 ;
    END
  END sram_addr0[1]
  PIN sram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 496.000 30.270 500.000 ;
    END
  END sram_addr0[2]
  PIN sram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 496.000 42.690 500.000 ;
    END
  END sram_addr0[3]
  PIN sram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 496.000 55.110 500.000 ;
    END
  END sram_addr0[4]
  PIN sram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 496.000 62.930 500.000 ;
    END
  END sram_addr0[5]
  PIN sram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 496.000 70.750 500.000 ;
    END
  END sram_addr0[6]
  PIN sram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 496.000 78.570 500.000 ;
    END
  END sram_addr0[7]
  PIN sram_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 496.000 86.390 500.000 ;
    END
  END sram_addr0[8]
  PIN sram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 496.000 6.810 500.000 ;
    END
  END sram_addr1[0]
  PIN sram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 496.000 19.230 500.000 ;
    END
  END sram_addr1[1]
  PIN sram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 496.000 31.650 500.000 ;
    END
  END sram_addr1[2]
  PIN sram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 496.000 44.070 500.000 ;
    END
  END sram_addr1[3]
  PIN sram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 496.000 56.490 500.000 ;
    END
  END sram_addr1[4]
  PIN sram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 496.000 64.310 500.000 ;
    END
  END sram_addr1[5]
  PIN sram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 496.000 72.130 500.000 ;
    END
  END sram_addr1[6]
  PIN sram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 496.000 79.950 500.000 ;
    END
  END sram_addr1[7]
  PIN sram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 496.000 87.770 500.000 ;
    END
  END sram_addr1[8]
  PIN sram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 496.000 0.830 500.000 ;
    END
  END sram_clk0
  PIN sram_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 496.000 2.210 500.000 ;
    END
  END sram_clk1
  PIN sram_csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 496.000 8.190 500.000 ;
    END
  END sram_csb0[0]
  PIN sram_csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 496.000 21.070 500.000 ;
    END
  END sram_csb0[1]
  PIN sram_csb0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 496.000 33.490 500.000 ;
    END
  END sram_csb0[2]
  PIN sram_csb0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 496.000 45.910 500.000 ;
    END
  END sram_csb0[3]
  PIN sram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 496.000 10.030 500.000 ;
    END
  END sram_csb1[0]
  PIN sram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 496.000 22.450 500.000 ;
    END
  END sram_csb1[1]
  PIN sram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 496.000 34.870 500.000 ;
    END
  END sram_csb1[2]
  PIN sram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 496.000 47.290 500.000 ;
    END
  END sram_csb1[3]
  PIN sram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 496.000 11.410 500.000 ;
    END
  END sram_din0[0]
  PIN sram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 496.000 98.810 500.000 ;
    END
  END sram_din0[10]
  PIN sram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 496.000 103.410 500.000 ;
    END
  END sram_din0[11]
  PIN sram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 496.000 108.010 500.000 ;
    END
  END sram_din0[12]
  PIN sram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 496.000 112.610 500.000 ;
    END
  END sram_din0[13]
  PIN sram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 496.000 117.210 500.000 ;
    END
  END sram_din0[14]
  PIN sram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 496.000 122.270 500.000 ;
    END
  END sram_din0[15]
  PIN sram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 496.000 126.870 500.000 ;
    END
  END sram_din0[16]
  PIN sram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 496.000 131.470 500.000 ;
    END
  END sram_din0[17]
  PIN sram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 496.000 136.070 500.000 ;
    END
  END sram_din0[18]
  PIN sram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 496.000 140.670 500.000 ;
    END
  END sram_din0[19]
  PIN sram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 496.000 23.830 500.000 ;
    END
  END sram_din0[1]
  PIN sram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 496.000 145.270 500.000 ;
    END
  END sram_din0[20]
  PIN sram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 496.000 150.330 500.000 ;
    END
  END sram_din0[21]
  PIN sram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 496.000 154.930 500.000 ;
    END
  END sram_din0[22]
  PIN sram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 496.000 159.530 500.000 ;
    END
  END sram_din0[23]
  PIN sram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 496.000 164.130 500.000 ;
    END
  END sram_din0[24]
  PIN sram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 496.000 168.730 500.000 ;
    END
  END sram_din0[25]
  PIN sram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 496.000 173.330 500.000 ;
    END
  END sram_din0[26]
  PIN sram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 496.000 178.390 500.000 ;
    END
  END sram_din0[27]
  PIN sram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 496.000 182.990 500.000 ;
    END
  END sram_din0[28]
  PIN sram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 496.000 187.590 500.000 ;
    END
  END sram_din0[29]
  PIN sram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 496.000 36.250 500.000 ;
    END
  END sram_din0[2]
  PIN sram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 496.000 192.190 500.000 ;
    END
  END sram_din0[30]
  PIN sram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 496.000 196.790 500.000 ;
    END
  END sram_din0[31]
  PIN sram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 496.000 48.670 500.000 ;
    END
  END sram_din0[3]
  PIN sram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 496.000 58.330 500.000 ;
    END
  END sram_din0[4]
  PIN sram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 496.000 66.150 500.000 ;
    END
  END sram_din0[5]
  PIN sram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 496.000 73.970 500.000 ;
    END
  END sram_din0[6]
  PIN sram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 496.000 81.790 500.000 ;
    END
  END sram_din0[7]
  PIN sram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 496.000 89.610 500.000 ;
    END
  END sram_din0[8]
  PIN sram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 496.000 94.210 500.000 ;
    END
  END sram_din0[9]
  PIN sram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 496.000 13.250 500.000 ;
    END
  END sram_dout0[0]
  PIN sram_dout0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 496.000 413.450 500.000 ;
    END
  END sram_dout0[100]
  PIN sram_dout0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 496.000 416.670 500.000 ;
    END
  END sram_dout0[101]
  PIN sram_dout0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 496.000 419.430 500.000 ;
    END
  END sram_dout0[102]
  PIN sram_dout0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 496.000 422.650 500.000 ;
    END
  END sram_dout0[103]
  PIN sram_dout0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 496.000 425.870 500.000 ;
    END
  END sram_dout0[104]
  PIN sram_dout0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 496.000 429.090 500.000 ;
    END
  END sram_dout0[105]
  PIN sram_dout0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 496.000 432.310 500.000 ;
    END
  END sram_dout0[106]
  PIN sram_dout0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 496.000 435.070 500.000 ;
    END
  END sram_dout0[107]
  PIN sram_dout0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 496.000 438.290 500.000 ;
    END
  END sram_dout0[108]
  PIN sram_dout0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 496.000 441.510 500.000 ;
    END
  END sram_dout0[109]
  PIN sram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 496.000 100.190 500.000 ;
    END
  END sram_dout0[10]
  PIN sram_dout0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 496.000 444.730 500.000 ;
    END
  END sram_dout0[110]
  PIN sram_dout0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 496.000 447.490 500.000 ;
    END
  END sram_dout0[111]
  PIN sram_dout0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 496.000 450.710 500.000 ;
    END
  END sram_dout0[112]
  PIN sram_dout0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 496.000 453.930 500.000 ;
    END
  END sram_dout0[113]
  PIN sram_dout0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 496.000 457.150 500.000 ;
    END
  END sram_dout0[114]
  PIN sram_dout0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 496.000 459.910 500.000 ;
    END
  END sram_dout0[115]
  PIN sram_dout0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 496.000 463.130 500.000 ;
    END
  END sram_dout0[116]
  PIN sram_dout0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 496.000 466.350 500.000 ;
    END
  END sram_dout0[117]
  PIN sram_dout0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 496.000 469.570 500.000 ;
    END
  END sram_dout0[118]
  PIN sram_dout0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 496.000 472.790 500.000 ;
    END
  END sram_dout0[119]
  PIN sram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 496.000 104.790 500.000 ;
    END
  END sram_dout0[11]
  PIN sram_dout0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 496.000 475.550 500.000 ;
    END
  END sram_dout0[120]
  PIN sram_dout0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 496.000 478.770 500.000 ;
    END
  END sram_dout0[121]
  PIN sram_dout0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 496.000 481.990 500.000 ;
    END
  END sram_dout0[122]
  PIN sram_dout0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 496.000 485.210 500.000 ;
    END
  END sram_dout0[123]
  PIN sram_dout0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 496.000 487.970 500.000 ;
    END
  END sram_dout0[124]
  PIN sram_dout0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 496.000 491.190 500.000 ;
    END
  END sram_dout0[125]
  PIN sram_dout0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 496.000 494.410 500.000 ;
    END
  END sram_dout0[126]
  PIN sram_dout0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 496.000 497.630 500.000 ;
    END
  END sram_dout0[127]
  PIN sram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 496.000 109.850 500.000 ;
    END
  END sram_dout0[12]
  PIN sram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 496.000 114.450 500.000 ;
    END
  END sram_dout0[13]
  PIN sram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 496.000 119.050 500.000 ;
    END
  END sram_dout0[14]
  PIN sram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 496.000 123.650 500.000 ;
    END
  END sram_dout0[15]
  PIN sram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 496.000 128.250 500.000 ;
    END
  END sram_dout0[16]
  PIN sram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 496.000 132.850 500.000 ;
    END
  END sram_dout0[17]
  PIN sram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 496.000 137.450 500.000 ;
    END
  END sram_dout0[18]
  PIN sram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 496.000 142.510 500.000 ;
    END
  END sram_dout0[19]
  PIN sram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 496.000 25.670 500.000 ;
    END
  END sram_dout0[1]
  PIN sram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 496.000 147.110 500.000 ;
    END
  END sram_dout0[20]
  PIN sram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 496.000 151.710 500.000 ;
    END
  END sram_dout0[21]
  PIN sram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 496.000 156.310 500.000 ;
    END
  END sram_dout0[22]
  PIN sram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 496.000 160.910 500.000 ;
    END
  END sram_dout0[23]
  PIN sram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 496.000 165.510 500.000 ;
    END
  END sram_dout0[24]
  PIN sram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 496.000 170.570 500.000 ;
    END
  END sram_dout0[25]
  PIN sram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 496.000 175.170 500.000 ;
    END
  END sram_dout0[26]
  PIN sram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 496.000 179.770 500.000 ;
    END
  END sram_dout0[27]
  PIN sram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 496.000 184.370 500.000 ;
    END
  END sram_dout0[28]
  PIN sram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 496.000 188.970 500.000 ;
    END
  END sram_dout0[29]
  PIN sram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 496.000 38.090 500.000 ;
    END
  END sram_dout0[2]
  PIN sram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 496.000 193.570 500.000 ;
    END
  END sram_dout0[30]
  PIN sram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 496.000 198.630 500.000 ;
    END
  END sram_dout0[31]
  PIN sram_dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 496.000 201.390 500.000 ;
    END
  END sram_dout0[32]
  PIN sram_dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 496.000 204.610 500.000 ;
    END
  END sram_dout0[33]
  PIN sram_dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 496.000 207.830 500.000 ;
    END
  END sram_dout0[34]
  PIN sram_dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 496.000 211.050 500.000 ;
    END
  END sram_dout0[35]
  PIN sram_dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 496.000 213.810 500.000 ;
    END
  END sram_dout0[36]
  PIN sram_dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 496.000 217.030 500.000 ;
    END
  END sram_dout0[37]
  PIN sram_dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 496.000 220.250 500.000 ;
    END
  END sram_dout0[38]
  PIN sram_dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 496.000 223.470 500.000 ;
    END
  END sram_dout0[39]
  PIN sram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 496.000 50.510 500.000 ;
    END
  END sram_dout0[3]
  PIN sram_dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 496.000 226.690 500.000 ;
    END
  END sram_dout0[40]
  PIN sram_dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 496.000 229.450 500.000 ;
    END
  END sram_dout0[41]
  PIN sram_dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 496.000 232.670 500.000 ;
    END
  END sram_dout0[42]
  PIN sram_dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 496.000 235.890 500.000 ;
    END
  END sram_dout0[43]
  PIN sram_dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 496.000 239.110 500.000 ;
    END
  END sram_dout0[44]
  PIN sram_dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 496.000 241.870 500.000 ;
    END
  END sram_dout0[45]
  PIN sram_dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 496.000 245.090 500.000 ;
    END
  END sram_dout0[46]
  PIN sram_dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 496.000 248.310 500.000 ;
    END
  END sram_dout0[47]
  PIN sram_dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 496.000 251.530 500.000 ;
    END
  END sram_dout0[48]
  PIN sram_dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 496.000 254.290 500.000 ;
    END
  END sram_dout0[49]
  PIN sram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 496.000 59.710 500.000 ;
    END
  END sram_dout0[4]
  PIN sram_dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 496.000 257.510 500.000 ;
    END
  END sram_dout0[50]
  PIN sram_dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 496.000 260.730 500.000 ;
    END
  END sram_dout0[51]
  PIN sram_dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 496.000 263.950 500.000 ;
    END
  END sram_dout0[52]
  PIN sram_dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 496.000 267.170 500.000 ;
    END
  END sram_dout0[53]
  PIN sram_dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 496.000 269.930 500.000 ;
    END
  END sram_dout0[54]
  PIN sram_dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 496.000 273.150 500.000 ;
    END
  END sram_dout0[55]
  PIN sram_dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 496.000 276.370 500.000 ;
    END
  END sram_dout0[56]
  PIN sram_dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 496.000 279.590 500.000 ;
    END
  END sram_dout0[57]
  PIN sram_dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 496.000 282.350 500.000 ;
    END
  END sram_dout0[58]
  PIN sram_dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 496.000 285.570 500.000 ;
    END
  END sram_dout0[59]
  PIN sram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 496.000 67.530 500.000 ;
    END
  END sram_dout0[5]
  PIN sram_dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 496.000 288.790 500.000 ;
    END
  END sram_dout0[60]
  PIN sram_dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 496.000 292.010 500.000 ;
    END
  END sram_dout0[61]
  PIN sram_dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 496.000 295.230 500.000 ;
    END
  END sram_dout0[62]
  PIN sram_dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 496.000 297.990 500.000 ;
    END
  END sram_dout0[63]
  PIN sram_dout0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 496.000 301.210 500.000 ;
    END
  END sram_dout0[64]
  PIN sram_dout0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 496.000 304.430 500.000 ;
    END
  END sram_dout0[65]
  PIN sram_dout0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 496.000 307.650 500.000 ;
    END
  END sram_dout0[66]
  PIN sram_dout0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 496.000 310.410 500.000 ;
    END
  END sram_dout0[67]
  PIN sram_dout0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 496.000 313.630 500.000 ;
    END
  END sram_dout0[68]
  PIN sram_dout0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 496.000 316.850 500.000 ;
    END
  END sram_dout0[69]
  PIN sram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 496.000 75.350 500.000 ;
    END
  END sram_dout0[6]
  PIN sram_dout0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 496.000 320.070 500.000 ;
    END
  END sram_dout0[70]
  PIN sram_dout0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 496.000 322.830 500.000 ;
    END
  END sram_dout0[71]
  PIN sram_dout0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 496.000 326.050 500.000 ;
    END
  END sram_dout0[72]
  PIN sram_dout0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 496.000 329.270 500.000 ;
    END
  END sram_dout0[73]
  PIN sram_dout0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 496.000 332.490 500.000 ;
    END
  END sram_dout0[74]
  PIN sram_dout0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 496.000 335.710 500.000 ;
    END
  END sram_dout0[75]
  PIN sram_dout0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 496.000 338.470 500.000 ;
    END
  END sram_dout0[76]
  PIN sram_dout0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 496.000 341.690 500.000 ;
    END
  END sram_dout0[77]
  PIN sram_dout0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 496.000 344.910 500.000 ;
    END
  END sram_dout0[78]
  PIN sram_dout0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 496.000 348.130 500.000 ;
    END
  END sram_dout0[79]
  PIN sram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 496.000 83.170 500.000 ;
    END
  END sram_dout0[7]
  PIN sram_dout0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 496.000 350.890 500.000 ;
    END
  END sram_dout0[80]
  PIN sram_dout0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 496.000 354.110 500.000 ;
    END
  END sram_dout0[81]
  PIN sram_dout0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 496.000 357.330 500.000 ;
    END
  END sram_dout0[82]
  PIN sram_dout0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 496.000 360.550 500.000 ;
    END
  END sram_dout0[83]
  PIN sram_dout0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 496.000 363.770 500.000 ;
    END
  END sram_dout0[84]
  PIN sram_dout0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 496.000 366.530 500.000 ;
    END
  END sram_dout0[85]
  PIN sram_dout0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 496.000 369.750 500.000 ;
    END
  END sram_dout0[86]
  PIN sram_dout0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 496.000 372.970 500.000 ;
    END
  END sram_dout0[87]
  PIN sram_dout0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 496.000 376.190 500.000 ;
    END
  END sram_dout0[88]
  PIN sram_dout0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 496.000 378.950 500.000 ;
    END
  END sram_dout0[89]
  PIN sram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 496.000 90.990 500.000 ;
    END
  END sram_dout0[8]
  PIN sram_dout0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 496.000 382.170 500.000 ;
    END
  END sram_dout0[90]
  PIN sram_dout0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 496.000 385.390 500.000 ;
    END
  END sram_dout0[91]
  PIN sram_dout0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 496.000 388.610 500.000 ;
    END
  END sram_dout0[92]
  PIN sram_dout0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 496.000 391.370 500.000 ;
    END
  END sram_dout0[93]
  PIN sram_dout0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 496.000 394.590 500.000 ;
    END
  END sram_dout0[94]
  PIN sram_dout0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 496.000 397.810 500.000 ;
    END
  END sram_dout0[95]
  PIN sram_dout0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 496.000 401.030 500.000 ;
    END
  END sram_dout0[96]
  PIN sram_dout0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 496.000 404.250 500.000 ;
    END
  END sram_dout0[97]
  PIN sram_dout0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 496.000 407.010 500.000 ;
    END
  END sram_dout0[98]
  PIN sram_dout0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 496.000 410.230 500.000 ;
    END
  END sram_dout0[99]
  PIN sram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 496.000 95.590 500.000 ;
    END
  END sram_dout0[9]
  PIN sram_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 496.000 14.630 500.000 ;
    END
  END sram_dout1[0]
  PIN sram_dout1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 496.000 414.830 500.000 ;
    END
  END sram_dout1[100]
  PIN sram_dout1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 496.000 418.050 500.000 ;
    END
  END sram_dout1[101]
  PIN sram_dout1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 496.000 421.270 500.000 ;
    END
  END sram_dout1[102]
  PIN sram_dout1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 496.000 424.490 500.000 ;
    END
  END sram_dout1[103]
  PIN sram_dout1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 496.000 427.250 500.000 ;
    END
  END sram_dout1[104]
  PIN sram_dout1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 496.000 430.470 500.000 ;
    END
  END sram_dout1[105]
  PIN sram_dout1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 496.000 433.690 500.000 ;
    END
  END sram_dout1[106]
  PIN sram_dout1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 496.000 436.910 500.000 ;
    END
  END sram_dout1[107]
  PIN sram_dout1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 496.000 439.670 500.000 ;
    END
  END sram_dout1[108]
  PIN sram_dout1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 496.000 442.890 500.000 ;
    END
  END sram_dout1[109]
  PIN sram_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 496.000 102.030 500.000 ;
    END
  END sram_dout1[10]
  PIN sram_dout1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 496.000 446.110 500.000 ;
    END
  END sram_dout1[110]
  PIN sram_dout1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 496.000 449.330 500.000 ;
    END
  END sram_dout1[111]
  PIN sram_dout1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 496.000 452.550 500.000 ;
    END
  END sram_dout1[112]
  PIN sram_dout1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 496.000 455.310 500.000 ;
    END
  END sram_dout1[113]
  PIN sram_dout1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 496.000 458.530 500.000 ;
    END
  END sram_dout1[114]
  PIN sram_dout1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 496.000 461.750 500.000 ;
    END
  END sram_dout1[115]
  PIN sram_dout1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 496.000 464.970 500.000 ;
    END
  END sram_dout1[116]
  PIN sram_dout1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 496.000 467.730 500.000 ;
    END
  END sram_dout1[117]
  PIN sram_dout1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 496.000 470.950 500.000 ;
    END
  END sram_dout1[118]
  PIN sram_dout1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 496.000 474.170 500.000 ;
    END
  END sram_dout1[119]
  PIN sram_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 496.000 106.630 500.000 ;
    END
  END sram_dout1[11]
  PIN sram_dout1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 496.000 477.390 500.000 ;
    END
  END sram_dout1[120]
  PIN sram_dout1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 496.000 480.150 500.000 ;
    END
  END sram_dout1[121]
  PIN sram_dout1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 496.000 483.370 500.000 ;
    END
  END sram_dout1[122]
  PIN sram_dout1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 496.000 486.590 500.000 ;
    END
  END sram_dout1[123]
  PIN sram_dout1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 496.000 489.810 500.000 ;
    END
  END sram_dout1[124]
  PIN sram_dout1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 496.000 493.030 500.000 ;
    END
  END sram_dout1[125]
  PIN sram_dout1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 496.000 495.790 500.000 ;
    END
  END sram_dout1[126]
  PIN sram_dout1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 496.000 499.010 500.000 ;
    END
  END sram_dout1[127]
  PIN sram_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 496.000 111.230 500.000 ;
    END
  END sram_dout1[12]
  PIN sram_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 496.000 115.830 500.000 ;
    END
  END sram_dout1[13]
  PIN sram_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 496.000 120.430 500.000 ;
    END
  END sram_dout1[14]
  PIN sram_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 496.000 125.030 500.000 ;
    END
  END sram_dout1[15]
  PIN sram_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 496.000 130.090 500.000 ;
    END
  END sram_dout1[16]
  PIN sram_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 496.000 134.690 500.000 ;
    END
  END sram_dout1[17]
  PIN sram_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 496.000 139.290 500.000 ;
    END
  END sram_dout1[18]
  PIN sram_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 496.000 143.890 500.000 ;
    END
  END sram_dout1[19]
  PIN sram_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 496.000 27.050 500.000 ;
    END
  END sram_dout1[1]
  PIN sram_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 496.000 148.490 500.000 ;
    END
  END sram_dout1[20]
  PIN sram_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 496.000 153.090 500.000 ;
    END
  END sram_dout1[21]
  PIN sram_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 496.000 158.150 500.000 ;
    END
  END sram_dout1[22]
  PIN sram_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 496.000 162.750 500.000 ;
    END
  END sram_dout1[23]
  PIN sram_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 496.000 167.350 500.000 ;
    END
  END sram_dout1[24]
  PIN sram_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 496.000 171.950 500.000 ;
    END
  END sram_dout1[25]
  PIN sram_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 496.000 176.550 500.000 ;
    END
  END sram_dout1[26]
  PIN sram_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 496.000 181.150 500.000 ;
    END
  END sram_dout1[27]
  PIN sram_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 496.000 185.750 500.000 ;
    END
  END sram_dout1[28]
  PIN sram_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 496.000 190.810 500.000 ;
    END
  END sram_dout1[29]
  PIN sram_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 496.000 39.470 500.000 ;
    END
  END sram_dout1[2]
  PIN sram_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 496.000 195.410 500.000 ;
    END
  END sram_dout1[30]
  PIN sram_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 496.000 200.010 500.000 ;
    END
  END sram_dout1[31]
  PIN sram_dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 496.000 203.230 500.000 ;
    END
  END sram_dout1[32]
  PIN sram_dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 496.000 205.990 500.000 ;
    END
  END sram_dout1[33]
  PIN sram_dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 496.000 209.210 500.000 ;
    END
  END sram_dout1[34]
  PIN sram_dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 496.000 212.430 500.000 ;
    END
  END sram_dout1[35]
  PIN sram_dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 496.000 215.650 500.000 ;
    END
  END sram_dout1[36]
  PIN sram_dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 496.000 218.870 500.000 ;
    END
  END sram_dout1[37]
  PIN sram_dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 496.000 221.630 500.000 ;
    END
  END sram_dout1[38]
  PIN sram_dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 496.000 224.850 500.000 ;
    END
  END sram_dout1[39]
  PIN sram_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 496.000 51.890 500.000 ;
    END
  END sram_dout1[3]
  PIN sram_dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 496.000 228.070 500.000 ;
    END
  END sram_dout1[40]
  PIN sram_dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 496.000 231.290 500.000 ;
    END
  END sram_dout1[41]
  PIN sram_dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 496.000 234.050 500.000 ;
    END
  END sram_dout1[42]
  PIN sram_dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 496.000 237.270 500.000 ;
    END
  END sram_dout1[43]
  PIN sram_dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 496.000 240.490 500.000 ;
    END
  END sram_dout1[44]
  PIN sram_dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 496.000 243.710 500.000 ;
    END
  END sram_dout1[45]
  PIN sram_dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 496.000 246.930 500.000 ;
    END
  END sram_dout1[46]
  PIN sram_dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 496.000 249.690 500.000 ;
    END
  END sram_dout1[47]
  PIN sram_dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 496.000 252.910 500.000 ;
    END
  END sram_dout1[48]
  PIN sram_dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 496.000 256.130 500.000 ;
    END
  END sram_dout1[49]
  PIN sram_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 496.000 61.550 500.000 ;
    END
  END sram_dout1[4]
  PIN sram_dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 496.000 259.350 500.000 ;
    END
  END sram_dout1[50]
  PIN sram_dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 496.000 262.110 500.000 ;
    END
  END sram_dout1[51]
  PIN sram_dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 496.000 265.330 500.000 ;
    END
  END sram_dout1[52]
  PIN sram_dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 496.000 268.550 500.000 ;
    END
  END sram_dout1[53]
  PIN sram_dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 496.000 271.770 500.000 ;
    END
  END sram_dout1[54]
  PIN sram_dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 496.000 274.530 500.000 ;
    END
  END sram_dout1[55]
  PIN sram_dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 496.000 277.750 500.000 ;
    END
  END sram_dout1[56]
  PIN sram_dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 496.000 280.970 500.000 ;
    END
  END sram_dout1[57]
  PIN sram_dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 496.000 284.190 500.000 ;
    END
  END sram_dout1[58]
  PIN sram_dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 496.000 287.410 500.000 ;
    END
  END sram_dout1[59]
  PIN sram_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 496.000 68.910 500.000 ;
    END
  END sram_dout1[5]
  PIN sram_dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 496.000 290.170 500.000 ;
    END
  END sram_dout1[60]
  PIN sram_dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 496.000 293.390 500.000 ;
    END
  END sram_dout1[61]
  PIN sram_dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 496.000 296.610 500.000 ;
    END
  END sram_dout1[62]
  PIN sram_dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 496.000 299.830 500.000 ;
    END
  END sram_dout1[63]
  PIN sram_dout1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 496.000 302.590 500.000 ;
    END
  END sram_dout1[64]
  PIN sram_dout1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 496.000 305.810 500.000 ;
    END
  END sram_dout1[65]
  PIN sram_dout1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 496.000 309.030 500.000 ;
    END
  END sram_dout1[66]
  PIN sram_dout1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 496.000 312.250 500.000 ;
    END
  END sram_dout1[67]
  PIN sram_dout1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 496.000 315.470 500.000 ;
    END
  END sram_dout1[68]
  PIN sram_dout1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 496.000 318.230 500.000 ;
    END
  END sram_dout1[69]
  PIN sram_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 496.000 76.730 500.000 ;
    END
  END sram_dout1[6]
  PIN sram_dout1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 496.000 321.450 500.000 ;
    END
  END sram_dout1[70]
  PIN sram_dout1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 496.000 324.670 500.000 ;
    END
  END sram_dout1[71]
  PIN sram_dout1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 496.000 327.890 500.000 ;
    END
  END sram_dout1[72]
  PIN sram_dout1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 496.000 330.650 500.000 ;
    END
  END sram_dout1[73]
  PIN sram_dout1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 496.000 333.870 500.000 ;
    END
  END sram_dout1[74]
  PIN sram_dout1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 496.000 337.090 500.000 ;
    END
  END sram_dout1[75]
  PIN sram_dout1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 496.000 340.310 500.000 ;
    END
  END sram_dout1[76]
  PIN sram_dout1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 496.000 343.070 500.000 ;
    END
  END sram_dout1[77]
  PIN sram_dout1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 496.000 346.290 500.000 ;
    END
  END sram_dout1[78]
  PIN sram_dout1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 496.000 349.510 500.000 ;
    END
  END sram_dout1[79]
  PIN sram_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 496.000 84.550 500.000 ;
    END
  END sram_dout1[7]
  PIN sram_dout1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 496.000 352.730 500.000 ;
    END
  END sram_dout1[80]
  PIN sram_dout1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 496.000 355.950 500.000 ;
    END
  END sram_dout1[81]
  PIN sram_dout1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 496.000 358.710 500.000 ;
    END
  END sram_dout1[82]
  PIN sram_dout1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 496.000 361.930 500.000 ;
    END
  END sram_dout1[83]
  PIN sram_dout1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 496.000 365.150 500.000 ;
    END
  END sram_dout1[84]
  PIN sram_dout1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 496.000 368.370 500.000 ;
    END
  END sram_dout1[85]
  PIN sram_dout1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 496.000 371.130 500.000 ;
    END
  END sram_dout1[86]
  PIN sram_dout1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 496.000 374.350 500.000 ;
    END
  END sram_dout1[87]
  PIN sram_dout1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 496.000 377.570 500.000 ;
    END
  END sram_dout1[88]
  PIN sram_dout1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 496.000 380.790 500.000 ;
    END
  END sram_dout1[89]
  PIN sram_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 496.000 92.370 500.000 ;
    END
  END sram_dout1[8]
  PIN sram_dout1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 496.000 384.010 500.000 ;
    END
  END sram_dout1[90]
  PIN sram_dout1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 496.000 386.770 500.000 ;
    END
  END sram_dout1[91]
  PIN sram_dout1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 496.000 389.990 500.000 ;
    END
  END sram_dout1[92]
  PIN sram_dout1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 496.000 393.210 500.000 ;
    END
  END sram_dout1[93]
  PIN sram_dout1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 496.000 396.430 500.000 ;
    END
  END sram_dout1[94]
  PIN sram_dout1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 496.000 399.190 500.000 ;
    END
  END sram_dout1[95]
  PIN sram_dout1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 496.000 402.410 500.000 ;
    END
  END sram_dout1[96]
  PIN sram_dout1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 496.000 405.630 500.000 ;
    END
  END sram_dout1[97]
  PIN sram_dout1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 496.000 408.850 500.000 ;
    END
  END sram_dout1[98]
  PIN sram_dout1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 496.000 411.610 500.000 ;
    END
  END sram_dout1[99]
  PIN sram_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 496.000 96.970 500.000 ;
    END
  END sram_dout1[9]
  PIN sram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 496.000 3.590 500.000 ;
    END
  END sram_web0
  PIN sram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 496.000 16.010 500.000 ;
    END
  END sram_wmask0[0]
  PIN sram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 496.000 28.430 500.000 ;
    END
  END sram_wmask0[1]
  PIN sram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 496.000 41.310 500.000 ;
    END
  END sram_wmask0[2]
  PIN sram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 496.000 53.730 500.000 ;
    END
  END sram_wmask0[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.080 500.000 155.680 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 342.760 500.000 343.360 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 217.640 500.000 218.240 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 405.320 500.000 405.920 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 30.640 500.000 31.240 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 280.200 500.000 280.800 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 467.880 500.000 468.480 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 92.520 500.000 93.120 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.070 8.880 497.650 497.380 ;
      LAYER met2 ;
        RECT 0.100 495.720 0.270 497.410 ;
        RECT 1.110 495.720 1.650 497.410 ;
        RECT 2.490 495.720 3.030 497.410 ;
        RECT 3.870 495.720 4.870 497.410 ;
        RECT 5.710 495.720 6.250 497.410 ;
        RECT 7.090 495.720 7.630 497.410 ;
        RECT 8.470 495.720 9.470 497.410 ;
        RECT 10.310 495.720 10.850 497.410 ;
        RECT 11.690 495.720 12.690 497.410 ;
        RECT 13.530 495.720 14.070 497.410 ;
        RECT 14.910 495.720 15.450 497.410 ;
        RECT 16.290 495.720 17.290 497.410 ;
        RECT 18.130 495.720 18.670 497.410 ;
        RECT 19.510 495.720 20.510 497.410 ;
        RECT 21.350 495.720 21.890 497.410 ;
        RECT 22.730 495.720 23.270 497.410 ;
        RECT 24.110 495.720 25.110 497.410 ;
        RECT 25.950 495.720 26.490 497.410 ;
        RECT 27.330 495.720 27.870 497.410 ;
        RECT 28.710 495.720 29.710 497.410 ;
        RECT 30.550 495.720 31.090 497.410 ;
        RECT 31.930 495.720 32.930 497.410 ;
        RECT 33.770 495.720 34.310 497.410 ;
        RECT 35.150 495.720 35.690 497.410 ;
        RECT 36.530 495.720 37.530 497.410 ;
        RECT 38.370 495.720 38.910 497.410 ;
        RECT 39.750 495.720 40.750 497.410 ;
        RECT 41.590 495.720 42.130 497.410 ;
        RECT 42.970 495.720 43.510 497.410 ;
        RECT 44.350 495.720 45.350 497.410 ;
        RECT 46.190 495.720 46.730 497.410 ;
        RECT 47.570 495.720 48.110 497.410 ;
        RECT 48.950 495.720 49.950 497.410 ;
        RECT 50.790 495.720 51.330 497.410 ;
        RECT 52.170 495.720 53.170 497.410 ;
        RECT 54.010 495.720 54.550 497.410 ;
        RECT 55.390 495.720 55.930 497.410 ;
        RECT 56.770 495.720 57.770 497.410 ;
        RECT 58.610 495.720 59.150 497.410 ;
        RECT 59.990 495.720 60.990 497.410 ;
        RECT 61.830 495.720 62.370 497.410 ;
        RECT 63.210 495.720 63.750 497.410 ;
        RECT 64.590 495.720 65.590 497.410 ;
        RECT 66.430 495.720 66.970 497.410 ;
        RECT 67.810 495.720 68.350 497.410 ;
        RECT 69.190 495.720 70.190 497.410 ;
        RECT 71.030 495.720 71.570 497.410 ;
        RECT 72.410 495.720 73.410 497.410 ;
        RECT 74.250 495.720 74.790 497.410 ;
        RECT 75.630 495.720 76.170 497.410 ;
        RECT 77.010 495.720 78.010 497.410 ;
        RECT 78.850 495.720 79.390 497.410 ;
        RECT 80.230 495.720 81.230 497.410 ;
        RECT 82.070 495.720 82.610 497.410 ;
        RECT 83.450 495.720 83.990 497.410 ;
        RECT 84.830 495.720 85.830 497.410 ;
        RECT 86.670 495.720 87.210 497.410 ;
        RECT 88.050 495.720 89.050 497.410 ;
        RECT 89.890 495.720 90.430 497.410 ;
        RECT 91.270 495.720 91.810 497.410 ;
        RECT 92.650 495.720 93.650 497.410 ;
        RECT 94.490 495.720 95.030 497.410 ;
        RECT 95.870 495.720 96.410 497.410 ;
        RECT 97.250 495.720 98.250 497.410 ;
        RECT 99.090 495.720 99.630 497.410 ;
        RECT 100.470 495.720 101.470 497.410 ;
        RECT 102.310 495.720 102.850 497.410 ;
        RECT 103.690 495.720 104.230 497.410 ;
        RECT 105.070 495.720 106.070 497.410 ;
        RECT 106.910 495.720 107.450 497.410 ;
        RECT 108.290 495.720 109.290 497.410 ;
        RECT 110.130 495.720 110.670 497.410 ;
        RECT 111.510 495.720 112.050 497.410 ;
        RECT 112.890 495.720 113.890 497.410 ;
        RECT 114.730 495.720 115.270 497.410 ;
        RECT 116.110 495.720 116.650 497.410 ;
        RECT 117.490 495.720 118.490 497.410 ;
        RECT 119.330 495.720 119.870 497.410 ;
        RECT 120.710 495.720 121.710 497.410 ;
        RECT 122.550 495.720 123.090 497.410 ;
        RECT 123.930 495.720 124.470 497.410 ;
        RECT 125.310 495.720 126.310 497.410 ;
        RECT 127.150 495.720 127.690 497.410 ;
        RECT 128.530 495.720 129.530 497.410 ;
        RECT 130.370 495.720 130.910 497.410 ;
        RECT 131.750 495.720 132.290 497.410 ;
        RECT 133.130 495.720 134.130 497.410 ;
        RECT 134.970 495.720 135.510 497.410 ;
        RECT 136.350 495.720 136.890 497.410 ;
        RECT 137.730 495.720 138.730 497.410 ;
        RECT 139.570 495.720 140.110 497.410 ;
        RECT 140.950 495.720 141.950 497.410 ;
        RECT 142.790 495.720 143.330 497.410 ;
        RECT 144.170 495.720 144.710 497.410 ;
        RECT 145.550 495.720 146.550 497.410 ;
        RECT 147.390 495.720 147.930 497.410 ;
        RECT 148.770 495.720 149.770 497.410 ;
        RECT 150.610 495.720 151.150 497.410 ;
        RECT 151.990 495.720 152.530 497.410 ;
        RECT 153.370 495.720 154.370 497.410 ;
        RECT 155.210 495.720 155.750 497.410 ;
        RECT 156.590 495.720 157.590 497.410 ;
        RECT 158.430 495.720 158.970 497.410 ;
        RECT 159.810 495.720 160.350 497.410 ;
        RECT 161.190 495.720 162.190 497.410 ;
        RECT 163.030 495.720 163.570 497.410 ;
        RECT 164.410 495.720 164.950 497.410 ;
        RECT 165.790 495.720 166.790 497.410 ;
        RECT 167.630 495.720 168.170 497.410 ;
        RECT 169.010 495.720 170.010 497.410 ;
        RECT 170.850 495.720 171.390 497.410 ;
        RECT 172.230 495.720 172.770 497.410 ;
        RECT 173.610 495.720 174.610 497.410 ;
        RECT 175.450 495.720 175.990 497.410 ;
        RECT 176.830 495.720 177.830 497.410 ;
        RECT 178.670 495.720 179.210 497.410 ;
        RECT 180.050 495.720 180.590 497.410 ;
        RECT 181.430 495.720 182.430 497.410 ;
        RECT 183.270 495.720 183.810 497.410 ;
        RECT 184.650 495.720 185.190 497.410 ;
        RECT 186.030 495.720 187.030 497.410 ;
        RECT 187.870 495.720 188.410 497.410 ;
        RECT 189.250 495.720 190.250 497.410 ;
        RECT 191.090 495.720 191.630 497.410 ;
        RECT 192.470 495.720 193.010 497.410 ;
        RECT 193.850 495.720 194.850 497.410 ;
        RECT 195.690 495.720 196.230 497.410 ;
        RECT 197.070 495.720 198.070 497.410 ;
        RECT 198.910 495.720 199.450 497.410 ;
        RECT 200.290 495.720 200.830 497.410 ;
        RECT 201.670 495.720 202.670 497.410 ;
        RECT 203.510 495.720 204.050 497.410 ;
        RECT 204.890 495.720 205.430 497.410 ;
        RECT 206.270 495.720 207.270 497.410 ;
        RECT 208.110 495.720 208.650 497.410 ;
        RECT 209.490 495.720 210.490 497.410 ;
        RECT 211.330 495.720 211.870 497.410 ;
        RECT 212.710 495.720 213.250 497.410 ;
        RECT 214.090 495.720 215.090 497.410 ;
        RECT 215.930 495.720 216.470 497.410 ;
        RECT 217.310 495.720 218.310 497.410 ;
        RECT 219.150 495.720 219.690 497.410 ;
        RECT 220.530 495.720 221.070 497.410 ;
        RECT 221.910 495.720 222.910 497.410 ;
        RECT 223.750 495.720 224.290 497.410 ;
        RECT 225.130 495.720 226.130 497.410 ;
        RECT 226.970 495.720 227.510 497.410 ;
        RECT 228.350 495.720 228.890 497.410 ;
        RECT 229.730 495.720 230.730 497.410 ;
        RECT 231.570 495.720 232.110 497.410 ;
        RECT 232.950 495.720 233.490 497.410 ;
        RECT 234.330 495.720 235.330 497.410 ;
        RECT 236.170 495.720 236.710 497.410 ;
        RECT 237.550 495.720 238.550 497.410 ;
        RECT 239.390 495.720 239.930 497.410 ;
        RECT 240.770 495.720 241.310 497.410 ;
        RECT 242.150 495.720 243.150 497.410 ;
        RECT 243.990 495.720 244.530 497.410 ;
        RECT 245.370 495.720 246.370 497.410 ;
        RECT 247.210 495.720 247.750 497.410 ;
        RECT 248.590 495.720 249.130 497.410 ;
        RECT 249.970 495.720 250.970 497.410 ;
        RECT 251.810 495.720 252.350 497.410 ;
        RECT 253.190 495.720 253.730 497.410 ;
        RECT 254.570 495.720 255.570 497.410 ;
        RECT 256.410 495.720 256.950 497.410 ;
        RECT 257.790 495.720 258.790 497.410 ;
        RECT 259.630 495.720 260.170 497.410 ;
        RECT 261.010 495.720 261.550 497.410 ;
        RECT 262.390 495.720 263.390 497.410 ;
        RECT 264.230 495.720 264.770 497.410 ;
        RECT 265.610 495.720 266.610 497.410 ;
        RECT 267.450 495.720 267.990 497.410 ;
        RECT 268.830 495.720 269.370 497.410 ;
        RECT 270.210 495.720 271.210 497.410 ;
        RECT 272.050 495.720 272.590 497.410 ;
        RECT 273.430 495.720 273.970 497.410 ;
        RECT 274.810 495.720 275.810 497.410 ;
        RECT 276.650 495.720 277.190 497.410 ;
        RECT 278.030 495.720 279.030 497.410 ;
        RECT 279.870 495.720 280.410 497.410 ;
        RECT 281.250 495.720 281.790 497.410 ;
        RECT 282.630 495.720 283.630 497.410 ;
        RECT 284.470 495.720 285.010 497.410 ;
        RECT 285.850 495.720 286.850 497.410 ;
        RECT 287.690 495.720 288.230 497.410 ;
        RECT 289.070 495.720 289.610 497.410 ;
        RECT 290.450 495.720 291.450 497.410 ;
        RECT 292.290 495.720 292.830 497.410 ;
        RECT 293.670 495.720 294.670 497.410 ;
        RECT 295.510 495.720 296.050 497.410 ;
        RECT 296.890 495.720 297.430 497.410 ;
        RECT 298.270 495.720 299.270 497.410 ;
        RECT 300.110 495.720 300.650 497.410 ;
        RECT 301.490 495.720 302.030 497.410 ;
        RECT 302.870 495.720 303.870 497.410 ;
        RECT 304.710 495.720 305.250 497.410 ;
        RECT 306.090 495.720 307.090 497.410 ;
        RECT 307.930 495.720 308.470 497.410 ;
        RECT 309.310 495.720 309.850 497.410 ;
        RECT 310.690 495.720 311.690 497.410 ;
        RECT 312.530 495.720 313.070 497.410 ;
        RECT 313.910 495.720 314.910 497.410 ;
        RECT 315.750 495.720 316.290 497.410 ;
        RECT 317.130 495.720 317.670 497.410 ;
        RECT 318.510 495.720 319.510 497.410 ;
        RECT 320.350 495.720 320.890 497.410 ;
        RECT 321.730 495.720 322.270 497.410 ;
        RECT 323.110 495.720 324.110 497.410 ;
        RECT 324.950 495.720 325.490 497.410 ;
        RECT 326.330 495.720 327.330 497.410 ;
        RECT 328.170 495.720 328.710 497.410 ;
        RECT 329.550 495.720 330.090 497.410 ;
        RECT 330.930 495.720 331.930 497.410 ;
        RECT 332.770 495.720 333.310 497.410 ;
        RECT 334.150 495.720 335.150 497.410 ;
        RECT 335.990 495.720 336.530 497.410 ;
        RECT 337.370 495.720 337.910 497.410 ;
        RECT 338.750 495.720 339.750 497.410 ;
        RECT 340.590 495.720 341.130 497.410 ;
        RECT 341.970 495.720 342.510 497.410 ;
        RECT 343.350 495.720 344.350 497.410 ;
        RECT 345.190 495.720 345.730 497.410 ;
        RECT 346.570 495.720 347.570 497.410 ;
        RECT 348.410 495.720 348.950 497.410 ;
        RECT 349.790 495.720 350.330 497.410 ;
        RECT 351.170 495.720 352.170 497.410 ;
        RECT 353.010 495.720 353.550 497.410 ;
        RECT 354.390 495.720 355.390 497.410 ;
        RECT 356.230 495.720 356.770 497.410 ;
        RECT 357.610 495.720 358.150 497.410 ;
        RECT 358.990 495.720 359.990 497.410 ;
        RECT 360.830 495.720 361.370 497.410 ;
        RECT 362.210 495.720 363.210 497.410 ;
        RECT 364.050 495.720 364.590 497.410 ;
        RECT 365.430 495.720 365.970 497.410 ;
        RECT 366.810 495.720 367.810 497.410 ;
        RECT 368.650 495.720 369.190 497.410 ;
        RECT 370.030 495.720 370.570 497.410 ;
        RECT 371.410 495.720 372.410 497.410 ;
        RECT 373.250 495.720 373.790 497.410 ;
        RECT 374.630 495.720 375.630 497.410 ;
        RECT 376.470 495.720 377.010 497.410 ;
        RECT 377.850 495.720 378.390 497.410 ;
        RECT 379.230 495.720 380.230 497.410 ;
        RECT 381.070 495.720 381.610 497.410 ;
        RECT 382.450 495.720 383.450 497.410 ;
        RECT 384.290 495.720 384.830 497.410 ;
        RECT 385.670 495.720 386.210 497.410 ;
        RECT 387.050 495.720 388.050 497.410 ;
        RECT 388.890 495.720 389.430 497.410 ;
        RECT 390.270 495.720 390.810 497.410 ;
        RECT 391.650 495.720 392.650 497.410 ;
        RECT 393.490 495.720 394.030 497.410 ;
        RECT 394.870 495.720 395.870 497.410 ;
        RECT 396.710 495.720 397.250 497.410 ;
        RECT 398.090 495.720 398.630 497.410 ;
        RECT 399.470 495.720 400.470 497.410 ;
        RECT 401.310 495.720 401.850 497.410 ;
        RECT 402.690 495.720 403.690 497.410 ;
        RECT 404.530 495.720 405.070 497.410 ;
        RECT 405.910 495.720 406.450 497.410 ;
        RECT 407.290 495.720 408.290 497.410 ;
        RECT 409.130 495.720 409.670 497.410 ;
        RECT 410.510 495.720 411.050 497.410 ;
        RECT 411.890 495.720 412.890 497.410 ;
        RECT 413.730 495.720 414.270 497.410 ;
        RECT 415.110 495.720 416.110 497.410 ;
        RECT 416.950 495.720 417.490 497.410 ;
        RECT 418.330 495.720 418.870 497.410 ;
        RECT 419.710 495.720 420.710 497.410 ;
        RECT 421.550 495.720 422.090 497.410 ;
        RECT 422.930 495.720 423.930 497.410 ;
        RECT 424.770 495.720 425.310 497.410 ;
        RECT 426.150 495.720 426.690 497.410 ;
        RECT 427.530 495.720 428.530 497.410 ;
        RECT 429.370 495.720 429.910 497.410 ;
        RECT 430.750 495.720 431.750 497.410 ;
        RECT 432.590 495.720 433.130 497.410 ;
        RECT 433.970 495.720 434.510 497.410 ;
        RECT 435.350 495.720 436.350 497.410 ;
        RECT 437.190 495.720 437.730 497.410 ;
        RECT 438.570 495.720 439.110 497.410 ;
        RECT 439.950 495.720 440.950 497.410 ;
        RECT 441.790 495.720 442.330 497.410 ;
        RECT 443.170 495.720 444.170 497.410 ;
        RECT 445.010 495.720 445.550 497.410 ;
        RECT 446.390 495.720 446.930 497.410 ;
        RECT 447.770 495.720 448.770 497.410 ;
        RECT 449.610 495.720 450.150 497.410 ;
        RECT 450.990 495.720 451.990 497.410 ;
        RECT 452.830 495.720 453.370 497.410 ;
        RECT 454.210 495.720 454.750 497.410 ;
        RECT 455.590 495.720 456.590 497.410 ;
        RECT 457.430 495.720 457.970 497.410 ;
        RECT 458.810 495.720 459.350 497.410 ;
        RECT 460.190 495.720 461.190 497.410 ;
        RECT 462.030 495.720 462.570 497.410 ;
        RECT 463.410 495.720 464.410 497.410 ;
        RECT 465.250 495.720 465.790 497.410 ;
        RECT 466.630 495.720 467.170 497.410 ;
        RECT 468.010 495.720 469.010 497.410 ;
        RECT 469.850 495.720 470.390 497.410 ;
        RECT 471.230 495.720 472.230 497.410 ;
        RECT 473.070 495.720 473.610 497.410 ;
        RECT 474.450 495.720 474.990 497.410 ;
        RECT 475.830 495.720 476.830 497.410 ;
        RECT 477.670 495.720 478.210 497.410 ;
        RECT 479.050 495.720 479.590 497.410 ;
        RECT 480.430 495.720 481.430 497.410 ;
        RECT 482.270 495.720 482.810 497.410 ;
        RECT 483.650 495.720 484.650 497.410 ;
        RECT 485.490 495.720 486.030 497.410 ;
        RECT 486.870 495.720 487.410 497.410 ;
        RECT 488.250 495.720 489.250 497.410 ;
        RECT 490.090 495.720 490.630 497.410 ;
        RECT 491.470 495.720 492.470 497.410 ;
        RECT 493.310 495.720 493.850 497.410 ;
        RECT 494.690 495.720 495.230 497.410 ;
        RECT 496.070 495.720 497.070 497.410 ;
        RECT 0.100 4.280 497.620 495.720 ;
        RECT 0.100 3.670 2.110 4.280 ;
        RECT 2.950 3.670 6.710 4.280 ;
        RECT 7.550 3.670 11.770 4.280 ;
        RECT 12.610 3.670 16.830 4.280 ;
        RECT 17.670 3.670 21.890 4.280 ;
        RECT 22.730 3.670 26.950 4.280 ;
        RECT 27.790 3.670 32.010 4.280 ;
        RECT 32.850 3.670 37.070 4.280 ;
        RECT 37.910 3.670 41.670 4.280 ;
        RECT 42.510 3.670 46.730 4.280 ;
        RECT 47.570 3.670 51.790 4.280 ;
        RECT 52.630 3.670 56.850 4.280 ;
        RECT 57.690 3.670 61.910 4.280 ;
        RECT 62.750 3.670 66.970 4.280 ;
        RECT 67.810 3.670 72.030 4.280 ;
        RECT 72.870 3.670 77.090 4.280 ;
        RECT 77.930 3.670 81.690 4.280 ;
        RECT 82.530 3.670 86.750 4.280 ;
        RECT 87.590 3.670 91.810 4.280 ;
        RECT 92.650 3.670 96.870 4.280 ;
        RECT 97.710 3.670 101.930 4.280 ;
        RECT 102.770 3.670 106.990 4.280 ;
        RECT 107.830 3.670 112.050 4.280 ;
        RECT 112.890 3.670 117.110 4.280 ;
        RECT 117.950 3.670 121.710 4.280 ;
        RECT 122.550 3.670 126.770 4.280 ;
        RECT 127.610 3.670 131.830 4.280 ;
        RECT 132.670 3.670 136.890 4.280 ;
        RECT 137.730 3.670 141.950 4.280 ;
        RECT 142.790 3.670 147.010 4.280 ;
        RECT 147.850 3.670 152.070 4.280 ;
        RECT 152.910 3.670 156.670 4.280 ;
        RECT 157.510 3.670 161.730 4.280 ;
        RECT 162.570 3.670 166.790 4.280 ;
        RECT 167.630 3.670 171.850 4.280 ;
        RECT 172.690 3.670 176.910 4.280 ;
        RECT 177.750 3.670 181.970 4.280 ;
        RECT 182.810 3.670 187.030 4.280 ;
        RECT 187.870 3.670 192.090 4.280 ;
        RECT 192.930 3.670 196.690 4.280 ;
        RECT 197.530 3.670 201.750 4.280 ;
        RECT 202.590 3.670 206.810 4.280 ;
        RECT 207.650 3.670 211.870 4.280 ;
        RECT 212.710 3.670 216.930 4.280 ;
        RECT 217.770 3.670 221.990 4.280 ;
        RECT 222.830 3.670 227.050 4.280 ;
        RECT 227.890 3.670 232.110 4.280 ;
        RECT 232.950 3.670 236.710 4.280 ;
        RECT 237.550 3.670 241.770 4.280 ;
        RECT 242.610 3.670 246.830 4.280 ;
        RECT 247.670 3.670 251.890 4.280 ;
        RECT 252.730 3.670 256.950 4.280 ;
        RECT 257.790 3.670 262.010 4.280 ;
        RECT 262.850 3.670 267.070 4.280 ;
        RECT 267.910 3.670 271.670 4.280 ;
        RECT 272.510 3.670 276.730 4.280 ;
        RECT 277.570 3.670 281.790 4.280 ;
        RECT 282.630 3.670 286.850 4.280 ;
        RECT 287.690 3.670 291.910 4.280 ;
        RECT 292.750 3.670 296.970 4.280 ;
        RECT 297.810 3.670 302.030 4.280 ;
        RECT 302.870 3.670 307.090 4.280 ;
        RECT 307.930 3.670 311.690 4.280 ;
        RECT 312.530 3.670 316.750 4.280 ;
        RECT 317.590 3.670 321.810 4.280 ;
        RECT 322.650 3.670 326.870 4.280 ;
        RECT 327.710 3.670 331.930 4.280 ;
        RECT 332.770 3.670 336.990 4.280 ;
        RECT 337.830 3.670 342.050 4.280 ;
        RECT 342.890 3.670 347.110 4.280 ;
        RECT 347.950 3.670 351.710 4.280 ;
        RECT 352.550 3.670 356.770 4.280 ;
        RECT 357.610 3.670 361.830 4.280 ;
        RECT 362.670 3.670 366.890 4.280 ;
        RECT 367.730 3.670 371.950 4.280 ;
        RECT 372.790 3.670 377.010 4.280 ;
        RECT 377.850 3.670 382.070 4.280 ;
        RECT 382.910 3.670 386.670 4.280 ;
        RECT 387.510 3.670 391.730 4.280 ;
        RECT 392.570 3.670 396.790 4.280 ;
        RECT 397.630 3.670 401.850 4.280 ;
        RECT 402.690 3.670 406.910 4.280 ;
        RECT 407.750 3.670 411.970 4.280 ;
        RECT 412.810 3.670 417.030 4.280 ;
        RECT 417.870 3.670 422.090 4.280 ;
        RECT 422.930 3.670 426.690 4.280 ;
        RECT 427.530 3.670 431.750 4.280 ;
        RECT 432.590 3.670 436.810 4.280 ;
        RECT 437.650 3.670 441.870 4.280 ;
        RECT 442.710 3.670 446.930 4.280 ;
        RECT 447.770 3.670 451.990 4.280 ;
        RECT 452.830 3.670 457.050 4.280 ;
        RECT 457.890 3.670 462.110 4.280 ;
        RECT 462.950 3.670 466.710 4.280 ;
        RECT 467.550 3.670 471.770 4.280 ;
        RECT 472.610 3.670 476.830 4.280 ;
        RECT 477.670 3.670 481.890 4.280 ;
        RECT 482.730 3.670 486.950 4.280 ;
        RECT 487.790 3.670 492.010 4.280 ;
        RECT 492.850 3.670 497.070 4.280 ;
      LAYER met3 ;
        RECT 21.050 468.880 496.000 496.225 ;
        RECT 21.050 467.480 495.600 468.880 ;
        RECT 21.050 406.320 496.000 467.480 ;
        RECT 21.050 404.920 495.600 406.320 ;
        RECT 21.050 343.760 496.000 404.920 ;
        RECT 21.050 342.360 495.600 343.760 ;
        RECT 21.050 281.200 496.000 342.360 ;
        RECT 21.050 279.800 495.600 281.200 ;
        RECT 21.050 218.640 496.000 279.800 ;
        RECT 21.050 217.240 495.600 218.640 ;
        RECT 21.050 156.080 496.000 217.240 ;
        RECT 21.050 154.680 495.600 156.080 ;
        RECT 21.050 93.520 496.000 154.680 ;
        RECT 21.050 92.120 495.600 93.520 ;
        RECT 21.050 31.640 496.000 92.120 ;
        RECT 21.050 30.240 495.600 31.640 ;
        RECT 21.050 10.715 496.000 30.240 ;
      LAYER met4 ;
        RECT 100.575 487.520 402.665 494.865 ;
        RECT 100.575 251.095 174.240 487.520 ;
        RECT 176.640 251.095 251.040 487.520 ;
        RECT 253.440 251.095 327.840 487.520 ;
        RECT 330.240 251.095 402.665 487.520 ;
  END
END Video
END LIBRARY

