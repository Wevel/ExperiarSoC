magic
tech sky130A
magscale 1 2
timestamp 1652993164
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 14 1776 99530 99476
<< metal2 >>
rect 110 99200 166 100000
rect 386 99200 442 100000
rect 662 99200 718 100000
rect 1030 99200 1086 100000
rect 1306 99200 1362 100000
rect 1582 99200 1638 100000
rect 1950 99200 2006 100000
rect 2226 99200 2282 100000
rect 2594 99200 2650 100000
rect 2870 99200 2926 100000
rect 3146 99200 3202 100000
rect 3514 99200 3570 100000
rect 3790 99200 3846 100000
rect 4158 99200 4214 100000
rect 4434 99200 4490 100000
rect 4710 99200 4766 100000
rect 5078 99200 5134 100000
rect 5354 99200 5410 100000
rect 5630 99200 5686 100000
rect 5998 99200 6054 100000
rect 6274 99200 6330 100000
rect 6642 99200 6698 100000
rect 6918 99200 6974 100000
rect 7194 99200 7250 100000
rect 7562 99200 7618 100000
rect 7838 99200 7894 100000
rect 8206 99200 8262 100000
rect 8482 99200 8538 100000
rect 8758 99200 8814 100000
rect 9126 99200 9182 100000
rect 9402 99200 9458 100000
rect 9678 99200 9734 100000
rect 10046 99200 10102 100000
rect 10322 99200 10378 100000
rect 10690 99200 10746 100000
rect 10966 99200 11022 100000
rect 11242 99200 11298 100000
rect 11610 99200 11666 100000
rect 11886 99200 11942 100000
rect 12254 99200 12310 100000
rect 12530 99200 12586 100000
rect 12806 99200 12862 100000
rect 13174 99200 13230 100000
rect 13450 99200 13506 100000
rect 13726 99200 13782 100000
rect 14094 99200 14150 100000
rect 14370 99200 14426 100000
rect 14738 99200 14794 100000
rect 15014 99200 15070 100000
rect 15290 99200 15346 100000
rect 15658 99200 15714 100000
rect 15934 99200 15990 100000
rect 16302 99200 16358 100000
rect 16578 99200 16634 100000
rect 16854 99200 16910 100000
rect 17222 99200 17278 100000
rect 17498 99200 17554 100000
rect 17866 99200 17922 100000
rect 18142 99200 18198 100000
rect 18418 99200 18474 100000
rect 18786 99200 18842 100000
rect 19062 99200 19118 100000
rect 19338 99200 19394 100000
rect 19706 99200 19762 100000
rect 19982 99200 20038 100000
rect 20350 99200 20406 100000
rect 20626 99200 20682 100000
rect 20902 99200 20958 100000
rect 21270 99200 21326 100000
rect 21546 99200 21602 100000
rect 21914 99200 21970 100000
rect 22190 99200 22246 100000
rect 22466 99200 22522 100000
rect 22834 99200 22890 100000
rect 23110 99200 23166 100000
rect 23386 99200 23442 100000
rect 23754 99200 23810 100000
rect 24030 99200 24086 100000
rect 24398 99200 24454 100000
rect 24674 99200 24730 100000
rect 24950 99200 25006 100000
rect 25318 99200 25374 100000
rect 25594 99200 25650 100000
rect 25962 99200 26018 100000
rect 26238 99200 26294 100000
rect 26514 99200 26570 100000
rect 26882 99200 26938 100000
rect 27158 99200 27214 100000
rect 27434 99200 27490 100000
rect 27802 99200 27858 100000
rect 28078 99200 28134 100000
rect 28446 99200 28502 100000
rect 28722 99200 28778 100000
rect 28998 99200 29054 100000
rect 29366 99200 29422 100000
rect 29642 99200 29698 100000
rect 30010 99200 30066 100000
rect 30286 99200 30342 100000
rect 30562 99200 30618 100000
rect 30930 99200 30986 100000
rect 31206 99200 31262 100000
rect 31574 99200 31630 100000
rect 31850 99200 31906 100000
rect 32126 99200 32182 100000
rect 32494 99200 32550 100000
rect 32770 99200 32826 100000
rect 33046 99200 33102 100000
rect 33414 99200 33470 100000
rect 33690 99200 33746 100000
rect 34058 99200 34114 100000
rect 34334 99200 34390 100000
rect 34610 99200 34666 100000
rect 34978 99200 35034 100000
rect 35254 99200 35310 100000
rect 35622 99200 35678 100000
rect 35898 99200 35954 100000
rect 36174 99200 36230 100000
rect 36542 99200 36598 100000
rect 36818 99200 36874 100000
rect 37094 99200 37150 100000
rect 37462 99200 37518 100000
rect 37738 99200 37794 100000
rect 38106 99200 38162 100000
rect 38382 99200 38438 100000
rect 38658 99200 38714 100000
rect 39026 99200 39082 100000
rect 39302 99200 39358 100000
rect 39670 99200 39726 100000
rect 39946 99200 40002 100000
rect 40222 99200 40278 100000
rect 40590 99200 40646 100000
rect 40866 99200 40922 100000
rect 41142 99200 41198 100000
rect 41510 99200 41566 100000
rect 41786 99200 41842 100000
rect 42154 99200 42210 100000
rect 42430 99200 42486 100000
rect 42706 99200 42762 100000
rect 43074 99200 43130 100000
rect 43350 99200 43406 100000
rect 43718 99200 43774 100000
rect 43994 99200 44050 100000
rect 44270 99200 44326 100000
rect 44638 99200 44694 100000
rect 44914 99200 44970 100000
rect 45282 99200 45338 100000
rect 45558 99200 45614 100000
rect 45834 99200 45890 100000
rect 46202 99200 46258 100000
rect 46478 99200 46534 100000
rect 46754 99200 46810 100000
rect 47122 99200 47178 100000
rect 47398 99200 47454 100000
rect 47766 99200 47822 100000
rect 48042 99200 48098 100000
rect 48318 99200 48374 100000
rect 48686 99200 48742 100000
rect 48962 99200 49018 100000
rect 49330 99200 49386 100000
rect 49606 99200 49662 100000
rect 49882 99200 49938 100000
rect 50250 99200 50306 100000
rect 50526 99200 50582 100000
rect 50802 99200 50858 100000
rect 51170 99200 51226 100000
rect 51446 99200 51502 100000
rect 51814 99200 51870 100000
rect 52090 99200 52146 100000
rect 52366 99200 52422 100000
rect 52734 99200 52790 100000
rect 53010 99200 53066 100000
rect 53378 99200 53434 100000
rect 53654 99200 53710 100000
rect 53930 99200 53986 100000
rect 54298 99200 54354 100000
rect 54574 99200 54630 100000
rect 54850 99200 54906 100000
rect 55218 99200 55274 100000
rect 55494 99200 55550 100000
rect 55862 99200 55918 100000
rect 56138 99200 56194 100000
rect 56414 99200 56470 100000
rect 56782 99200 56838 100000
rect 57058 99200 57114 100000
rect 57426 99200 57482 100000
rect 57702 99200 57758 100000
rect 57978 99200 58034 100000
rect 58346 99200 58402 100000
rect 58622 99200 58678 100000
rect 58990 99200 59046 100000
rect 59266 99200 59322 100000
rect 59542 99200 59598 100000
rect 59910 99200 59966 100000
rect 60186 99200 60242 100000
rect 60462 99200 60518 100000
rect 60830 99200 60886 100000
rect 61106 99200 61162 100000
rect 61474 99200 61530 100000
rect 61750 99200 61806 100000
rect 62026 99200 62082 100000
rect 62394 99200 62450 100000
rect 62670 99200 62726 100000
rect 63038 99200 63094 100000
rect 63314 99200 63370 100000
rect 63590 99200 63646 100000
rect 63958 99200 64014 100000
rect 64234 99200 64290 100000
rect 64510 99200 64566 100000
rect 64878 99200 64934 100000
rect 65154 99200 65210 100000
rect 65522 99200 65578 100000
rect 65798 99200 65854 100000
rect 66074 99200 66130 100000
rect 66442 99200 66498 100000
rect 66718 99200 66774 100000
rect 67086 99200 67142 100000
rect 67362 99200 67418 100000
rect 67638 99200 67694 100000
rect 68006 99200 68062 100000
rect 68282 99200 68338 100000
rect 68558 99200 68614 100000
rect 68926 99200 68982 100000
rect 69202 99200 69258 100000
rect 69570 99200 69626 100000
rect 69846 99200 69902 100000
rect 70122 99200 70178 100000
rect 70490 99200 70546 100000
rect 70766 99200 70822 100000
rect 71134 99200 71190 100000
rect 71410 99200 71466 100000
rect 71686 99200 71742 100000
rect 72054 99200 72110 100000
rect 72330 99200 72386 100000
rect 72698 99200 72754 100000
rect 72974 99200 73030 100000
rect 73250 99200 73306 100000
rect 73618 99200 73674 100000
rect 73894 99200 73950 100000
rect 74170 99200 74226 100000
rect 74538 99200 74594 100000
rect 74814 99200 74870 100000
rect 75182 99200 75238 100000
rect 75458 99200 75514 100000
rect 75734 99200 75790 100000
rect 76102 99200 76158 100000
rect 76378 99200 76434 100000
rect 76746 99200 76802 100000
rect 77022 99200 77078 100000
rect 77298 99200 77354 100000
rect 77666 99200 77722 100000
rect 77942 99200 77998 100000
rect 78218 99200 78274 100000
rect 78586 99200 78642 100000
rect 78862 99200 78918 100000
rect 79230 99200 79286 100000
rect 79506 99200 79562 100000
rect 79782 99200 79838 100000
rect 80150 99200 80206 100000
rect 80426 99200 80482 100000
rect 80794 99200 80850 100000
rect 81070 99200 81126 100000
rect 81346 99200 81402 100000
rect 81714 99200 81770 100000
rect 81990 99200 82046 100000
rect 82266 99200 82322 100000
rect 82634 99200 82690 100000
rect 82910 99200 82966 100000
rect 83278 99200 83334 100000
rect 83554 99200 83610 100000
rect 83830 99200 83886 100000
rect 84198 99200 84254 100000
rect 84474 99200 84530 100000
rect 84842 99200 84898 100000
rect 85118 99200 85174 100000
rect 85394 99200 85450 100000
rect 85762 99200 85818 100000
rect 86038 99200 86094 100000
rect 86406 99200 86462 100000
rect 86682 99200 86738 100000
rect 86958 99200 87014 100000
rect 87326 99200 87382 100000
rect 87602 99200 87658 100000
rect 87878 99200 87934 100000
rect 88246 99200 88302 100000
rect 88522 99200 88578 100000
rect 88890 99200 88946 100000
rect 89166 99200 89222 100000
rect 89442 99200 89498 100000
rect 89810 99200 89866 100000
rect 90086 99200 90142 100000
rect 90454 99200 90510 100000
rect 90730 99200 90786 100000
rect 91006 99200 91062 100000
rect 91374 99200 91430 100000
rect 91650 99200 91706 100000
rect 91926 99200 91982 100000
rect 92294 99200 92350 100000
rect 92570 99200 92626 100000
rect 92938 99200 92994 100000
rect 93214 99200 93270 100000
rect 93490 99200 93546 100000
rect 93858 99200 93914 100000
rect 94134 99200 94190 100000
rect 94502 99200 94558 100000
rect 94778 99200 94834 100000
rect 95054 99200 95110 100000
rect 95422 99200 95478 100000
rect 95698 99200 95754 100000
rect 95974 99200 96030 100000
rect 96342 99200 96398 100000
rect 96618 99200 96674 100000
rect 96986 99200 97042 100000
rect 97262 99200 97318 100000
rect 97538 99200 97594 100000
rect 97906 99200 97962 100000
rect 98182 99200 98238 100000
rect 98550 99200 98606 100000
rect 98826 99200 98882 100000
rect 99102 99200 99158 100000
rect 99470 99200 99526 100000
rect 99746 99200 99802 100000
rect 478 0 534 800
rect 1398 0 1454 800
rect 2410 0 2466 800
rect 3422 0 3478 800
rect 4434 0 4490 800
rect 5446 0 5502 800
rect 6458 0 6514 800
rect 7470 0 7526 800
rect 8390 0 8446 800
rect 9402 0 9458 800
rect 10414 0 10470 800
rect 11426 0 11482 800
rect 12438 0 12494 800
rect 13450 0 13506 800
rect 14462 0 14518 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17406 0 17462 800
rect 18418 0 18474 800
rect 19430 0 19486 800
rect 20442 0 20498 800
rect 21454 0 21510 800
rect 22466 0 22522 800
rect 23478 0 23534 800
rect 24398 0 24454 800
rect 25410 0 25466 800
rect 26422 0 26478 800
rect 27434 0 27490 800
rect 28446 0 28502 800
rect 29458 0 29514 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32402 0 32458 800
rect 33414 0 33470 800
rect 34426 0 34482 800
rect 35438 0 35494 800
rect 36450 0 36506 800
rect 37462 0 37518 800
rect 38474 0 38530 800
rect 39394 0 39450 800
rect 40406 0 40462 800
rect 41418 0 41474 800
rect 42430 0 42486 800
rect 43442 0 43498 800
rect 44454 0 44510 800
rect 45466 0 45522 800
rect 46478 0 46534 800
rect 47398 0 47454 800
rect 48410 0 48466 800
rect 49422 0 49478 800
rect 50434 0 50490 800
rect 51446 0 51502 800
rect 52458 0 52514 800
rect 53470 0 53526 800
rect 54390 0 54446 800
rect 55402 0 55458 800
rect 56414 0 56470 800
rect 57426 0 57482 800
rect 58438 0 58494 800
rect 59450 0 59506 800
rect 60462 0 60518 800
rect 61474 0 61530 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68466 0 68522 800
rect 69478 0 69534 800
rect 70398 0 70454 800
rect 71410 0 71466 800
rect 72422 0 72478 800
rect 73434 0 73490 800
rect 74446 0 74502 800
rect 75458 0 75514 800
rect 76470 0 76526 800
rect 77390 0 77446 800
rect 78402 0 78458 800
rect 79414 0 79470 800
rect 80426 0 80482 800
rect 81438 0 81494 800
rect 82450 0 82506 800
rect 83462 0 83518 800
rect 84474 0 84530 800
rect 85394 0 85450 800
rect 86406 0 86462 800
rect 87418 0 87474 800
rect 88430 0 88486 800
rect 89442 0 89498 800
rect 90454 0 90510 800
rect 91466 0 91522 800
rect 92478 0 92534 800
rect 93398 0 93454 800
rect 94410 0 94466 800
rect 95422 0 95478 800
rect 96434 0 96490 800
rect 97446 0 97502 800
rect 98458 0 98514 800
rect 99470 0 99526 800
<< obsm2 >>
rect 20 99144 54 99482
rect 222 99144 330 99482
rect 498 99144 606 99482
rect 774 99144 974 99482
rect 1142 99144 1250 99482
rect 1418 99144 1526 99482
rect 1694 99144 1894 99482
rect 2062 99144 2170 99482
rect 2338 99144 2538 99482
rect 2706 99144 2814 99482
rect 2982 99144 3090 99482
rect 3258 99144 3458 99482
rect 3626 99144 3734 99482
rect 3902 99144 4102 99482
rect 4270 99144 4378 99482
rect 4546 99144 4654 99482
rect 4822 99144 5022 99482
rect 5190 99144 5298 99482
rect 5466 99144 5574 99482
rect 5742 99144 5942 99482
rect 6110 99144 6218 99482
rect 6386 99144 6586 99482
rect 6754 99144 6862 99482
rect 7030 99144 7138 99482
rect 7306 99144 7506 99482
rect 7674 99144 7782 99482
rect 7950 99144 8150 99482
rect 8318 99144 8426 99482
rect 8594 99144 8702 99482
rect 8870 99144 9070 99482
rect 9238 99144 9346 99482
rect 9514 99144 9622 99482
rect 9790 99144 9990 99482
rect 10158 99144 10266 99482
rect 10434 99144 10634 99482
rect 10802 99144 10910 99482
rect 11078 99144 11186 99482
rect 11354 99144 11554 99482
rect 11722 99144 11830 99482
rect 11998 99144 12198 99482
rect 12366 99144 12474 99482
rect 12642 99144 12750 99482
rect 12918 99144 13118 99482
rect 13286 99144 13394 99482
rect 13562 99144 13670 99482
rect 13838 99144 14038 99482
rect 14206 99144 14314 99482
rect 14482 99144 14682 99482
rect 14850 99144 14958 99482
rect 15126 99144 15234 99482
rect 15402 99144 15602 99482
rect 15770 99144 15878 99482
rect 16046 99144 16246 99482
rect 16414 99144 16522 99482
rect 16690 99144 16798 99482
rect 16966 99144 17166 99482
rect 17334 99144 17442 99482
rect 17610 99144 17810 99482
rect 17978 99144 18086 99482
rect 18254 99144 18362 99482
rect 18530 99144 18730 99482
rect 18898 99144 19006 99482
rect 19174 99144 19282 99482
rect 19450 99144 19650 99482
rect 19818 99144 19926 99482
rect 20094 99144 20294 99482
rect 20462 99144 20570 99482
rect 20738 99144 20846 99482
rect 21014 99144 21214 99482
rect 21382 99144 21490 99482
rect 21658 99144 21858 99482
rect 22026 99144 22134 99482
rect 22302 99144 22410 99482
rect 22578 99144 22778 99482
rect 22946 99144 23054 99482
rect 23222 99144 23330 99482
rect 23498 99144 23698 99482
rect 23866 99144 23974 99482
rect 24142 99144 24342 99482
rect 24510 99144 24618 99482
rect 24786 99144 24894 99482
rect 25062 99144 25262 99482
rect 25430 99144 25538 99482
rect 25706 99144 25906 99482
rect 26074 99144 26182 99482
rect 26350 99144 26458 99482
rect 26626 99144 26826 99482
rect 26994 99144 27102 99482
rect 27270 99144 27378 99482
rect 27546 99144 27746 99482
rect 27914 99144 28022 99482
rect 28190 99144 28390 99482
rect 28558 99144 28666 99482
rect 28834 99144 28942 99482
rect 29110 99144 29310 99482
rect 29478 99144 29586 99482
rect 29754 99144 29954 99482
rect 30122 99144 30230 99482
rect 30398 99144 30506 99482
rect 30674 99144 30874 99482
rect 31042 99144 31150 99482
rect 31318 99144 31518 99482
rect 31686 99144 31794 99482
rect 31962 99144 32070 99482
rect 32238 99144 32438 99482
rect 32606 99144 32714 99482
rect 32882 99144 32990 99482
rect 33158 99144 33358 99482
rect 33526 99144 33634 99482
rect 33802 99144 34002 99482
rect 34170 99144 34278 99482
rect 34446 99144 34554 99482
rect 34722 99144 34922 99482
rect 35090 99144 35198 99482
rect 35366 99144 35566 99482
rect 35734 99144 35842 99482
rect 36010 99144 36118 99482
rect 36286 99144 36486 99482
rect 36654 99144 36762 99482
rect 36930 99144 37038 99482
rect 37206 99144 37406 99482
rect 37574 99144 37682 99482
rect 37850 99144 38050 99482
rect 38218 99144 38326 99482
rect 38494 99144 38602 99482
rect 38770 99144 38970 99482
rect 39138 99144 39246 99482
rect 39414 99144 39614 99482
rect 39782 99144 39890 99482
rect 40058 99144 40166 99482
rect 40334 99144 40534 99482
rect 40702 99144 40810 99482
rect 40978 99144 41086 99482
rect 41254 99144 41454 99482
rect 41622 99144 41730 99482
rect 41898 99144 42098 99482
rect 42266 99144 42374 99482
rect 42542 99144 42650 99482
rect 42818 99144 43018 99482
rect 43186 99144 43294 99482
rect 43462 99144 43662 99482
rect 43830 99144 43938 99482
rect 44106 99144 44214 99482
rect 44382 99144 44582 99482
rect 44750 99144 44858 99482
rect 45026 99144 45226 99482
rect 45394 99144 45502 99482
rect 45670 99144 45778 99482
rect 45946 99144 46146 99482
rect 46314 99144 46422 99482
rect 46590 99144 46698 99482
rect 46866 99144 47066 99482
rect 47234 99144 47342 99482
rect 47510 99144 47710 99482
rect 47878 99144 47986 99482
rect 48154 99144 48262 99482
rect 48430 99144 48630 99482
rect 48798 99144 48906 99482
rect 49074 99144 49274 99482
rect 49442 99144 49550 99482
rect 49718 99144 49826 99482
rect 49994 99144 50194 99482
rect 50362 99144 50470 99482
rect 50638 99144 50746 99482
rect 50914 99144 51114 99482
rect 51282 99144 51390 99482
rect 51558 99144 51758 99482
rect 51926 99144 52034 99482
rect 52202 99144 52310 99482
rect 52478 99144 52678 99482
rect 52846 99144 52954 99482
rect 53122 99144 53322 99482
rect 53490 99144 53598 99482
rect 53766 99144 53874 99482
rect 54042 99144 54242 99482
rect 54410 99144 54518 99482
rect 54686 99144 54794 99482
rect 54962 99144 55162 99482
rect 55330 99144 55438 99482
rect 55606 99144 55806 99482
rect 55974 99144 56082 99482
rect 56250 99144 56358 99482
rect 56526 99144 56726 99482
rect 56894 99144 57002 99482
rect 57170 99144 57370 99482
rect 57538 99144 57646 99482
rect 57814 99144 57922 99482
rect 58090 99144 58290 99482
rect 58458 99144 58566 99482
rect 58734 99144 58934 99482
rect 59102 99144 59210 99482
rect 59378 99144 59486 99482
rect 59654 99144 59854 99482
rect 60022 99144 60130 99482
rect 60298 99144 60406 99482
rect 60574 99144 60774 99482
rect 60942 99144 61050 99482
rect 61218 99144 61418 99482
rect 61586 99144 61694 99482
rect 61862 99144 61970 99482
rect 62138 99144 62338 99482
rect 62506 99144 62614 99482
rect 62782 99144 62982 99482
rect 63150 99144 63258 99482
rect 63426 99144 63534 99482
rect 63702 99144 63902 99482
rect 64070 99144 64178 99482
rect 64346 99144 64454 99482
rect 64622 99144 64822 99482
rect 64990 99144 65098 99482
rect 65266 99144 65466 99482
rect 65634 99144 65742 99482
rect 65910 99144 66018 99482
rect 66186 99144 66386 99482
rect 66554 99144 66662 99482
rect 66830 99144 67030 99482
rect 67198 99144 67306 99482
rect 67474 99144 67582 99482
rect 67750 99144 67950 99482
rect 68118 99144 68226 99482
rect 68394 99144 68502 99482
rect 68670 99144 68870 99482
rect 69038 99144 69146 99482
rect 69314 99144 69514 99482
rect 69682 99144 69790 99482
rect 69958 99144 70066 99482
rect 70234 99144 70434 99482
rect 70602 99144 70710 99482
rect 70878 99144 71078 99482
rect 71246 99144 71354 99482
rect 71522 99144 71630 99482
rect 71798 99144 71998 99482
rect 72166 99144 72274 99482
rect 72442 99144 72642 99482
rect 72810 99144 72918 99482
rect 73086 99144 73194 99482
rect 73362 99144 73562 99482
rect 73730 99144 73838 99482
rect 74006 99144 74114 99482
rect 74282 99144 74482 99482
rect 74650 99144 74758 99482
rect 74926 99144 75126 99482
rect 75294 99144 75402 99482
rect 75570 99144 75678 99482
rect 75846 99144 76046 99482
rect 76214 99144 76322 99482
rect 76490 99144 76690 99482
rect 76858 99144 76966 99482
rect 77134 99144 77242 99482
rect 77410 99144 77610 99482
rect 77778 99144 77886 99482
rect 78054 99144 78162 99482
rect 78330 99144 78530 99482
rect 78698 99144 78806 99482
rect 78974 99144 79174 99482
rect 79342 99144 79450 99482
rect 79618 99144 79726 99482
rect 79894 99144 80094 99482
rect 80262 99144 80370 99482
rect 80538 99144 80738 99482
rect 80906 99144 81014 99482
rect 81182 99144 81290 99482
rect 81458 99144 81658 99482
rect 81826 99144 81934 99482
rect 82102 99144 82210 99482
rect 82378 99144 82578 99482
rect 82746 99144 82854 99482
rect 83022 99144 83222 99482
rect 83390 99144 83498 99482
rect 83666 99144 83774 99482
rect 83942 99144 84142 99482
rect 84310 99144 84418 99482
rect 84586 99144 84786 99482
rect 84954 99144 85062 99482
rect 85230 99144 85338 99482
rect 85506 99144 85706 99482
rect 85874 99144 85982 99482
rect 86150 99144 86350 99482
rect 86518 99144 86626 99482
rect 86794 99144 86902 99482
rect 87070 99144 87270 99482
rect 87438 99144 87546 99482
rect 87714 99144 87822 99482
rect 87990 99144 88190 99482
rect 88358 99144 88466 99482
rect 88634 99144 88834 99482
rect 89002 99144 89110 99482
rect 89278 99144 89386 99482
rect 89554 99144 89754 99482
rect 89922 99144 90030 99482
rect 90198 99144 90398 99482
rect 90566 99144 90674 99482
rect 90842 99144 90950 99482
rect 91118 99144 91318 99482
rect 91486 99144 91594 99482
rect 91762 99144 91870 99482
rect 92038 99144 92238 99482
rect 92406 99144 92514 99482
rect 92682 99144 92882 99482
rect 93050 99144 93158 99482
rect 93326 99144 93434 99482
rect 93602 99144 93802 99482
rect 93970 99144 94078 99482
rect 94246 99144 94446 99482
rect 94614 99144 94722 99482
rect 94890 99144 94998 99482
rect 95166 99144 95366 99482
rect 95534 99144 95642 99482
rect 95810 99144 95918 99482
rect 96086 99144 96286 99482
rect 96454 99144 96562 99482
rect 96730 99144 96930 99482
rect 97098 99144 97206 99482
rect 97374 99144 97482 99482
rect 97650 99144 97850 99482
rect 98018 99144 98126 99482
rect 98294 99144 98494 99482
rect 98662 99144 98770 99482
rect 98938 99144 99046 99482
rect 99214 99144 99414 99482
rect 20 856 99524 99144
rect 20 734 422 856
rect 590 734 1342 856
rect 1510 734 2354 856
rect 2522 734 3366 856
rect 3534 734 4378 856
rect 4546 734 5390 856
rect 5558 734 6402 856
rect 6570 734 7414 856
rect 7582 734 8334 856
rect 8502 734 9346 856
rect 9514 734 10358 856
rect 10526 734 11370 856
rect 11538 734 12382 856
rect 12550 734 13394 856
rect 13562 734 14406 856
rect 14574 734 15418 856
rect 15586 734 16338 856
rect 16506 734 17350 856
rect 17518 734 18362 856
rect 18530 734 19374 856
rect 19542 734 20386 856
rect 20554 734 21398 856
rect 21566 734 22410 856
rect 22578 734 23422 856
rect 23590 734 24342 856
rect 24510 734 25354 856
rect 25522 734 26366 856
rect 26534 734 27378 856
rect 27546 734 28390 856
rect 28558 734 29402 856
rect 29570 734 30414 856
rect 30582 734 31334 856
rect 31502 734 32346 856
rect 32514 734 33358 856
rect 33526 734 34370 856
rect 34538 734 35382 856
rect 35550 734 36394 856
rect 36562 734 37406 856
rect 37574 734 38418 856
rect 38586 734 39338 856
rect 39506 734 40350 856
rect 40518 734 41362 856
rect 41530 734 42374 856
rect 42542 734 43386 856
rect 43554 734 44398 856
rect 44566 734 45410 856
rect 45578 734 46422 856
rect 46590 734 47342 856
rect 47510 734 48354 856
rect 48522 734 49366 856
rect 49534 734 50378 856
rect 50546 734 51390 856
rect 51558 734 52402 856
rect 52570 734 53414 856
rect 53582 734 54334 856
rect 54502 734 55346 856
rect 55514 734 56358 856
rect 56526 734 57370 856
rect 57538 734 58382 856
rect 58550 734 59394 856
rect 59562 734 60406 856
rect 60574 734 61418 856
rect 61586 734 62338 856
rect 62506 734 63350 856
rect 63518 734 64362 856
rect 64530 734 65374 856
rect 65542 734 66386 856
rect 66554 734 67398 856
rect 67566 734 68410 856
rect 68578 734 69422 856
rect 69590 734 70342 856
rect 70510 734 71354 856
rect 71522 734 72366 856
rect 72534 734 73378 856
rect 73546 734 74390 856
rect 74558 734 75402 856
rect 75570 734 76414 856
rect 76582 734 77334 856
rect 77502 734 78346 856
rect 78514 734 79358 856
rect 79526 734 80370 856
rect 80538 734 81382 856
rect 81550 734 82394 856
rect 82562 734 83406 856
rect 83574 734 84418 856
rect 84586 734 85338 856
rect 85506 734 86350 856
rect 86518 734 87362 856
rect 87530 734 88374 856
rect 88542 734 89386 856
rect 89554 734 90398 856
rect 90566 734 91410 856
rect 91578 734 92422 856
rect 92590 734 93342 856
rect 93510 734 94354 856
rect 94522 734 95366 856
rect 95534 734 96378 856
rect 96546 734 97390 856
rect 97558 734 98402 856
rect 98570 734 99414 856
<< metal3 >>
rect 99200 93576 100000 93696
rect 99200 81064 100000 81184
rect 99200 68552 100000 68672
rect 99200 56040 100000 56160
rect 99200 43528 100000 43648
rect 99200 31016 100000 31136
rect 99200 18504 100000 18624
rect 99200 6128 100000 6248
<< obsm3 >>
rect 4210 93776 99200 99245
rect 4210 93496 99120 93776
rect 4210 81264 99200 93496
rect 4210 80984 99120 81264
rect 4210 68752 99200 80984
rect 4210 68472 99120 68752
rect 4210 56240 99200 68472
rect 4210 55960 99120 56240
rect 4210 43728 99200 55960
rect 4210 43448 99120 43728
rect 4210 31216 99200 43448
rect 4210 30936 99120 31216
rect 4210 18704 99200 30936
rect 4210 18424 99120 18704
rect 4210 6328 99200 18424
rect 4210 6048 99120 6328
rect 4210 2143 99200 6048
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 20115 97504 80533 98973
rect 20115 50219 34848 97504
rect 35328 50219 50208 97504
rect 50688 50219 65568 97504
rect 66048 50219 80533 97504
<< labels >>
rlabel metal2 s 1030 99200 1086 100000 6 sram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 3514 99200 3570 100000 6 sram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 5998 99200 6054 100000 6 sram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 8482 99200 8538 100000 6 sram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 10966 99200 11022 100000 6 sram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 12530 99200 12586 100000 6 sram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 14094 99200 14150 100000 6 sram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 15658 99200 15714 100000 6 sram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 17222 99200 17278 100000 6 sram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 1306 99200 1362 100000 6 sram_addr1[0]
port 10 nsew signal output
rlabel metal2 s 3790 99200 3846 100000 6 sram_addr1[1]
port 11 nsew signal output
rlabel metal2 s 6274 99200 6330 100000 6 sram_addr1[2]
port 12 nsew signal output
rlabel metal2 s 8758 99200 8814 100000 6 sram_addr1[3]
port 13 nsew signal output
rlabel metal2 s 11242 99200 11298 100000 6 sram_addr1[4]
port 14 nsew signal output
rlabel metal2 s 12806 99200 12862 100000 6 sram_addr1[5]
port 15 nsew signal output
rlabel metal2 s 14370 99200 14426 100000 6 sram_addr1[6]
port 16 nsew signal output
rlabel metal2 s 15934 99200 15990 100000 6 sram_addr1[7]
port 17 nsew signal output
rlabel metal2 s 17498 99200 17554 100000 6 sram_addr1[8]
port 18 nsew signal output
rlabel metal2 s 110 99200 166 100000 6 sram_clk0
port 19 nsew signal output
rlabel metal2 s 386 99200 442 100000 6 sram_clk1
port 20 nsew signal output
rlabel metal2 s 1582 99200 1638 100000 6 sram_csb0[0]
port 21 nsew signal output
rlabel metal2 s 4158 99200 4214 100000 6 sram_csb0[1]
port 22 nsew signal output
rlabel metal2 s 6642 99200 6698 100000 6 sram_csb0[2]
port 23 nsew signal output
rlabel metal2 s 9126 99200 9182 100000 6 sram_csb0[3]
port 24 nsew signal output
rlabel metal2 s 1950 99200 2006 100000 6 sram_csb1[0]
port 25 nsew signal output
rlabel metal2 s 4434 99200 4490 100000 6 sram_csb1[1]
port 26 nsew signal output
rlabel metal2 s 6918 99200 6974 100000 6 sram_csb1[2]
port 27 nsew signal output
rlabel metal2 s 9402 99200 9458 100000 6 sram_csb1[3]
port 28 nsew signal output
rlabel metal2 s 2226 99200 2282 100000 6 sram_din0[0]
port 29 nsew signal output
rlabel metal2 s 19706 99200 19762 100000 6 sram_din0[10]
port 30 nsew signal output
rlabel metal2 s 20626 99200 20682 100000 6 sram_din0[11]
port 31 nsew signal output
rlabel metal2 s 21546 99200 21602 100000 6 sram_din0[12]
port 32 nsew signal output
rlabel metal2 s 22466 99200 22522 100000 6 sram_din0[13]
port 33 nsew signal output
rlabel metal2 s 23386 99200 23442 100000 6 sram_din0[14]
port 34 nsew signal output
rlabel metal2 s 24398 99200 24454 100000 6 sram_din0[15]
port 35 nsew signal output
rlabel metal2 s 25318 99200 25374 100000 6 sram_din0[16]
port 36 nsew signal output
rlabel metal2 s 26238 99200 26294 100000 6 sram_din0[17]
port 37 nsew signal output
rlabel metal2 s 27158 99200 27214 100000 6 sram_din0[18]
port 38 nsew signal output
rlabel metal2 s 28078 99200 28134 100000 6 sram_din0[19]
port 39 nsew signal output
rlabel metal2 s 4710 99200 4766 100000 6 sram_din0[1]
port 40 nsew signal output
rlabel metal2 s 28998 99200 29054 100000 6 sram_din0[20]
port 41 nsew signal output
rlabel metal2 s 30010 99200 30066 100000 6 sram_din0[21]
port 42 nsew signal output
rlabel metal2 s 30930 99200 30986 100000 6 sram_din0[22]
port 43 nsew signal output
rlabel metal2 s 31850 99200 31906 100000 6 sram_din0[23]
port 44 nsew signal output
rlabel metal2 s 32770 99200 32826 100000 6 sram_din0[24]
port 45 nsew signal output
rlabel metal2 s 33690 99200 33746 100000 6 sram_din0[25]
port 46 nsew signal output
rlabel metal2 s 34610 99200 34666 100000 6 sram_din0[26]
port 47 nsew signal output
rlabel metal2 s 35622 99200 35678 100000 6 sram_din0[27]
port 48 nsew signal output
rlabel metal2 s 36542 99200 36598 100000 6 sram_din0[28]
port 49 nsew signal output
rlabel metal2 s 37462 99200 37518 100000 6 sram_din0[29]
port 50 nsew signal output
rlabel metal2 s 7194 99200 7250 100000 6 sram_din0[2]
port 51 nsew signal output
rlabel metal2 s 38382 99200 38438 100000 6 sram_din0[30]
port 52 nsew signal output
rlabel metal2 s 39302 99200 39358 100000 6 sram_din0[31]
port 53 nsew signal output
rlabel metal2 s 9678 99200 9734 100000 6 sram_din0[3]
port 54 nsew signal output
rlabel metal2 s 11610 99200 11666 100000 6 sram_din0[4]
port 55 nsew signal output
rlabel metal2 s 13174 99200 13230 100000 6 sram_din0[5]
port 56 nsew signal output
rlabel metal2 s 14738 99200 14794 100000 6 sram_din0[6]
port 57 nsew signal output
rlabel metal2 s 16302 99200 16358 100000 6 sram_din0[7]
port 58 nsew signal output
rlabel metal2 s 17866 99200 17922 100000 6 sram_din0[8]
port 59 nsew signal output
rlabel metal2 s 18786 99200 18842 100000 6 sram_din0[9]
port 60 nsew signal output
rlabel metal2 s 2594 99200 2650 100000 6 sram_dout0[0]
port 61 nsew signal input
rlabel metal2 s 82634 99200 82690 100000 6 sram_dout0[100]
port 62 nsew signal input
rlabel metal2 s 83278 99200 83334 100000 6 sram_dout0[101]
port 63 nsew signal input
rlabel metal2 s 83830 99200 83886 100000 6 sram_dout0[102]
port 64 nsew signal input
rlabel metal2 s 84474 99200 84530 100000 6 sram_dout0[103]
port 65 nsew signal input
rlabel metal2 s 85118 99200 85174 100000 6 sram_dout0[104]
port 66 nsew signal input
rlabel metal2 s 85762 99200 85818 100000 6 sram_dout0[105]
port 67 nsew signal input
rlabel metal2 s 86406 99200 86462 100000 6 sram_dout0[106]
port 68 nsew signal input
rlabel metal2 s 86958 99200 87014 100000 6 sram_dout0[107]
port 69 nsew signal input
rlabel metal2 s 87602 99200 87658 100000 6 sram_dout0[108]
port 70 nsew signal input
rlabel metal2 s 88246 99200 88302 100000 6 sram_dout0[109]
port 71 nsew signal input
rlabel metal2 s 19982 99200 20038 100000 6 sram_dout0[10]
port 72 nsew signal input
rlabel metal2 s 88890 99200 88946 100000 6 sram_dout0[110]
port 73 nsew signal input
rlabel metal2 s 89442 99200 89498 100000 6 sram_dout0[111]
port 74 nsew signal input
rlabel metal2 s 90086 99200 90142 100000 6 sram_dout0[112]
port 75 nsew signal input
rlabel metal2 s 90730 99200 90786 100000 6 sram_dout0[113]
port 76 nsew signal input
rlabel metal2 s 91374 99200 91430 100000 6 sram_dout0[114]
port 77 nsew signal input
rlabel metal2 s 91926 99200 91982 100000 6 sram_dout0[115]
port 78 nsew signal input
rlabel metal2 s 92570 99200 92626 100000 6 sram_dout0[116]
port 79 nsew signal input
rlabel metal2 s 93214 99200 93270 100000 6 sram_dout0[117]
port 80 nsew signal input
rlabel metal2 s 93858 99200 93914 100000 6 sram_dout0[118]
port 81 nsew signal input
rlabel metal2 s 94502 99200 94558 100000 6 sram_dout0[119]
port 82 nsew signal input
rlabel metal2 s 20902 99200 20958 100000 6 sram_dout0[11]
port 83 nsew signal input
rlabel metal2 s 95054 99200 95110 100000 6 sram_dout0[120]
port 84 nsew signal input
rlabel metal2 s 95698 99200 95754 100000 6 sram_dout0[121]
port 85 nsew signal input
rlabel metal2 s 96342 99200 96398 100000 6 sram_dout0[122]
port 86 nsew signal input
rlabel metal2 s 96986 99200 97042 100000 6 sram_dout0[123]
port 87 nsew signal input
rlabel metal2 s 97538 99200 97594 100000 6 sram_dout0[124]
port 88 nsew signal input
rlabel metal2 s 98182 99200 98238 100000 6 sram_dout0[125]
port 89 nsew signal input
rlabel metal2 s 98826 99200 98882 100000 6 sram_dout0[126]
port 90 nsew signal input
rlabel metal2 s 99470 99200 99526 100000 6 sram_dout0[127]
port 91 nsew signal input
rlabel metal2 s 21914 99200 21970 100000 6 sram_dout0[12]
port 92 nsew signal input
rlabel metal2 s 22834 99200 22890 100000 6 sram_dout0[13]
port 93 nsew signal input
rlabel metal2 s 23754 99200 23810 100000 6 sram_dout0[14]
port 94 nsew signal input
rlabel metal2 s 24674 99200 24730 100000 6 sram_dout0[15]
port 95 nsew signal input
rlabel metal2 s 25594 99200 25650 100000 6 sram_dout0[16]
port 96 nsew signal input
rlabel metal2 s 26514 99200 26570 100000 6 sram_dout0[17]
port 97 nsew signal input
rlabel metal2 s 27434 99200 27490 100000 6 sram_dout0[18]
port 98 nsew signal input
rlabel metal2 s 28446 99200 28502 100000 6 sram_dout0[19]
port 99 nsew signal input
rlabel metal2 s 5078 99200 5134 100000 6 sram_dout0[1]
port 100 nsew signal input
rlabel metal2 s 29366 99200 29422 100000 6 sram_dout0[20]
port 101 nsew signal input
rlabel metal2 s 30286 99200 30342 100000 6 sram_dout0[21]
port 102 nsew signal input
rlabel metal2 s 31206 99200 31262 100000 6 sram_dout0[22]
port 103 nsew signal input
rlabel metal2 s 32126 99200 32182 100000 6 sram_dout0[23]
port 104 nsew signal input
rlabel metal2 s 33046 99200 33102 100000 6 sram_dout0[24]
port 105 nsew signal input
rlabel metal2 s 34058 99200 34114 100000 6 sram_dout0[25]
port 106 nsew signal input
rlabel metal2 s 34978 99200 35034 100000 6 sram_dout0[26]
port 107 nsew signal input
rlabel metal2 s 35898 99200 35954 100000 6 sram_dout0[27]
port 108 nsew signal input
rlabel metal2 s 36818 99200 36874 100000 6 sram_dout0[28]
port 109 nsew signal input
rlabel metal2 s 37738 99200 37794 100000 6 sram_dout0[29]
port 110 nsew signal input
rlabel metal2 s 7562 99200 7618 100000 6 sram_dout0[2]
port 111 nsew signal input
rlabel metal2 s 38658 99200 38714 100000 6 sram_dout0[30]
port 112 nsew signal input
rlabel metal2 s 39670 99200 39726 100000 6 sram_dout0[31]
port 113 nsew signal input
rlabel metal2 s 40222 99200 40278 100000 6 sram_dout0[32]
port 114 nsew signal input
rlabel metal2 s 40866 99200 40922 100000 6 sram_dout0[33]
port 115 nsew signal input
rlabel metal2 s 41510 99200 41566 100000 6 sram_dout0[34]
port 116 nsew signal input
rlabel metal2 s 42154 99200 42210 100000 6 sram_dout0[35]
port 117 nsew signal input
rlabel metal2 s 42706 99200 42762 100000 6 sram_dout0[36]
port 118 nsew signal input
rlabel metal2 s 43350 99200 43406 100000 6 sram_dout0[37]
port 119 nsew signal input
rlabel metal2 s 43994 99200 44050 100000 6 sram_dout0[38]
port 120 nsew signal input
rlabel metal2 s 44638 99200 44694 100000 6 sram_dout0[39]
port 121 nsew signal input
rlabel metal2 s 10046 99200 10102 100000 6 sram_dout0[3]
port 122 nsew signal input
rlabel metal2 s 45282 99200 45338 100000 6 sram_dout0[40]
port 123 nsew signal input
rlabel metal2 s 45834 99200 45890 100000 6 sram_dout0[41]
port 124 nsew signal input
rlabel metal2 s 46478 99200 46534 100000 6 sram_dout0[42]
port 125 nsew signal input
rlabel metal2 s 47122 99200 47178 100000 6 sram_dout0[43]
port 126 nsew signal input
rlabel metal2 s 47766 99200 47822 100000 6 sram_dout0[44]
port 127 nsew signal input
rlabel metal2 s 48318 99200 48374 100000 6 sram_dout0[45]
port 128 nsew signal input
rlabel metal2 s 48962 99200 49018 100000 6 sram_dout0[46]
port 129 nsew signal input
rlabel metal2 s 49606 99200 49662 100000 6 sram_dout0[47]
port 130 nsew signal input
rlabel metal2 s 50250 99200 50306 100000 6 sram_dout0[48]
port 131 nsew signal input
rlabel metal2 s 50802 99200 50858 100000 6 sram_dout0[49]
port 132 nsew signal input
rlabel metal2 s 11886 99200 11942 100000 6 sram_dout0[4]
port 133 nsew signal input
rlabel metal2 s 51446 99200 51502 100000 6 sram_dout0[50]
port 134 nsew signal input
rlabel metal2 s 52090 99200 52146 100000 6 sram_dout0[51]
port 135 nsew signal input
rlabel metal2 s 52734 99200 52790 100000 6 sram_dout0[52]
port 136 nsew signal input
rlabel metal2 s 53378 99200 53434 100000 6 sram_dout0[53]
port 137 nsew signal input
rlabel metal2 s 53930 99200 53986 100000 6 sram_dout0[54]
port 138 nsew signal input
rlabel metal2 s 54574 99200 54630 100000 6 sram_dout0[55]
port 139 nsew signal input
rlabel metal2 s 55218 99200 55274 100000 6 sram_dout0[56]
port 140 nsew signal input
rlabel metal2 s 55862 99200 55918 100000 6 sram_dout0[57]
port 141 nsew signal input
rlabel metal2 s 56414 99200 56470 100000 6 sram_dout0[58]
port 142 nsew signal input
rlabel metal2 s 57058 99200 57114 100000 6 sram_dout0[59]
port 143 nsew signal input
rlabel metal2 s 13450 99200 13506 100000 6 sram_dout0[5]
port 144 nsew signal input
rlabel metal2 s 57702 99200 57758 100000 6 sram_dout0[60]
port 145 nsew signal input
rlabel metal2 s 58346 99200 58402 100000 6 sram_dout0[61]
port 146 nsew signal input
rlabel metal2 s 58990 99200 59046 100000 6 sram_dout0[62]
port 147 nsew signal input
rlabel metal2 s 59542 99200 59598 100000 6 sram_dout0[63]
port 148 nsew signal input
rlabel metal2 s 60186 99200 60242 100000 6 sram_dout0[64]
port 149 nsew signal input
rlabel metal2 s 60830 99200 60886 100000 6 sram_dout0[65]
port 150 nsew signal input
rlabel metal2 s 61474 99200 61530 100000 6 sram_dout0[66]
port 151 nsew signal input
rlabel metal2 s 62026 99200 62082 100000 6 sram_dout0[67]
port 152 nsew signal input
rlabel metal2 s 62670 99200 62726 100000 6 sram_dout0[68]
port 153 nsew signal input
rlabel metal2 s 63314 99200 63370 100000 6 sram_dout0[69]
port 154 nsew signal input
rlabel metal2 s 15014 99200 15070 100000 6 sram_dout0[6]
port 155 nsew signal input
rlabel metal2 s 63958 99200 64014 100000 6 sram_dout0[70]
port 156 nsew signal input
rlabel metal2 s 64510 99200 64566 100000 6 sram_dout0[71]
port 157 nsew signal input
rlabel metal2 s 65154 99200 65210 100000 6 sram_dout0[72]
port 158 nsew signal input
rlabel metal2 s 65798 99200 65854 100000 6 sram_dout0[73]
port 159 nsew signal input
rlabel metal2 s 66442 99200 66498 100000 6 sram_dout0[74]
port 160 nsew signal input
rlabel metal2 s 67086 99200 67142 100000 6 sram_dout0[75]
port 161 nsew signal input
rlabel metal2 s 67638 99200 67694 100000 6 sram_dout0[76]
port 162 nsew signal input
rlabel metal2 s 68282 99200 68338 100000 6 sram_dout0[77]
port 163 nsew signal input
rlabel metal2 s 68926 99200 68982 100000 6 sram_dout0[78]
port 164 nsew signal input
rlabel metal2 s 69570 99200 69626 100000 6 sram_dout0[79]
port 165 nsew signal input
rlabel metal2 s 16578 99200 16634 100000 6 sram_dout0[7]
port 166 nsew signal input
rlabel metal2 s 70122 99200 70178 100000 6 sram_dout0[80]
port 167 nsew signal input
rlabel metal2 s 70766 99200 70822 100000 6 sram_dout0[81]
port 168 nsew signal input
rlabel metal2 s 71410 99200 71466 100000 6 sram_dout0[82]
port 169 nsew signal input
rlabel metal2 s 72054 99200 72110 100000 6 sram_dout0[83]
port 170 nsew signal input
rlabel metal2 s 72698 99200 72754 100000 6 sram_dout0[84]
port 171 nsew signal input
rlabel metal2 s 73250 99200 73306 100000 6 sram_dout0[85]
port 172 nsew signal input
rlabel metal2 s 73894 99200 73950 100000 6 sram_dout0[86]
port 173 nsew signal input
rlabel metal2 s 74538 99200 74594 100000 6 sram_dout0[87]
port 174 nsew signal input
rlabel metal2 s 75182 99200 75238 100000 6 sram_dout0[88]
port 175 nsew signal input
rlabel metal2 s 75734 99200 75790 100000 6 sram_dout0[89]
port 176 nsew signal input
rlabel metal2 s 18142 99200 18198 100000 6 sram_dout0[8]
port 177 nsew signal input
rlabel metal2 s 76378 99200 76434 100000 6 sram_dout0[90]
port 178 nsew signal input
rlabel metal2 s 77022 99200 77078 100000 6 sram_dout0[91]
port 179 nsew signal input
rlabel metal2 s 77666 99200 77722 100000 6 sram_dout0[92]
port 180 nsew signal input
rlabel metal2 s 78218 99200 78274 100000 6 sram_dout0[93]
port 181 nsew signal input
rlabel metal2 s 78862 99200 78918 100000 6 sram_dout0[94]
port 182 nsew signal input
rlabel metal2 s 79506 99200 79562 100000 6 sram_dout0[95]
port 183 nsew signal input
rlabel metal2 s 80150 99200 80206 100000 6 sram_dout0[96]
port 184 nsew signal input
rlabel metal2 s 80794 99200 80850 100000 6 sram_dout0[97]
port 185 nsew signal input
rlabel metal2 s 81346 99200 81402 100000 6 sram_dout0[98]
port 186 nsew signal input
rlabel metal2 s 81990 99200 82046 100000 6 sram_dout0[99]
port 187 nsew signal input
rlabel metal2 s 19062 99200 19118 100000 6 sram_dout0[9]
port 188 nsew signal input
rlabel metal2 s 2870 99200 2926 100000 6 sram_dout1[0]
port 189 nsew signal input
rlabel metal2 s 82910 99200 82966 100000 6 sram_dout1[100]
port 190 nsew signal input
rlabel metal2 s 83554 99200 83610 100000 6 sram_dout1[101]
port 191 nsew signal input
rlabel metal2 s 84198 99200 84254 100000 6 sram_dout1[102]
port 192 nsew signal input
rlabel metal2 s 84842 99200 84898 100000 6 sram_dout1[103]
port 193 nsew signal input
rlabel metal2 s 85394 99200 85450 100000 6 sram_dout1[104]
port 194 nsew signal input
rlabel metal2 s 86038 99200 86094 100000 6 sram_dout1[105]
port 195 nsew signal input
rlabel metal2 s 86682 99200 86738 100000 6 sram_dout1[106]
port 196 nsew signal input
rlabel metal2 s 87326 99200 87382 100000 6 sram_dout1[107]
port 197 nsew signal input
rlabel metal2 s 87878 99200 87934 100000 6 sram_dout1[108]
port 198 nsew signal input
rlabel metal2 s 88522 99200 88578 100000 6 sram_dout1[109]
port 199 nsew signal input
rlabel metal2 s 20350 99200 20406 100000 6 sram_dout1[10]
port 200 nsew signal input
rlabel metal2 s 89166 99200 89222 100000 6 sram_dout1[110]
port 201 nsew signal input
rlabel metal2 s 89810 99200 89866 100000 6 sram_dout1[111]
port 202 nsew signal input
rlabel metal2 s 90454 99200 90510 100000 6 sram_dout1[112]
port 203 nsew signal input
rlabel metal2 s 91006 99200 91062 100000 6 sram_dout1[113]
port 204 nsew signal input
rlabel metal2 s 91650 99200 91706 100000 6 sram_dout1[114]
port 205 nsew signal input
rlabel metal2 s 92294 99200 92350 100000 6 sram_dout1[115]
port 206 nsew signal input
rlabel metal2 s 92938 99200 92994 100000 6 sram_dout1[116]
port 207 nsew signal input
rlabel metal2 s 93490 99200 93546 100000 6 sram_dout1[117]
port 208 nsew signal input
rlabel metal2 s 94134 99200 94190 100000 6 sram_dout1[118]
port 209 nsew signal input
rlabel metal2 s 94778 99200 94834 100000 6 sram_dout1[119]
port 210 nsew signal input
rlabel metal2 s 21270 99200 21326 100000 6 sram_dout1[11]
port 211 nsew signal input
rlabel metal2 s 95422 99200 95478 100000 6 sram_dout1[120]
port 212 nsew signal input
rlabel metal2 s 95974 99200 96030 100000 6 sram_dout1[121]
port 213 nsew signal input
rlabel metal2 s 96618 99200 96674 100000 6 sram_dout1[122]
port 214 nsew signal input
rlabel metal2 s 97262 99200 97318 100000 6 sram_dout1[123]
port 215 nsew signal input
rlabel metal2 s 97906 99200 97962 100000 6 sram_dout1[124]
port 216 nsew signal input
rlabel metal2 s 98550 99200 98606 100000 6 sram_dout1[125]
port 217 nsew signal input
rlabel metal2 s 99102 99200 99158 100000 6 sram_dout1[126]
port 218 nsew signal input
rlabel metal2 s 99746 99200 99802 100000 6 sram_dout1[127]
port 219 nsew signal input
rlabel metal2 s 22190 99200 22246 100000 6 sram_dout1[12]
port 220 nsew signal input
rlabel metal2 s 23110 99200 23166 100000 6 sram_dout1[13]
port 221 nsew signal input
rlabel metal2 s 24030 99200 24086 100000 6 sram_dout1[14]
port 222 nsew signal input
rlabel metal2 s 24950 99200 25006 100000 6 sram_dout1[15]
port 223 nsew signal input
rlabel metal2 s 25962 99200 26018 100000 6 sram_dout1[16]
port 224 nsew signal input
rlabel metal2 s 26882 99200 26938 100000 6 sram_dout1[17]
port 225 nsew signal input
rlabel metal2 s 27802 99200 27858 100000 6 sram_dout1[18]
port 226 nsew signal input
rlabel metal2 s 28722 99200 28778 100000 6 sram_dout1[19]
port 227 nsew signal input
rlabel metal2 s 5354 99200 5410 100000 6 sram_dout1[1]
port 228 nsew signal input
rlabel metal2 s 29642 99200 29698 100000 6 sram_dout1[20]
port 229 nsew signal input
rlabel metal2 s 30562 99200 30618 100000 6 sram_dout1[21]
port 230 nsew signal input
rlabel metal2 s 31574 99200 31630 100000 6 sram_dout1[22]
port 231 nsew signal input
rlabel metal2 s 32494 99200 32550 100000 6 sram_dout1[23]
port 232 nsew signal input
rlabel metal2 s 33414 99200 33470 100000 6 sram_dout1[24]
port 233 nsew signal input
rlabel metal2 s 34334 99200 34390 100000 6 sram_dout1[25]
port 234 nsew signal input
rlabel metal2 s 35254 99200 35310 100000 6 sram_dout1[26]
port 235 nsew signal input
rlabel metal2 s 36174 99200 36230 100000 6 sram_dout1[27]
port 236 nsew signal input
rlabel metal2 s 37094 99200 37150 100000 6 sram_dout1[28]
port 237 nsew signal input
rlabel metal2 s 38106 99200 38162 100000 6 sram_dout1[29]
port 238 nsew signal input
rlabel metal2 s 7838 99200 7894 100000 6 sram_dout1[2]
port 239 nsew signal input
rlabel metal2 s 39026 99200 39082 100000 6 sram_dout1[30]
port 240 nsew signal input
rlabel metal2 s 39946 99200 40002 100000 6 sram_dout1[31]
port 241 nsew signal input
rlabel metal2 s 40590 99200 40646 100000 6 sram_dout1[32]
port 242 nsew signal input
rlabel metal2 s 41142 99200 41198 100000 6 sram_dout1[33]
port 243 nsew signal input
rlabel metal2 s 41786 99200 41842 100000 6 sram_dout1[34]
port 244 nsew signal input
rlabel metal2 s 42430 99200 42486 100000 6 sram_dout1[35]
port 245 nsew signal input
rlabel metal2 s 43074 99200 43130 100000 6 sram_dout1[36]
port 246 nsew signal input
rlabel metal2 s 43718 99200 43774 100000 6 sram_dout1[37]
port 247 nsew signal input
rlabel metal2 s 44270 99200 44326 100000 6 sram_dout1[38]
port 248 nsew signal input
rlabel metal2 s 44914 99200 44970 100000 6 sram_dout1[39]
port 249 nsew signal input
rlabel metal2 s 10322 99200 10378 100000 6 sram_dout1[3]
port 250 nsew signal input
rlabel metal2 s 45558 99200 45614 100000 6 sram_dout1[40]
port 251 nsew signal input
rlabel metal2 s 46202 99200 46258 100000 6 sram_dout1[41]
port 252 nsew signal input
rlabel metal2 s 46754 99200 46810 100000 6 sram_dout1[42]
port 253 nsew signal input
rlabel metal2 s 47398 99200 47454 100000 6 sram_dout1[43]
port 254 nsew signal input
rlabel metal2 s 48042 99200 48098 100000 6 sram_dout1[44]
port 255 nsew signal input
rlabel metal2 s 48686 99200 48742 100000 6 sram_dout1[45]
port 256 nsew signal input
rlabel metal2 s 49330 99200 49386 100000 6 sram_dout1[46]
port 257 nsew signal input
rlabel metal2 s 49882 99200 49938 100000 6 sram_dout1[47]
port 258 nsew signal input
rlabel metal2 s 50526 99200 50582 100000 6 sram_dout1[48]
port 259 nsew signal input
rlabel metal2 s 51170 99200 51226 100000 6 sram_dout1[49]
port 260 nsew signal input
rlabel metal2 s 12254 99200 12310 100000 6 sram_dout1[4]
port 261 nsew signal input
rlabel metal2 s 51814 99200 51870 100000 6 sram_dout1[50]
port 262 nsew signal input
rlabel metal2 s 52366 99200 52422 100000 6 sram_dout1[51]
port 263 nsew signal input
rlabel metal2 s 53010 99200 53066 100000 6 sram_dout1[52]
port 264 nsew signal input
rlabel metal2 s 53654 99200 53710 100000 6 sram_dout1[53]
port 265 nsew signal input
rlabel metal2 s 54298 99200 54354 100000 6 sram_dout1[54]
port 266 nsew signal input
rlabel metal2 s 54850 99200 54906 100000 6 sram_dout1[55]
port 267 nsew signal input
rlabel metal2 s 55494 99200 55550 100000 6 sram_dout1[56]
port 268 nsew signal input
rlabel metal2 s 56138 99200 56194 100000 6 sram_dout1[57]
port 269 nsew signal input
rlabel metal2 s 56782 99200 56838 100000 6 sram_dout1[58]
port 270 nsew signal input
rlabel metal2 s 57426 99200 57482 100000 6 sram_dout1[59]
port 271 nsew signal input
rlabel metal2 s 13726 99200 13782 100000 6 sram_dout1[5]
port 272 nsew signal input
rlabel metal2 s 57978 99200 58034 100000 6 sram_dout1[60]
port 273 nsew signal input
rlabel metal2 s 58622 99200 58678 100000 6 sram_dout1[61]
port 274 nsew signal input
rlabel metal2 s 59266 99200 59322 100000 6 sram_dout1[62]
port 275 nsew signal input
rlabel metal2 s 59910 99200 59966 100000 6 sram_dout1[63]
port 276 nsew signal input
rlabel metal2 s 60462 99200 60518 100000 6 sram_dout1[64]
port 277 nsew signal input
rlabel metal2 s 61106 99200 61162 100000 6 sram_dout1[65]
port 278 nsew signal input
rlabel metal2 s 61750 99200 61806 100000 6 sram_dout1[66]
port 279 nsew signal input
rlabel metal2 s 62394 99200 62450 100000 6 sram_dout1[67]
port 280 nsew signal input
rlabel metal2 s 63038 99200 63094 100000 6 sram_dout1[68]
port 281 nsew signal input
rlabel metal2 s 63590 99200 63646 100000 6 sram_dout1[69]
port 282 nsew signal input
rlabel metal2 s 15290 99200 15346 100000 6 sram_dout1[6]
port 283 nsew signal input
rlabel metal2 s 64234 99200 64290 100000 6 sram_dout1[70]
port 284 nsew signal input
rlabel metal2 s 64878 99200 64934 100000 6 sram_dout1[71]
port 285 nsew signal input
rlabel metal2 s 65522 99200 65578 100000 6 sram_dout1[72]
port 286 nsew signal input
rlabel metal2 s 66074 99200 66130 100000 6 sram_dout1[73]
port 287 nsew signal input
rlabel metal2 s 66718 99200 66774 100000 6 sram_dout1[74]
port 288 nsew signal input
rlabel metal2 s 67362 99200 67418 100000 6 sram_dout1[75]
port 289 nsew signal input
rlabel metal2 s 68006 99200 68062 100000 6 sram_dout1[76]
port 290 nsew signal input
rlabel metal2 s 68558 99200 68614 100000 6 sram_dout1[77]
port 291 nsew signal input
rlabel metal2 s 69202 99200 69258 100000 6 sram_dout1[78]
port 292 nsew signal input
rlabel metal2 s 69846 99200 69902 100000 6 sram_dout1[79]
port 293 nsew signal input
rlabel metal2 s 16854 99200 16910 100000 6 sram_dout1[7]
port 294 nsew signal input
rlabel metal2 s 70490 99200 70546 100000 6 sram_dout1[80]
port 295 nsew signal input
rlabel metal2 s 71134 99200 71190 100000 6 sram_dout1[81]
port 296 nsew signal input
rlabel metal2 s 71686 99200 71742 100000 6 sram_dout1[82]
port 297 nsew signal input
rlabel metal2 s 72330 99200 72386 100000 6 sram_dout1[83]
port 298 nsew signal input
rlabel metal2 s 72974 99200 73030 100000 6 sram_dout1[84]
port 299 nsew signal input
rlabel metal2 s 73618 99200 73674 100000 6 sram_dout1[85]
port 300 nsew signal input
rlabel metal2 s 74170 99200 74226 100000 6 sram_dout1[86]
port 301 nsew signal input
rlabel metal2 s 74814 99200 74870 100000 6 sram_dout1[87]
port 302 nsew signal input
rlabel metal2 s 75458 99200 75514 100000 6 sram_dout1[88]
port 303 nsew signal input
rlabel metal2 s 76102 99200 76158 100000 6 sram_dout1[89]
port 304 nsew signal input
rlabel metal2 s 18418 99200 18474 100000 6 sram_dout1[8]
port 305 nsew signal input
rlabel metal2 s 76746 99200 76802 100000 6 sram_dout1[90]
port 306 nsew signal input
rlabel metal2 s 77298 99200 77354 100000 6 sram_dout1[91]
port 307 nsew signal input
rlabel metal2 s 77942 99200 77998 100000 6 sram_dout1[92]
port 308 nsew signal input
rlabel metal2 s 78586 99200 78642 100000 6 sram_dout1[93]
port 309 nsew signal input
rlabel metal2 s 79230 99200 79286 100000 6 sram_dout1[94]
port 310 nsew signal input
rlabel metal2 s 79782 99200 79838 100000 6 sram_dout1[95]
port 311 nsew signal input
rlabel metal2 s 80426 99200 80482 100000 6 sram_dout1[96]
port 312 nsew signal input
rlabel metal2 s 81070 99200 81126 100000 6 sram_dout1[97]
port 313 nsew signal input
rlabel metal2 s 81714 99200 81770 100000 6 sram_dout1[98]
port 314 nsew signal input
rlabel metal2 s 82266 99200 82322 100000 6 sram_dout1[99]
port 315 nsew signal input
rlabel metal2 s 19338 99200 19394 100000 6 sram_dout1[9]
port 316 nsew signal input
rlabel metal2 s 662 99200 718 100000 6 sram_web0
port 317 nsew signal output
rlabel metal2 s 3146 99200 3202 100000 6 sram_wmask0[0]
port 318 nsew signal output
rlabel metal2 s 5630 99200 5686 100000 6 sram_wmask0[1]
port 319 nsew signal output
rlabel metal2 s 8206 99200 8262 100000 6 sram_wmask0[2]
port 320 nsew signal output
rlabel metal2 s 10690 99200 10746 100000 6 sram_wmask0[3]
port 321 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 322 nsew power bidirectional
rlabel metal3 s 99200 31016 100000 31136 6 vga_b[0]
port 323 nsew signal output
rlabel metal3 s 99200 68552 100000 68672 6 vga_b[1]
port 324 nsew signal output
rlabel metal3 s 99200 43528 100000 43648 6 vga_g[0]
port 325 nsew signal output
rlabel metal3 s 99200 81064 100000 81184 6 vga_g[1]
port 326 nsew signal output
rlabel metal3 s 99200 6128 100000 6248 6 vga_hsync
port 327 nsew signal output
rlabel metal3 s 99200 56040 100000 56160 6 vga_r[0]
port 328 nsew signal output
rlabel metal3 s 99200 93576 100000 93696 6 vga_r[1]
port 329 nsew signal output
rlabel metal3 s 99200 18504 100000 18624 6 vga_vsync
port 330 nsew signal output
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 331 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 331 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 331 nsew ground bidirectional
rlabel metal2 s 478 0 534 800 6 wb_ack_o
port 332 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wb_adr_i[0]
port 333 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wb_adr_i[10]
port 334 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wb_adr_i[11]
port 335 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wb_adr_i[12]
port 336 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 wb_adr_i[13]
port 337 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wb_adr_i[14]
port 338 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wb_adr_i[15]
port 339 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wb_adr_i[16]
port 340 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wb_adr_i[17]
port 341 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wb_adr_i[18]
port 342 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wb_adr_i[19]
port 343 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wb_adr_i[1]
port 344 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 wb_adr_i[20]
port 345 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 wb_adr_i[21]
port 346 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 wb_adr_i[22]
port 347 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 wb_adr_i[23]
port 348 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wb_adr_i[2]
port 349 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wb_adr_i[3]
port 350 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wb_adr_i[4]
port 351 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wb_adr_i[5]
port 352 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wb_adr_i[6]
port 353 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wb_adr_i[7]
port 354 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wb_adr_i[8]
port 355 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wb_adr_i[9]
port 356 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_clk_i
port 357 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wb_cyc_i
port 358 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wb_data_i[0]
port 359 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wb_data_i[10]
port 360 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wb_data_i[11]
port 361 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wb_data_i[12]
port 362 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wb_data_i[13]
port 363 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wb_data_i[14]
port 364 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wb_data_i[15]
port 365 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wb_data_i[16]
port 366 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wb_data_i[17]
port 367 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wb_data_i[18]
port 368 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wb_data_i[19]
port 369 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wb_data_i[1]
port 370 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 wb_data_i[20]
port 371 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 wb_data_i[21]
port 372 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 wb_data_i[22]
port 373 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wb_data_i[23]
port 374 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 wb_data_i[24]
port 375 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 wb_data_i[25]
port 376 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 wb_data_i[26]
port 377 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 wb_data_i[27]
port 378 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wb_data_i[28]
port 379 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 wb_data_i[29]
port 380 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wb_data_i[2]
port 381 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 wb_data_i[30]
port 382 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 wb_data_i[31]
port 383 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wb_data_i[3]
port 384 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wb_data_i[4]
port 385 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wb_data_i[5]
port 386 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wb_data_i[6]
port 387 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wb_data_i[7]
port 388 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wb_data_i[8]
port 389 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wb_data_i[9]
port 390 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wb_data_o[0]
port 391 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 wb_data_o[10]
port 392 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 wb_data_o[11]
port 393 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 wb_data_o[12]
port 394 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 wb_data_o[13]
port 395 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 wb_data_o[14]
port 396 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 wb_data_o[15]
port 397 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 wb_data_o[16]
port 398 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 wb_data_o[17]
port 399 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 wb_data_o[18]
port 400 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 wb_data_o[19]
port 401 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wb_data_o[1]
port 402 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 wb_data_o[20]
port 403 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 wb_data_o[21]
port 404 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 wb_data_o[22]
port 405 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 wb_data_o[23]
port 406 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 wb_data_o[24]
port 407 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wb_data_o[25]
port 408 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 wb_data_o[26]
port 409 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 wb_data_o[27]
port 410 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 wb_data_o[28]
port 411 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 wb_data_o[29]
port 412 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wb_data_o[2]
port 413 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 wb_data_o[30]
port 414 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 wb_data_o[31]
port 415 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wb_data_o[3]
port 416 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wb_data_o[4]
port 417 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wb_data_o[5]
port 418 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wb_data_o[6]
port 419 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wb_data_o[7]
port 420 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wb_data_o[8]
port 421 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wb_data_o[9]
port 422 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 wb_error_o
port 423 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wb_rst_i
port 424 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wb_sel_i[0]
port 425 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wb_sel_i[1]
port 426 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wb_sel_i[2]
port 427 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wb_sel_i[3]
port 428 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wb_stall_o
port 429 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wb_stb_i
port 430 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wb_we_i
port 431 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7552660
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Video/runs/Video/results/signoff/Video.magic.gds
string GDS_START 694590
<< end >>

