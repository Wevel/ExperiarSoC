VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WishboneInterconnect
  CLASS BLOCK ;
  FOREIGN WishboneInterconnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 1100.000 ;
  PIN master0_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END master0_wb_ack_i
  PIN master0_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END master0_wb_adr_o[0]
  PIN master0_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END master0_wb_adr_o[10]
  PIN master0_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END master0_wb_adr_o[11]
  PIN master0_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END master0_wb_adr_o[12]
  PIN master0_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END master0_wb_adr_o[13]
  PIN master0_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END master0_wb_adr_o[14]
  PIN master0_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END master0_wb_adr_o[15]
  PIN master0_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END master0_wb_adr_o[16]
  PIN master0_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END master0_wb_adr_o[17]
  PIN master0_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END master0_wb_adr_o[18]
  PIN master0_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END master0_wb_adr_o[19]
  PIN master0_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END master0_wb_adr_o[1]
  PIN master0_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END master0_wb_adr_o[20]
  PIN master0_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END master0_wb_adr_o[21]
  PIN master0_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END master0_wb_adr_o[22]
  PIN master0_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END master0_wb_adr_o[23]
  PIN master0_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END master0_wb_adr_o[24]
  PIN master0_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END master0_wb_adr_o[25]
  PIN master0_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END master0_wb_adr_o[26]
  PIN master0_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END master0_wb_adr_o[27]
  PIN master0_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END master0_wb_adr_o[2]
  PIN master0_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END master0_wb_adr_o[3]
  PIN master0_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END master0_wb_adr_o[4]
  PIN master0_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END master0_wb_adr_o[5]
  PIN master0_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END master0_wb_adr_o[6]
  PIN master0_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END master0_wb_adr_o[7]
  PIN master0_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END master0_wb_adr_o[8]
  PIN master0_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END master0_wb_adr_o[9]
  PIN master0_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END master0_wb_cyc_o
  PIN master0_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END master0_wb_data_i[0]
  PIN master0_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END master0_wb_data_i[10]
  PIN master0_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END master0_wb_data_i[11]
  PIN master0_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END master0_wb_data_i[12]
  PIN master0_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END master0_wb_data_i[13]
  PIN master0_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END master0_wb_data_i[14]
  PIN master0_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END master0_wb_data_i[15]
  PIN master0_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END master0_wb_data_i[16]
  PIN master0_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END master0_wb_data_i[17]
  PIN master0_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END master0_wb_data_i[18]
  PIN master0_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END master0_wb_data_i[19]
  PIN master0_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END master0_wb_data_i[1]
  PIN master0_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END master0_wb_data_i[20]
  PIN master0_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END master0_wb_data_i[21]
  PIN master0_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END master0_wb_data_i[22]
  PIN master0_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END master0_wb_data_i[23]
  PIN master0_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END master0_wb_data_i[24]
  PIN master0_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END master0_wb_data_i[25]
  PIN master0_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END master0_wb_data_i[26]
  PIN master0_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END master0_wb_data_i[27]
  PIN master0_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END master0_wb_data_i[28]
  PIN master0_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END master0_wb_data_i[29]
  PIN master0_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END master0_wb_data_i[2]
  PIN master0_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END master0_wb_data_i[30]
  PIN master0_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END master0_wb_data_i[31]
  PIN master0_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END master0_wb_data_i[3]
  PIN master0_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END master0_wb_data_i[4]
  PIN master0_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END master0_wb_data_i[5]
  PIN master0_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END master0_wb_data_i[6]
  PIN master0_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END master0_wb_data_i[7]
  PIN master0_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END master0_wb_data_i[8]
  PIN master0_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END master0_wb_data_i[9]
  PIN master0_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END master0_wb_data_o[0]
  PIN master0_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END master0_wb_data_o[10]
  PIN master0_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END master0_wb_data_o[11]
  PIN master0_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END master0_wb_data_o[12]
  PIN master0_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END master0_wb_data_o[13]
  PIN master0_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END master0_wb_data_o[14]
  PIN master0_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END master0_wb_data_o[15]
  PIN master0_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END master0_wb_data_o[16]
  PIN master0_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END master0_wb_data_o[17]
  PIN master0_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END master0_wb_data_o[18]
  PIN master0_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END master0_wb_data_o[19]
  PIN master0_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END master0_wb_data_o[1]
  PIN master0_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END master0_wb_data_o[20]
  PIN master0_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END master0_wb_data_o[21]
  PIN master0_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END master0_wb_data_o[22]
  PIN master0_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END master0_wb_data_o[23]
  PIN master0_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END master0_wb_data_o[24]
  PIN master0_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END master0_wb_data_o[25]
  PIN master0_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END master0_wb_data_o[26]
  PIN master0_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END master0_wb_data_o[27]
  PIN master0_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END master0_wb_data_o[28]
  PIN master0_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END master0_wb_data_o[29]
  PIN master0_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END master0_wb_data_o[2]
  PIN master0_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END master0_wb_data_o[30]
  PIN master0_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END master0_wb_data_o[31]
  PIN master0_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END master0_wb_data_o[3]
  PIN master0_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END master0_wb_data_o[4]
  PIN master0_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END master0_wb_data_o[5]
  PIN master0_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END master0_wb_data_o[6]
  PIN master0_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END master0_wb_data_o[7]
  PIN master0_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END master0_wb_data_o[8]
  PIN master0_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END master0_wb_data_o[9]
  PIN master0_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END master0_wb_error_i
  PIN master0_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END master0_wb_sel_o[0]
  PIN master0_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END master0_wb_sel_o[1]
  PIN master0_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END master0_wb_sel_o[2]
  PIN master0_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END master0_wb_sel_o[3]
  PIN master0_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END master0_wb_stall_i
  PIN master0_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END master0_wb_stb_o
  PIN master0_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END master0_wb_we_o
  PIN master1_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 551.520 4.000 552.120 ;
    END
  END master1_wb_ack_i
  PIN master1_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END master1_wb_adr_o[0]
  PIN master1_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END master1_wb_adr_o[10]
  PIN master1_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END master1_wb_adr_o[11]
  PIN master1_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END master1_wb_adr_o[12]
  PIN master1_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END master1_wb_adr_o[13]
  PIN master1_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 694.320 4.000 694.920 ;
    END
  END master1_wb_adr_o[14]
  PIN master1_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END master1_wb_adr_o[15]
  PIN master1_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END master1_wb_adr_o[16]
  PIN master1_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.800 4.000 719.400 ;
    END
  END master1_wb_adr_o[17]
  PIN master1_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END master1_wb_adr_o[18]
  PIN master1_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END master1_wb_adr_o[19]
  PIN master1_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END master1_wb_adr_o[1]
  PIN master1_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END master1_wb_adr_o[20]
  PIN master1_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END master1_wb_adr_o[21]
  PIN master1_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END master1_wb_adr_o[22]
  PIN master1_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END master1_wb_adr_o[23]
  PIN master1_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END master1_wb_adr_o[24]
  PIN master1_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END master1_wb_adr_o[25]
  PIN master1_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END master1_wb_adr_o[26]
  PIN master1_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END master1_wb_adr_o[27]
  PIN master1_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END master1_wb_adr_o[2]
  PIN master1_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 600.480 4.000 601.080 ;
    END
  END master1_wb_adr_o[3]
  PIN master1_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 611.360 4.000 611.960 ;
    END
  END master1_wb_adr_o[4]
  PIN master1_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END master1_wb_adr_o[5]
  PIN master1_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END master1_wb_adr_o[6]
  PIN master1_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END master1_wb_adr_o[7]
  PIN master1_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END master1_wb_adr_o[8]
  PIN master1_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END master1_wb_adr_o[9]
  PIN master1_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END master1_wb_cyc_o
  PIN master1_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END master1_wb_data_i[0]
  PIN master1_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END master1_wb_data_i[10]
  PIN master1_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END master1_wb_data_i[11]
  PIN master1_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END master1_wb_data_i[12]
  PIN master1_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END master1_wb_data_i[13]
  PIN master1_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END master1_wb_data_i[14]
  PIN master1_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END master1_wb_data_i[15]
  PIN master1_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END master1_wb_data_i[16]
  PIN master1_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END master1_wb_data_i[17]
  PIN master1_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END master1_wb_data_i[18]
  PIN master1_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END master1_wb_data_i[19]
  PIN master1_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END master1_wb_data_i[1]
  PIN master1_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END master1_wb_data_i[20]
  PIN master1_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END master1_wb_data_i[21]
  PIN master1_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END master1_wb_data_i[22]
  PIN master1_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END master1_wb_data_i[23]
  PIN master1_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END master1_wb_data_i[24]
  PIN master1_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END master1_wb_data_i[25]
  PIN master1_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 796.320 4.000 796.920 ;
    END
  END master1_wb_data_i[26]
  PIN master1_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 804.480 4.000 805.080 ;
    END
  END master1_wb_data_i[27]
  PIN master1_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.920 4.000 810.520 ;
    END
  END master1_wb_data_i[28]
  PIN master1_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END master1_wb_data_i[29]
  PIN master1_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END master1_wb_data_i[2]
  PIN master1_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END master1_wb_data_i[30]
  PIN master1_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END master1_wb_data_i[31]
  PIN master1_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END master1_wb_data_i[3]
  PIN master1_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END master1_wb_data_i[4]
  PIN master1_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END master1_wb_data_i[5]
  PIN master1_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END master1_wb_data_i[6]
  PIN master1_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END master1_wb_data_i[7]
  PIN master1_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END master1_wb_data_i[8]
  PIN master1_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END master1_wb_data_i[9]
  PIN master1_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END master1_wb_data_o[0]
  PIN master1_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END master1_wb_data_o[10]
  PIN master1_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END master1_wb_data_o[11]
  PIN master1_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END master1_wb_data_o[12]
  PIN master1_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END master1_wb_data_o[13]
  PIN master1_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.760 4.000 700.360 ;
    END
  END master1_wb_data_o[14]
  PIN master1_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.920 4.000 708.520 ;
    END
  END master1_wb_data_o[15]
  PIN master1_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END master1_wb_data_o[16]
  PIN master1_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END master1_wb_data_o[17]
  PIN master1_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 732.400 4.000 733.000 ;
    END
  END master1_wb_data_o[18]
  PIN master1_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END master1_wb_data_o[19]
  PIN master1_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.160 4.000 584.760 ;
    END
  END master1_wb_data_o[1]
  PIN master1_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END master1_wb_data_o[20]
  PIN master1_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END master1_wb_data_o[21]
  PIN master1_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END master1_wb_data_o[22]
  PIN master1_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END master1_wb_data_o[23]
  PIN master1_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END master1_wb_data_o[24]
  PIN master1_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.200 4.000 790.800 ;
    END
  END master1_wb_data_o[25]
  PIN master1_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END master1_wb_data_o[26]
  PIN master1_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END master1_wb_data_o[27]
  PIN master1_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END master1_wb_data_o[28]
  PIN master1_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END master1_wb_data_o[29]
  PIN master1_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END master1_wb_data_o[2]
  PIN master1_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END master1_wb_data_o[30]
  PIN master1_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.960 4.000 829.560 ;
    END
  END master1_wb_data_o[31]
  PIN master1_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END master1_wb_data_o[3]
  PIN master1_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END master1_wb_data_o[4]
  PIN master1_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END master1_wb_data_o[5]
  PIN master1_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END master1_wb_data_o[6]
  PIN master1_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END master1_wb_data_o[7]
  PIN master1_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END master1_wb_data_o[8]
  PIN master1_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END master1_wb_data_o[9]
  PIN master1_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END master1_wb_error_i
  PIN master1_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.000 4.000 576.600 ;
    END
  END master1_wb_sel_o[0]
  PIN master1_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END master1_wb_sel_o[1]
  PIN master1_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END master1_wb_sel_o[2]
  PIN master1_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END master1_wb_sel_o[3]
  PIN master1_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END master1_wb_stall_i
  PIN master1_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END master1_wb_stb_o
  PIN master1_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.120 4.000 565.720 ;
    END
  END master1_wb_we_o
  PIN master2_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END master2_wb_ack_i
  PIN master2_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END master2_wb_adr_o[0]
  PIN master2_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END master2_wb_adr_o[10]
  PIN master2_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END master2_wb_adr_o[11]
  PIN master2_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END master2_wb_adr_o[12]
  PIN master2_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END master2_wb_adr_o[13]
  PIN master2_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END master2_wb_adr_o[14]
  PIN master2_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END master2_wb_adr_o[15]
  PIN master2_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END master2_wb_adr_o[16]
  PIN master2_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END master2_wb_adr_o[17]
  PIN master2_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END master2_wb_adr_o[18]
  PIN master2_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END master2_wb_adr_o[19]
  PIN master2_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END master2_wb_adr_o[1]
  PIN master2_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END master2_wb_adr_o[20]
  PIN master2_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END master2_wb_adr_o[21]
  PIN master2_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END master2_wb_adr_o[22]
  PIN master2_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END master2_wb_adr_o[23]
  PIN master2_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END master2_wb_adr_o[24]
  PIN master2_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END master2_wb_adr_o[25]
  PIN master2_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END master2_wb_adr_o[26]
  PIN master2_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END master2_wb_adr_o[27]
  PIN master2_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END master2_wb_adr_o[2]
  PIN master2_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END master2_wb_adr_o[3]
  PIN master2_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END master2_wb_adr_o[4]
  PIN master2_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END master2_wb_adr_o[5]
  PIN master2_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END master2_wb_adr_o[6]
  PIN master2_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END master2_wb_adr_o[7]
  PIN master2_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END master2_wb_adr_o[8]
  PIN master2_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END master2_wb_adr_o[9]
  PIN master2_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END master2_wb_cyc_o
  PIN master2_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END master2_wb_data_i[0]
  PIN master2_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END master2_wb_data_i[10]
  PIN master2_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END master2_wb_data_i[11]
  PIN master2_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END master2_wb_data_i[12]
  PIN master2_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END master2_wb_data_i[13]
  PIN master2_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END master2_wb_data_i[14]
  PIN master2_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END master2_wb_data_i[15]
  PIN master2_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END master2_wb_data_i[16]
  PIN master2_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END master2_wb_data_i[17]
  PIN master2_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END master2_wb_data_i[18]
  PIN master2_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END master2_wb_data_i[19]
  PIN master2_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END master2_wb_data_i[1]
  PIN master2_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END master2_wb_data_i[20]
  PIN master2_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END master2_wb_data_i[21]
  PIN master2_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END master2_wb_data_i[22]
  PIN master2_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END master2_wb_data_i[23]
  PIN master2_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END master2_wb_data_i[24]
  PIN master2_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END master2_wb_data_i[25]
  PIN master2_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END master2_wb_data_i[26]
  PIN master2_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END master2_wb_data_i[27]
  PIN master2_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END master2_wb_data_i[28]
  PIN master2_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END master2_wb_data_i[29]
  PIN master2_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END master2_wb_data_i[2]
  PIN master2_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END master2_wb_data_i[30]
  PIN master2_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END master2_wb_data_i[31]
  PIN master2_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END master2_wb_data_i[3]
  PIN master2_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END master2_wb_data_i[4]
  PIN master2_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END master2_wb_data_i[5]
  PIN master2_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END master2_wb_data_i[6]
  PIN master2_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END master2_wb_data_i[7]
  PIN master2_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END master2_wb_data_i[8]
  PIN master2_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END master2_wb_data_i[9]
  PIN master2_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END master2_wb_data_o[0]
  PIN master2_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END master2_wb_data_o[10]
  PIN master2_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END master2_wb_data_o[11]
  PIN master2_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END master2_wb_data_o[12]
  PIN master2_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END master2_wb_data_o[13]
  PIN master2_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END master2_wb_data_o[14]
  PIN master2_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END master2_wb_data_o[15]
  PIN master2_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END master2_wb_data_o[16]
  PIN master2_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END master2_wb_data_o[17]
  PIN master2_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END master2_wb_data_o[18]
  PIN master2_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END master2_wb_data_o[19]
  PIN master2_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END master2_wb_data_o[1]
  PIN master2_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END master2_wb_data_o[20]
  PIN master2_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END master2_wb_data_o[21]
  PIN master2_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END master2_wb_data_o[22]
  PIN master2_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END master2_wb_data_o[23]
  PIN master2_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END master2_wb_data_o[24]
  PIN master2_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END master2_wb_data_o[25]
  PIN master2_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END master2_wb_data_o[26]
  PIN master2_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END master2_wb_data_o[27]
  PIN master2_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END master2_wb_data_o[28]
  PIN master2_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END master2_wb_data_o[29]
  PIN master2_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END master2_wb_data_o[2]
  PIN master2_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END master2_wb_data_o[30]
  PIN master2_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END master2_wb_data_o[31]
  PIN master2_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END master2_wb_data_o[3]
  PIN master2_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END master2_wb_data_o[4]
  PIN master2_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END master2_wb_data_o[5]
  PIN master2_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END master2_wb_data_o[6]
  PIN master2_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END master2_wb_data_o[7]
  PIN master2_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END master2_wb_data_o[8]
  PIN master2_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END master2_wb_data_o[9]
  PIN master2_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END master2_wb_error_i
  PIN master2_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END master2_wb_sel_o[0]
  PIN master2_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END master2_wb_sel_o[1]
  PIN master2_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END master2_wb_sel_o[2]
  PIN master2_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END master2_wb_sel_o[3]
  PIN master2_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END master2_wb_stall_i
  PIN master2_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END master2_wb_stb_o
  PIN master2_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END master2_wb_we_o
  PIN probe_master0_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END probe_master0_currentSlave[0]
  PIN probe_master0_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END probe_master0_currentSlave[1]
  PIN probe_master1_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END probe_master1_currentSlave[0]
  PIN probe_master1_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END probe_master1_currentSlave[1]
  PIN probe_master2_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END probe_master2_currentSlave[0]
  PIN probe_master2_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END probe_master2_currentSlave[1]
  PIN probe_master3_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END probe_master3_currentSlave[0]
  PIN probe_master3_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END probe_master3_currentSlave[1]
  PIN probe_slave0_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END probe_slave0_currentMaster[0]
  PIN probe_slave0_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END probe_slave0_currentMaster[1]
  PIN probe_slave1_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END probe_slave1_currentMaster[0]
  PIN probe_slave1_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END probe_slave1_currentMaster[1]
  PIN probe_slave2_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END probe_slave2_currentMaster[0]
  PIN probe_slave2_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END probe_slave2_currentMaster[1]
  PIN probe_slave3_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END probe_slave3_currentMaster[0]
  PIN probe_slave3_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END probe_slave3_currentMaster[1]
  PIN slave0_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.680 4.000 832.280 ;
    END
  END slave0_wb_ack_o
  PIN slave0_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.000 4.000 848.600 ;
    END
  END slave0_wb_adr_i[0]
  PIN slave0_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END slave0_wb_adr_i[10]
  PIN slave0_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.000 4.000 950.600 ;
    END
  END slave0_wb_adr_i[11]
  PIN slave0_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.160 4.000 958.760 ;
    END
  END slave0_wb_adr_i[12]
  PIN slave0_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 966.320 4.000 966.920 ;
    END
  END slave0_wb_adr_i[13]
  PIN slave0_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END slave0_wb_adr_i[14]
  PIN slave0_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END slave0_wb_adr_i[15]
  PIN slave0_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END slave0_wb_adr_i[16]
  PIN slave0_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END slave0_wb_adr_i[17]
  PIN slave0_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END slave0_wb_adr_i[18]
  PIN slave0_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.960 4.000 1016.560 ;
    END
  END slave0_wb_adr_i[19]
  PIN slave0_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END slave0_wb_adr_i[1]
  PIN slave0_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END slave0_wb_adr_i[20]
  PIN slave0_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END slave0_wb_adr_i[21]
  PIN slave0_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.120 4.000 1041.720 ;
    END
  END slave0_wb_adr_i[22]
  PIN slave0_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END slave0_wb_adr_i[23]
  PIN slave0_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END slave0_wb_adr_i[2]
  PIN slave0_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END slave0_wb_adr_i[3]
  PIN slave0_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END slave0_wb_adr_i[4]
  PIN slave0_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 4.000 900.960 ;
    END
  END slave0_wb_adr_i[5]
  PIN slave0_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END slave0_wb_adr_i[6]
  PIN slave0_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END slave0_wb_adr_i[7]
  PIN slave0_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END slave0_wb_adr_i[8]
  PIN slave0_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.680 4.000 934.280 ;
    END
  END slave0_wb_adr_i[9]
  PIN slave0_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 834.400 4.000 835.000 ;
    END
  END slave0_wb_cyc_i
  PIN slave0_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.720 4.000 851.320 ;
    END
  END slave0_wb_data_i[0]
  PIN slave0_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END slave0_wb_data_i[10]
  PIN slave0_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.720 4.000 953.320 ;
    END
  END slave0_wb_data_i[11]
  PIN slave0_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END slave0_wb_data_i[12]
  PIN slave0_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END slave0_wb_data_i[13]
  PIN slave0_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.200 4.000 977.800 ;
    END
  END slave0_wb_data_i[14]
  PIN slave0_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END slave0_wb_data_i[15]
  PIN slave0_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END slave0_wb_data_i[16]
  PIN slave0_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1002.360 4.000 1002.960 ;
    END
  END slave0_wb_data_i[17]
  PIN slave0_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1010.520 4.000 1011.120 ;
    END
  END slave0_wb_data_i[18]
  PIN slave0_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END slave0_wb_data_i[19]
  PIN slave0_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END slave0_wb_data_i[1]
  PIN slave0_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END slave0_wb_data_i[20]
  PIN slave0_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.000 4.000 1035.600 ;
    END
  END slave0_wb_data_i[21]
  PIN slave0_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END slave0_wb_data_i[22]
  PIN slave0_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1052.000 4.000 1052.600 ;
    END
  END slave0_wb_data_i[23]
  PIN slave0_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END slave0_wb_data_i[24]
  PIN slave0_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.880 4.000 1063.480 ;
    END
  END slave0_wb_data_i[25]
  PIN slave0_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1068.320 4.000 1068.920 ;
    END
  END slave0_wb_data_i[26]
  PIN slave0_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.760 4.000 1074.360 ;
    END
  END slave0_wb_data_i[27]
  PIN slave0_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.200 4.000 1079.800 ;
    END
  END slave0_wb_data_i[28]
  PIN slave0_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END slave0_wb_data_i[29]
  PIN slave0_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END slave0_wb_data_i[2]
  PIN slave0_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.080 4.000 1090.680 ;
    END
  END slave0_wb_data_i[30]
  PIN slave0_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1095.520 4.000 1096.120 ;
    END
  END slave0_wb_data_i[31]
  PIN slave0_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END slave0_wb_data_i[3]
  PIN slave0_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END slave0_wb_data_i[4]
  PIN slave0_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.080 4.000 903.680 ;
    END
  END slave0_wb_data_i[5]
  PIN slave0_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END slave0_wb_data_i[6]
  PIN slave0_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END slave0_wb_data_i[7]
  PIN slave0_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END slave0_wb_data_i[8]
  PIN slave0_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 936.400 4.000 937.000 ;
    END
  END slave0_wb_data_i[9]
  PIN slave0_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END slave0_wb_data_o[0]
  PIN slave0_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.280 4.000 947.880 ;
    END
  END slave0_wb_data_o[10]
  PIN slave0_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END slave0_wb_data_o[11]
  PIN slave0_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END slave0_wb_data_o[12]
  PIN slave0_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.760 4.000 972.360 ;
    END
  END slave0_wb_data_o[13]
  PIN slave0_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END slave0_wb_data_o[14]
  PIN slave0_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.760 4.000 989.360 ;
    END
  END slave0_wb_data_o[15]
  PIN slave0_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END slave0_wb_data_o[16]
  PIN slave0_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.080 4.000 1005.680 ;
    END
  END slave0_wb_data_o[17]
  PIN slave0_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END slave0_wb_data_o[18]
  PIN slave0_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1021.400 4.000 1022.000 ;
    END
  END slave0_wb_data_o[19]
  PIN slave0_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END slave0_wb_data_o[1]
  PIN slave0_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END slave0_wb_data_o[20]
  PIN slave0_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.720 4.000 1038.320 ;
    END
  END slave0_wb_data_o[21]
  PIN slave0_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END slave0_wb_data_o[22]
  PIN slave0_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.720 4.000 1055.320 ;
    END
  END slave0_wb_data_o[23]
  PIN slave0_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.160 4.000 1060.760 ;
    END
  END slave0_wb_data_o[24]
  PIN slave0_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1065.600 4.000 1066.200 ;
    END
  END slave0_wb_data_o[25]
  PIN slave0_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END slave0_wb_data_o[26]
  PIN slave0_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1076.480 4.000 1077.080 ;
    END
  END slave0_wb_data_o[27]
  PIN slave0_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.920 4.000 1082.520 ;
    END
  END slave0_wb_data_o[28]
  PIN slave0_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1087.360 4.000 1087.960 ;
    END
  END slave0_wb_data_o[29]
  PIN slave0_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END slave0_wb_data_o[2]
  PIN slave0_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1092.800 4.000 1093.400 ;
    END
  END slave0_wb_data_o[30]
  PIN slave0_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END slave0_wb_data_o[31]
  PIN slave0_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.760 4.000 887.360 ;
    END
  END slave0_wb_data_o[3]
  PIN slave0_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END slave0_wb_data_o[4]
  PIN slave0_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END slave0_wb_data_o[5]
  PIN slave0_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.960 4.000 914.560 ;
    END
  END slave0_wb_data_o[6]
  PIN slave0_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.800 4.000 923.400 ;
    END
  END slave0_wb_data_o[7]
  PIN slave0_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END slave0_wb_data_o[8]
  PIN slave0_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END slave0_wb_data_o[9]
  PIN slave0_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.120 4.000 837.720 ;
    END
  END slave0_wb_error_o
  PIN slave0_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.160 4.000 856.760 ;
    END
  END slave0_wb_sel_i[0]
  PIN slave0_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END slave0_wb_sel_i[1]
  PIN slave0_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END slave0_wb_sel_i[2]
  PIN slave0_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END slave0_wb_sel_i[3]
  PIN slave0_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END slave0_wb_stall_o
  PIN slave0_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 842.560 4.000 843.160 ;
    END
  END slave0_wb_stb_i
  PIN slave0_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.280 4.000 845.880 ;
    END
  END slave0_wb_we_i
  PIN slave1_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END slave1_wb_ack_o
  PIN slave1_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END slave1_wb_adr_i[0]
  PIN slave1_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END slave1_wb_adr_i[10]
  PIN slave1_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END slave1_wb_adr_i[11]
  PIN slave1_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END slave1_wb_adr_i[12]
  PIN slave1_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END slave1_wb_adr_i[13]
  PIN slave1_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END slave1_wb_adr_i[14]
  PIN slave1_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END slave1_wb_adr_i[15]
  PIN slave1_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END slave1_wb_adr_i[16]
  PIN slave1_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END slave1_wb_adr_i[17]
  PIN slave1_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END slave1_wb_adr_i[18]
  PIN slave1_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END slave1_wb_adr_i[19]
  PIN slave1_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END slave1_wb_adr_i[1]
  PIN slave1_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END slave1_wb_adr_i[20]
  PIN slave1_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END slave1_wb_adr_i[21]
  PIN slave1_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END slave1_wb_adr_i[22]
  PIN slave1_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END slave1_wb_adr_i[23]
  PIN slave1_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END slave1_wb_adr_i[2]
  PIN slave1_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END slave1_wb_adr_i[3]
  PIN slave1_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END slave1_wb_adr_i[4]
  PIN slave1_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END slave1_wb_adr_i[5]
  PIN slave1_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END slave1_wb_adr_i[6]
  PIN slave1_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END slave1_wb_adr_i[7]
  PIN slave1_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END slave1_wb_adr_i[8]
  PIN slave1_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END slave1_wb_adr_i[9]
  PIN slave1_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END slave1_wb_cyc_i
  PIN slave1_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END slave1_wb_data_i[0]
  PIN slave1_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END slave1_wb_data_i[10]
  PIN slave1_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END slave1_wb_data_i[11]
  PIN slave1_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END slave1_wb_data_i[12]
  PIN slave1_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END slave1_wb_data_i[13]
  PIN slave1_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END slave1_wb_data_i[14]
  PIN slave1_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END slave1_wb_data_i[15]
  PIN slave1_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END slave1_wb_data_i[16]
  PIN slave1_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END slave1_wb_data_i[17]
  PIN slave1_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END slave1_wb_data_i[18]
  PIN slave1_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END slave1_wb_data_i[19]
  PIN slave1_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END slave1_wb_data_i[1]
  PIN slave1_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END slave1_wb_data_i[20]
  PIN slave1_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END slave1_wb_data_i[21]
  PIN slave1_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END slave1_wb_data_i[22]
  PIN slave1_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END slave1_wb_data_i[23]
  PIN slave1_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END slave1_wb_data_i[24]
  PIN slave1_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END slave1_wb_data_i[25]
  PIN slave1_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END slave1_wb_data_i[26]
  PIN slave1_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END slave1_wb_data_i[27]
  PIN slave1_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END slave1_wb_data_i[28]
  PIN slave1_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END slave1_wb_data_i[29]
  PIN slave1_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END slave1_wb_data_i[2]
  PIN slave1_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END slave1_wb_data_i[30]
  PIN slave1_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END slave1_wb_data_i[31]
  PIN slave1_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END slave1_wb_data_i[3]
  PIN slave1_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END slave1_wb_data_i[4]
  PIN slave1_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END slave1_wb_data_i[5]
  PIN slave1_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END slave1_wb_data_i[6]
  PIN slave1_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END slave1_wb_data_i[7]
  PIN slave1_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END slave1_wb_data_i[8]
  PIN slave1_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END slave1_wb_data_i[9]
  PIN slave1_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END slave1_wb_data_o[0]
  PIN slave1_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END slave1_wb_data_o[10]
  PIN slave1_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END slave1_wb_data_o[11]
  PIN slave1_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END slave1_wb_data_o[12]
  PIN slave1_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END slave1_wb_data_o[13]
  PIN slave1_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END slave1_wb_data_o[14]
  PIN slave1_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END slave1_wb_data_o[15]
  PIN slave1_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END slave1_wb_data_o[16]
  PIN slave1_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END slave1_wb_data_o[17]
  PIN slave1_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END slave1_wb_data_o[18]
  PIN slave1_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END slave1_wb_data_o[19]
  PIN slave1_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END slave1_wb_data_o[1]
  PIN slave1_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END slave1_wb_data_o[20]
  PIN slave1_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END slave1_wb_data_o[21]
  PIN slave1_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END slave1_wb_data_o[22]
  PIN slave1_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END slave1_wb_data_o[23]
  PIN slave1_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END slave1_wb_data_o[24]
  PIN slave1_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END slave1_wb_data_o[25]
  PIN slave1_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END slave1_wb_data_o[26]
  PIN slave1_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END slave1_wb_data_o[27]
  PIN slave1_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END slave1_wb_data_o[28]
  PIN slave1_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END slave1_wb_data_o[29]
  PIN slave1_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END slave1_wb_data_o[2]
  PIN slave1_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END slave1_wb_data_o[30]
  PIN slave1_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END slave1_wb_data_o[31]
  PIN slave1_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END slave1_wb_data_o[3]
  PIN slave1_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END slave1_wb_data_o[4]
  PIN slave1_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END slave1_wb_data_o[5]
  PIN slave1_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END slave1_wb_data_o[6]
  PIN slave1_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END slave1_wb_data_o[7]
  PIN slave1_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END slave1_wb_data_o[8]
  PIN slave1_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END slave1_wb_data_o[9]
  PIN slave1_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END slave1_wb_error_o
  PIN slave1_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END slave1_wb_sel_i[0]
  PIN slave1_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END slave1_wb_sel_i[1]
  PIN slave1_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END slave1_wb_sel_i[2]
  PIN slave1_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END slave1_wb_sel_i[3]
  PIN slave1_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END slave1_wb_stall_o
  PIN slave1_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END slave1_wb_stb_i
  PIN slave1_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END slave1_wb_we_i
  PIN slave2_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 1096.000 1.750 1100.000 ;
    END
  END slave2_wb_ack_o
  PIN slave2_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1096.000 22.910 1100.000 ;
    END
  END slave2_wb_adr_i[0]
  PIN slave2_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 1096.000 144.350 1100.000 ;
    END
  END slave2_wb_adr_i[10]
  PIN slave2_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1096.000 154.930 1100.000 ;
    END
  END slave2_wb_adr_i[11]
  PIN slave2_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 1096.000 165.970 1100.000 ;
    END
  END slave2_wb_adr_i[12]
  PIN slave2_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 1096.000 176.550 1100.000 ;
    END
  END slave2_wb_adr_i[13]
  PIN slave2_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 1096.000 187.130 1100.000 ;
    END
  END slave2_wb_adr_i[14]
  PIN slave2_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 1096.000 198.170 1100.000 ;
    END
  END slave2_wb_adr_i[15]
  PIN slave2_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 1096.000 208.750 1100.000 ;
    END
  END slave2_wb_adr_i[16]
  PIN slave2_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1096.000 219.330 1100.000 ;
    END
  END slave2_wb_adr_i[17]
  PIN slave2_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 1096.000 229.910 1100.000 ;
    END
  END slave2_wb_adr_i[18]
  PIN slave2_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 1096.000 240.950 1100.000 ;
    END
  END slave2_wb_adr_i[19]
  PIN slave2_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 1096.000 37.170 1100.000 ;
    END
  END slave2_wb_adr_i[1]
  PIN slave2_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1096.000 251.530 1100.000 ;
    END
  END slave2_wb_adr_i[20]
  PIN slave2_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 1096.000 262.110 1100.000 ;
    END
  END slave2_wb_adr_i[21]
  PIN slave2_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 1096.000 273.150 1100.000 ;
    END
  END slave2_wb_adr_i[22]
  PIN slave2_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1096.000 283.730 1100.000 ;
    END
  END slave2_wb_adr_i[23]
  PIN slave2_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 1096.000 51.430 1100.000 ;
    END
  END slave2_wb_adr_i[2]
  PIN slave2_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 1096.000 65.690 1100.000 ;
    END
  END slave2_wb_adr_i[3]
  PIN slave2_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 1096.000 79.950 1100.000 ;
    END
  END slave2_wb_adr_i[4]
  PIN slave2_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 1096.000 90.990 1100.000 ;
    END
  END slave2_wb_adr_i[5]
  PIN slave2_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 1096.000 101.570 1100.000 ;
    END
  END slave2_wb_adr_i[6]
  PIN slave2_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 1096.000 112.150 1100.000 ;
    END
  END slave2_wb_adr_i[7]
  PIN slave2_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 1096.000 123.190 1100.000 ;
    END
  END slave2_wb_adr_i[8]
  PIN slave2_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 1096.000 133.770 1100.000 ;
    END
  END slave2_wb_adr_i[9]
  PIN slave2_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 1096.000 4.970 1100.000 ;
    END
  END slave2_wb_cyc_i
  PIN slave2_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 1096.000 26.590 1100.000 ;
    END
  END slave2_wb_data_i[0]
  PIN slave2_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 1096.000 148.030 1100.000 ;
    END
  END slave2_wb_data_i[10]
  PIN slave2_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 1096.000 158.610 1100.000 ;
    END
  END slave2_wb_data_i[11]
  PIN slave2_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 1096.000 169.190 1100.000 ;
    END
  END slave2_wb_data_i[12]
  PIN slave2_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 1096.000 180.230 1100.000 ;
    END
  END slave2_wb_data_i[13]
  PIN slave2_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 1096.000 190.810 1100.000 ;
    END
  END slave2_wb_data_i[14]
  PIN slave2_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 1096.000 201.390 1100.000 ;
    END
  END slave2_wb_data_i[15]
  PIN slave2_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 1096.000 212.430 1100.000 ;
    END
  END slave2_wb_data_i[16]
  PIN slave2_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 1096.000 223.010 1100.000 ;
    END
  END slave2_wb_data_i[17]
  PIN slave2_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 1096.000 233.590 1100.000 ;
    END
  END slave2_wb_data_i[18]
  PIN slave2_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 1096.000 244.630 1100.000 ;
    END
  END slave2_wb_data_i[19]
  PIN slave2_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 1096.000 40.850 1100.000 ;
    END
  END slave2_wb_data_i[1]
  PIN slave2_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 1096.000 255.210 1100.000 ;
    END
  END slave2_wb_data_i[20]
  PIN slave2_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 1096.000 265.790 1100.000 ;
    END
  END slave2_wb_data_i[21]
  PIN slave2_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 1096.000 276.370 1100.000 ;
    END
  END slave2_wb_data_i[22]
  PIN slave2_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 1096.000 287.410 1100.000 ;
    END
  END slave2_wb_data_i[23]
  PIN slave2_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 1096.000 294.310 1100.000 ;
    END
  END slave2_wb_data_i[24]
  PIN slave2_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 1096.000 301.670 1100.000 ;
    END
  END slave2_wb_data_i[25]
  PIN slave2_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 1096.000 308.570 1100.000 ;
    END
  END slave2_wb_data_i[26]
  PIN slave2_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1096.000 315.930 1100.000 ;
    END
  END slave2_wb_data_i[27]
  PIN slave2_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 1096.000 322.830 1100.000 ;
    END
  END slave2_wb_data_i[28]
  PIN slave2_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 1096.000 330.190 1100.000 ;
    END
  END slave2_wb_data_i[29]
  PIN slave2_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1096.000 55.110 1100.000 ;
    END
  END slave2_wb_data_i[2]
  PIN slave2_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 1096.000 337.090 1100.000 ;
    END
  END slave2_wb_data_i[30]
  PIN slave2_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 1096.000 344.450 1100.000 ;
    END
  END slave2_wb_data_i[31]
  PIN slave2_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 1096.000 69.370 1100.000 ;
    END
  END slave2_wb_data_i[3]
  PIN slave2_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 1096.000 83.630 1100.000 ;
    END
  END slave2_wb_data_i[4]
  PIN slave2_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 1096.000 94.210 1100.000 ;
    END
  END slave2_wb_data_i[5]
  PIN slave2_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 1096.000 105.250 1100.000 ;
    END
  END slave2_wb_data_i[6]
  PIN slave2_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 1096.000 115.830 1100.000 ;
    END
  END slave2_wb_data_i[7]
  PIN slave2_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 1096.000 126.410 1100.000 ;
    END
  END slave2_wb_data_i[8]
  PIN slave2_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 1096.000 137.450 1100.000 ;
    END
  END slave2_wb_data_i[9]
  PIN slave2_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 1096.000 30.270 1100.000 ;
    END
  END slave2_wb_data_o[0]
  PIN slave2_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1096.000 151.710 1100.000 ;
    END
  END slave2_wb_data_o[10]
  PIN slave2_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 1096.000 162.290 1100.000 ;
    END
  END slave2_wb_data_o[11]
  PIN slave2_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 1096.000 172.870 1100.000 ;
    END
  END slave2_wb_data_o[12]
  PIN slave2_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1096.000 183.910 1100.000 ;
    END
  END slave2_wb_data_o[13]
  PIN slave2_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 1096.000 194.490 1100.000 ;
    END
  END slave2_wb_data_o[14]
  PIN slave2_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 1096.000 205.070 1100.000 ;
    END
  END slave2_wb_data_o[15]
  PIN slave2_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 1096.000 215.650 1100.000 ;
    END
  END slave2_wb_data_o[16]
  PIN slave2_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 1096.000 226.690 1100.000 ;
    END
  END slave2_wb_data_o[17]
  PIN slave2_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 1096.000 237.270 1100.000 ;
    END
  END slave2_wb_data_o[18]
  PIN slave2_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 1096.000 247.850 1100.000 ;
    END
  END slave2_wb_data_o[19]
  PIN slave2_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 1096.000 44.530 1100.000 ;
    END
  END slave2_wb_data_o[1]
  PIN slave2_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 1096.000 258.890 1100.000 ;
    END
  END slave2_wb_data_o[20]
  PIN slave2_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 1096.000 269.470 1100.000 ;
    END
  END slave2_wb_data_o[21]
  PIN slave2_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 1096.000 280.050 1100.000 ;
    END
  END slave2_wb_data_o[22]
  PIN slave2_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 1096.000 290.630 1100.000 ;
    END
  END slave2_wb_data_o[23]
  PIN slave2_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 1096.000 297.990 1100.000 ;
    END
  END slave2_wb_data_o[24]
  PIN slave2_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 1096.000 305.350 1100.000 ;
    END
  END slave2_wb_data_o[25]
  PIN slave2_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 1096.000 312.250 1100.000 ;
    END
  END slave2_wb_data_o[26]
  PIN slave2_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 1096.000 319.610 1100.000 ;
    END
  END slave2_wb_data_o[27]
  PIN slave2_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 1096.000 326.510 1100.000 ;
    END
  END slave2_wb_data_o[28]
  PIN slave2_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 1096.000 333.870 1100.000 ;
    END
  END slave2_wb_data_o[29]
  PIN slave2_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 1096.000 58.790 1100.000 ;
    END
  END slave2_wb_data_o[2]
  PIN slave2_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 1096.000 340.770 1100.000 ;
    END
  END slave2_wb_data_o[30]
  PIN slave2_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 1096.000 348.130 1100.000 ;
    END
  END slave2_wb_data_o[31]
  PIN slave2_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 1096.000 73.050 1100.000 ;
    END
  END slave2_wb_data_o[3]
  PIN slave2_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1096.000 87.310 1100.000 ;
    END
  END slave2_wb_data_o[4]
  PIN slave2_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 1096.000 97.890 1100.000 ;
    END
  END slave2_wb_data_o[5]
  PIN slave2_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 1096.000 108.470 1100.000 ;
    END
  END slave2_wb_data_o[6]
  PIN slave2_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1096.000 119.510 1100.000 ;
    END
  END slave2_wb_data_o[7]
  PIN slave2_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 1096.000 130.090 1100.000 ;
    END
  END slave2_wb_data_o[8]
  PIN slave2_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 1096.000 140.670 1100.000 ;
    END
  END slave2_wb_data_o[9]
  PIN slave2_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 1096.000 8.650 1100.000 ;
    END
  END slave2_wb_error_o
  PIN slave2_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 1096.000 33.490 1100.000 ;
    END
  END slave2_wb_sel_i[0]
  PIN slave2_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1096.000 47.750 1100.000 ;
    END
  END slave2_wb_sel_i[1]
  PIN slave2_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 1096.000 62.470 1100.000 ;
    END
  END slave2_wb_sel_i[2]
  PIN slave2_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 1096.000 76.730 1100.000 ;
    END
  END slave2_wb_sel_i[3]
  PIN slave2_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 1096.000 12.330 1100.000 ;
    END
  END slave2_wb_stall_o
  PIN slave2_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 1096.000 16.010 1100.000 ;
    END
  END slave2_wb_stb_i
  PIN slave2_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 1096.000 19.230 1100.000 ;
    END
  END slave2_wb_we_i
  PIN slave3_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 552.880 350.000 553.480 ;
    END
  END slave3_wb_ack_o
  PIN slave3_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 586.200 350.000 586.800 ;
    END
  END slave3_wb_adr_i[0]
  PIN slave3_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 777.280 350.000 777.880 ;
    END
  END slave3_wb_adr_i[10]
  PIN slave3_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 793.600 350.000 794.200 ;
    END
  END slave3_wb_adr_i[11]
  PIN slave3_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 810.600 350.000 811.200 ;
    END
  END slave3_wb_adr_i[12]
  PIN slave3_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 827.600 350.000 828.200 ;
    END
  END slave3_wb_adr_i[13]
  PIN slave3_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 844.600 350.000 845.200 ;
    END
  END slave3_wb_adr_i[14]
  PIN slave3_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 861.600 350.000 862.200 ;
    END
  END slave3_wb_adr_i[15]
  PIN slave3_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 877.920 350.000 878.520 ;
    END
  END slave3_wb_adr_i[16]
  PIN slave3_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 894.920 350.000 895.520 ;
    END
  END slave3_wb_adr_i[17]
  PIN slave3_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 911.920 350.000 912.520 ;
    END
  END slave3_wb_adr_i[18]
  PIN slave3_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 928.920 350.000 929.520 ;
    END
  END slave3_wb_adr_i[19]
  PIN slave3_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 608.640 350.000 609.240 ;
    END
  END slave3_wb_adr_i[1]
  PIN slave3_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 945.240 350.000 945.840 ;
    END
  END slave3_wb_adr_i[20]
  PIN slave3_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 962.240 350.000 962.840 ;
    END
  END slave3_wb_adr_i[21]
  PIN slave3_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 979.240 350.000 979.840 ;
    END
  END slave3_wb_adr_i[22]
  PIN slave3_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 996.240 350.000 996.840 ;
    END
  END slave3_wb_adr_i[23]
  PIN slave3_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 631.080 350.000 631.680 ;
    END
  END slave3_wb_adr_i[2]
  PIN slave3_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 653.520 350.000 654.120 ;
    END
  END slave3_wb_adr_i[3]
  PIN slave3_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 675.960 350.000 676.560 ;
    END
  END slave3_wb_adr_i[4]
  PIN slave3_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 692.960 350.000 693.560 ;
    END
  END slave3_wb_adr_i[5]
  PIN slave3_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 709.960 350.000 710.560 ;
    END
  END slave3_wb_adr_i[6]
  PIN slave3_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 726.280 350.000 726.880 ;
    END
  END slave3_wb_adr_i[7]
  PIN slave3_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 743.280 350.000 743.880 ;
    END
  END slave3_wb_adr_i[8]
  PIN slave3_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 760.280 350.000 760.880 ;
    END
  END slave3_wb_adr_i[9]
  PIN slave3_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 558.320 350.000 558.920 ;
    END
  END slave3_wb_cyc_i
  PIN slave3_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 591.640 350.000 592.240 ;
    END
  END slave3_wb_data_i[0]
  PIN slave3_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 782.720 350.000 783.320 ;
    END
  END slave3_wb_data_i[10]
  PIN slave3_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 799.720 350.000 800.320 ;
    END
  END slave3_wb_data_i[11]
  PIN slave3_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 816.040 350.000 816.640 ;
    END
  END slave3_wb_data_i[12]
  PIN slave3_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 833.040 350.000 833.640 ;
    END
  END slave3_wb_data_i[13]
  PIN slave3_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 850.040 350.000 850.640 ;
    END
  END slave3_wb_data_i[14]
  PIN slave3_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 867.040 350.000 867.640 ;
    END
  END slave3_wb_data_i[15]
  PIN slave3_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 884.040 350.000 884.640 ;
    END
  END slave3_wb_data_i[16]
  PIN slave3_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 900.360 350.000 900.960 ;
    END
  END slave3_wb_data_i[17]
  PIN slave3_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 917.360 350.000 917.960 ;
    END
  END slave3_wb_data_i[18]
  PIN slave3_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 934.360 350.000 934.960 ;
    END
  END slave3_wb_data_i[19]
  PIN slave3_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 614.080 350.000 614.680 ;
    END
  END slave3_wb_data_i[1]
  PIN slave3_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 951.360 350.000 951.960 ;
    END
  END slave3_wb_data_i[20]
  PIN slave3_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 967.680 350.000 968.280 ;
    END
  END slave3_wb_data_i[21]
  PIN slave3_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 984.680 350.000 985.280 ;
    END
  END slave3_wb_data_i[22]
  PIN slave3_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1001.680 350.000 1002.280 ;
    END
  END slave3_wb_data_i[23]
  PIN slave3_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1012.560 350.000 1013.160 ;
    END
  END slave3_wb_data_i[24]
  PIN slave3_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1024.120 350.000 1024.720 ;
    END
  END slave3_wb_data_i[25]
  PIN slave3_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1035.000 350.000 1035.600 ;
    END
  END slave3_wb_data_i[26]
  PIN slave3_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1046.560 350.000 1047.160 ;
    END
  END slave3_wb_data_i[27]
  PIN slave3_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1057.440 350.000 1058.040 ;
    END
  END slave3_wb_data_i[28]
  PIN slave3_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1069.000 350.000 1069.600 ;
    END
  END slave3_wb_data_i[29]
  PIN slave3_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 636.520 350.000 637.120 ;
    END
  END slave3_wb_data_i[2]
  PIN slave3_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1079.880 350.000 1080.480 ;
    END
  END slave3_wb_data_i[30]
  PIN slave3_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1091.440 350.000 1092.040 ;
    END
  END slave3_wb_data_i[31]
  PIN slave3_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 658.960 350.000 659.560 ;
    END
  END slave3_wb_data_i[3]
  PIN slave3_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 681.400 350.000 682.000 ;
    END
  END slave3_wb_data_i[4]
  PIN slave3_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 698.400 350.000 699.000 ;
    END
  END slave3_wb_data_i[5]
  PIN slave3_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 715.400 350.000 716.000 ;
    END
  END slave3_wb_data_i[6]
  PIN slave3_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 732.400 350.000 733.000 ;
    END
  END slave3_wb_data_i[7]
  PIN slave3_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 748.720 350.000 749.320 ;
    END
  END slave3_wb_data_i[8]
  PIN slave3_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 765.720 350.000 766.320 ;
    END
  END slave3_wb_data_i[9]
  PIN slave3_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 597.760 350.000 598.360 ;
    END
  END slave3_wb_data_o[0]
  PIN slave3_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 788.160 350.000 788.760 ;
    END
  END slave3_wb_data_o[10]
  PIN slave3_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 805.160 350.000 805.760 ;
    END
  END slave3_wb_data_o[11]
  PIN slave3_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 822.160 350.000 822.760 ;
    END
  END slave3_wb_data_o[12]
  PIN slave3_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 839.160 350.000 839.760 ;
    END
  END slave3_wb_data_o[13]
  PIN slave3_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 855.480 350.000 856.080 ;
    END
  END slave3_wb_data_o[14]
  PIN slave3_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 872.480 350.000 873.080 ;
    END
  END slave3_wb_data_o[15]
  PIN slave3_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 889.480 350.000 890.080 ;
    END
  END slave3_wb_data_o[16]
  PIN slave3_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 906.480 350.000 907.080 ;
    END
  END slave3_wb_data_o[17]
  PIN slave3_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 922.800 350.000 923.400 ;
    END
  END slave3_wb_data_o[18]
  PIN slave3_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 939.800 350.000 940.400 ;
    END
  END slave3_wb_data_o[19]
  PIN slave3_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 620.200 350.000 620.800 ;
    END
  END slave3_wb_data_o[1]
  PIN slave3_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 956.800 350.000 957.400 ;
    END
  END slave3_wb_data_o[20]
  PIN slave3_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 973.800 350.000 974.400 ;
    END
  END slave3_wb_data_o[21]
  PIN slave3_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 990.120 350.000 990.720 ;
    END
  END slave3_wb_data_o[22]
  PIN slave3_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1007.120 350.000 1007.720 ;
    END
  END slave3_wb_data_o[23]
  PIN slave3_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1018.680 350.000 1019.280 ;
    END
  END slave3_wb_data_o[24]
  PIN slave3_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1029.560 350.000 1030.160 ;
    END
  END slave3_wb_data_o[25]
  PIN slave3_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1041.120 350.000 1041.720 ;
    END
  END slave3_wb_data_o[26]
  PIN slave3_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1052.000 350.000 1052.600 ;
    END
  END slave3_wb_data_o[27]
  PIN slave3_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1063.560 350.000 1064.160 ;
    END
  END slave3_wb_data_o[28]
  PIN slave3_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1074.440 350.000 1075.040 ;
    END
  END slave3_wb_data_o[29]
  PIN slave3_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 642.640 350.000 643.240 ;
    END
  END slave3_wb_data_o[2]
  PIN slave3_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1086.000 350.000 1086.600 ;
    END
  END slave3_wb_data_o[30]
  PIN slave3_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1096.880 350.000 1097.480 ;
    END
  END slave3_wb_data_o[31]
  PIN slave3_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 665.080 350.000 665.680 ;
    END
  END slave3_wb_data_o[3]
  PIN slave3_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 687.520 350.000 688.120 ;
    END
  END slave3_wb_data_o[4]
  PIN slave3_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 703.840 350.000 704.440 ;
    END
  END slave3_wb_data_o[5]
  PIN slave3_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 720.840 350.000 721.440 ;
    END
  END slave3_wb_data_o[6]
  PIN slave3_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 737.840 350.000 738.440 ;
    END
  END slave3_wb_data_o[7]
  PIN slave3_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 754.840 350.000 755.440 ;
    END
  END slave3_wb_data_o[8]
  PIN slave3_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 771.160 350.000 771.760 ;
    END
  END slave3_wb_data_o[9]
  PIN slave3_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 563.760 350.000 564.360 ;
    END
  END slave3_wb_error_o
  PIN slave3_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 603.200 350.000 603.800 ;
    END
  END slave3_wb_sel_i[0]
  PIN slave3_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 625.640 350.000 626.240 ;
    END
  END slave3_wb_sel_i[1]
  PIN slave3_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 648.080 350.000 648.680 ;
    END
  END slave3_wb_sel_i[2]
  PIN slave3_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 670.520 350.000 671.120 ;
    END
  END slave3_wb_sel_i[3]
  PIN slave3_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 569.200 350.000 569.800 ;
    END
  END slave3_wb_stall_o
  PIN slave3_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 575.320 350.000 575.920 ;
    END
  END slave3_wb_stb_i
  PIN slave3_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 580.760 350.000 581.360 ;
    END
  END slave3_wb_we_i
  PIN slave4_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 2.760 350.000 3.360 ;
    END
  END slave4_wb_ack_o
  PIN slave4_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 36.080 350.000 36.680 ;
    END
  END slave4_wb_adr_i[0]
  PIN slave4_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 227.160 350.000 227.760 ;
    END
  END slave4_wb_adr_i[10]
  PIN slave4_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 243.480 350.000 244.080 ;
    END
  END slave4_wb_adr_i[11]
  PIN slave4_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 260.480 350.000 261.080 ;
    END
  END slave4_wb_adr_i[12]
  PIN slave4_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 277.480 350.000 278.080 ;
    END
  END slave4_wb_adr_i[13]
  PIN slave4_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 294.480 350.000 295.080 ;
    END
  END slave4_wb_adr_i[14]
  PIN slave4_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 311.480 350.000 312.080 ;
    END
  END slave4_wb_adr_i[15]
  PIN slave4_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 327.800 350.000 328.400 ;
    END
  END slave4_wb_adr_i[16]
  PIN slave4_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 344.800 350.000 345.400 ;
    END
  END slave4_wb_adr_i[17]
  PIN slave4_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 361.800 350.000 362.400 ;
    END
  END slave4_wb_adr_i[18]
  PIN slave4_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 378.800 350.000 379.400 ;
    END
  END slave4_wb_adr_i[19]
  PIN slave4_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 58.520 350.000 59.120 ;
    END
  END slave4_wb_adr_i[1]
  PIN slave4_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 395.120 350.000 395.720 ;
    END
  END slave4_wb_adr_i[20]
  PIN slave4_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 412.120 350.000 412.720 ;
    END
  END slave4_wb_adr_i[21]
  PIN slave4_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 429.120 350.000 429.720 ;
    END
  END slave4_wb_adr_i[22]
  PIN slave4_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 446.120 350.000 446.720 ;
    END
  END slave4_wb_adr_i[23]
  PIN slave4_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 80.960 350.000 81.560 ;
    END
  END slave4_wb_adr_i[2]
  PIN slave4_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 103.400 350.000 104.000 ;
    END
  END slave4_wb_adr_i[3]
  PIN slave4_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 125.840 350.000 126.440 ;
    END
  END slave4_wb_adr_i[4]
  PIN slave4_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 142.840 350.000 143.440 ;
    END
  END slave4_wb_adr_i[5]
  PIN slave4_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 159.840 350.000 160.440 ;
    END
  END slave4_wb_adr_i[6]
  PIN slave4_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 176.160 350.000 176.760 ;
    END
  END slave4_wb_adr_i[7]
  PIN slave4_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 193.160 350.000 193.760 ;
    END
  END slave4_wb_adr_i[8]
  PIN slave4_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 210.160 350.000 210.760 ;
    END
  END slave4_wb_adr_i[9]
  PIN slave4_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 8.200 350.000 8.800 ;
    END
  END slave4_wb_cyc_i
  PIN slave4_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 41.520 350.000 42.120 ;
    END
  END slave4_wb_data_i[0]
  PIN slave4_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 232.600 350.000 233.200 ;
    END
  END slave4_wb_data_i[10]
  PIN slave4_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 249.600 350.000 250.200 ;
    END
  END slave4_wb_data_i[11]
  PIN slave4_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 265.920 350.000 266.520 ;
    END
  END slave4_wb_data_i[12]
  PIN slave4_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 282.920 350.000 283.520 ;
    END
  END slave4_wb_data_i[13]
  PIN slave4_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 299.920 350.000 300.520 ;
    END
  END slave4_wb_data_i[14]
  PIN slave4_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 316.920 350.000 317.520 ;
    END
  END slave4_wb_data_i[15]
  PIN slave4_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 333.920 350.000 334.520 ;
    END
  END slave4_wb_data_i[16]
  PIN slave4_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 350.240 350.000 350.840 ;
    END
  END slave4_wb_data_i[17]
  PIN slave4_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 367.240 350.000 367.840 ;
    END
  END slave4_wb_data_i[18]
  PIN slave4_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 384.240 350.000 384.840 ;
    END
  END slave4_wb_data_i[19]
  PIN slave4_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 63.960 350.000 64.560 ;
    END
  END slave4_wb_data_i[1]
  PIN slave4_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 401.240 350.000 401.840 ;
    END
  END slave4_wb_data_i[20]
  PIN slave4_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 417.560 350.000 418.160 ;
    END
  END slave4_wb_data_i[21]
  PIN slave4_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 434.560 350.000 435.160 ;
    END
  END slave4_wb_data_i[22]
  PIN slave4_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 451.560 350.000 452.160 ;
    END
  END slave4_wb_data_i[23]
  PIN slave4_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 462.440 350.000 463.040 ;
    END
  END slave4_wb_data_i[24]
  PIN slave4_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 474.000 350.000 474.600 ;
    END
  END slave4_wb_data_i[25]
  PIN slave4_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 484.880 350.000 485.480 ;
    END
  END slave4_wb_data_i[26]
  PIN slave4_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 496.440 350.000 497.040 ;
    END
  END slave4_wb_data_i[27]
  PIN slave4_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 507.320 350.000 507.920 ;
    END
  END slave4_wb_data_i[28]
  PIN slave4_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 518.880 350.000 519.480 ;
    END
  END slave4_wb_data_i[29]
  PIN slave4_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 86.400 350.000 87.000 ;
    END
  END slave4_wb_data_i[2]
  PIN slave4_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 529.760 350.000 530.360 ;
    END
  END slave4_wb_data_i[30]
  PIN slave4_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 541.320 350.000 541.920 ;
    END
  END slave4_wb_data_i[31]
  PIN slave4_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 108.840 350.000 109.440 ;
    END
  END slave4_wb_data_i[3]
  PIN slave4_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 131.280 350.000 131.880 ;
    END
  END slave4_wb_data_i[4]
  PIN slave4_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 148.280 350.000 148.880 ;
    END
  END slave4_wb_data_i[5]
  PIN slave4_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 165.280 350.000 165.880 ;
    END
  END slave4_wb_data_i[6]
  PIN slave4_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 182.280 350.000 182.880 ;
    END
  END slave4_wb_data_i[7]
  PIN slave4_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 198.600 350.000 199.200 ;
    END
  END slave4_wb_data_i[8]
  PIN slave4_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 215.600 350.000 216.200 ;
    END
  END slave4_wb_data_i[9]
  PIN slave4_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 47.640 350.000 48.240 ;
    END
  END slave4_wb_data_o[0]
  PIN slave4_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 238.040 350.000 238.640 ;
    END
  END slave4_wb_data_o[10]
  PIN slave4_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 255.040 350.000 255.640 ;
    END
  END slave4_wb_data_o[11]
  PIN slave4_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 272.040 350.000 272.640 ;
    END
  END slave4_wb_data_o[12]
  PIN slave4_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 289.040 350.000 289.640 ;
    END
  END slave4_wb_data_o[13]
  PIN slave4_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 305.360 350.000 305.960 ;
    END
  END slave4_wb_data_o[14]
  PIN slave4_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 322.360 350.000 322.960 ;
    END
  END slave4_wb_data_o[15]
  PIN slave4_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 339.360 350.000 339.960 ;
    END
  END slave4_wb_data_o[16]
  PIN slave4_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 356.360 350.000 356.960 ;
    END
  END slave4_wb_data_o[17]
  PIN slave4_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 372.680 350.000 373.280 ;
    END
  END slave4_wb_data_o[18]
  PIN slave4_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 389.680 350.000 390.280 ;
    END
  END slave4_wb_data_o[19]
  PIN slave4_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 70.080 350.000 70.680 ;
    END
  END slave4_wb_data_o[1]
  PIN slave4_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 406.680 350.000 407.280 ;
    END
  END slave4_wb_data_o[20]
  PIN slave4_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 423.680 350.000 424.280 ;
    END
  END slave4_wb_data_o[21]
  PIN slave4_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 440.000 350.000 440.600 ;
    END
  END slave4_wb_data_o[22]
  PIN slave4_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 457.000 350.000 457.600 ;
    END
  END slave4_wb_data_o[23]
  PIN slave4_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 468.560 350.000 469.160 ;
    END
  END slave4_wb_data_o[24]
  PIN slave4_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 479.440 350.000 480.040 ;
    END
  END slave4_wb_data_o[25]
  PIN slave4_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 491.000 350.000 491.600 ;
    END
  END slave4_wb_data_o[26]
  PIN slave4_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 501.880 350.000 502.480 ;
    END
  END slave4_wb_data_o[27]
  PIN slave4_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 513.440 350.000 514.040 ;
    END
  END slave4_wb_data_o[28]
  PIN slave4_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 524.320 350.000 524.920 ;
    END
  END slave4_wb_data_o[29]
  PIN slave4_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 92.520 350.000 93.120 ;
    END
  END slave4_wb_data_o[2]
  PIN slave4_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 535.880 350.000 536.480 ;
    END
  END slave4_wb_data_o[30]
  PIN slave4_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 546.760 350.000 547.360 ;
    END
  END slave4_wb_data_o[31]
  PIN slave4_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 114.960 350.000 115.560 ;
    END
  END slave4_wb_data_o[3]
  PIN slave4_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 137.400 350.000 138.000 ;
    END
  END slave4_wb_data_o[4]
  PIN slave4_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 153.720 350.000 154.320 ;
    END
  END slave4_wb_data_o[5]
  PIN slave4_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 170.720 350.000 171.320 ;
    END
  END slave4_wb_data_o[6]
  PIN slave4_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 187.720 350.000 188.320 ;
    END
  END slave4_wb_data_o[7]
  PIN slave4_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 204.720 350.000 205.320 ;
    END
  END slave4_wb_data_o[8]
  PIN slave4_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 221.040 350.000 221.640 ;
    END
  END slave4_wb_data_o[9]
  PIN slave4_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 13.640 350.000 14.240 ;
    END
  END slave4_wb_error_o
  PIN slave4_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 53.080 350.000 53.680 ;
    END
  END slave4_wb_sel_i[0]
  PIN slave4_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 75.520 350.000 76.120 ;
    END
  END slave4_wb_sel_i[1]
  PIN slave4_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 97.960 350.000 98.560 ;
    END
  END slave4_wb_sel_i[2]
  PIN slave4_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 120.400 350.000 121.000 ;
    END
  END slave4_wb_sel_i[3]
  PIN slave4_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 19.080 350.000 19.680 ;
    END
  END slave4_wb_stall_o
  PIN slave4_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 25.200 350.000 25.800 ;
    END
  END slave4_wb_stb_i
  PIN slave4_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 30.640 350.000 31.240 ;
    END
  END slave4_wb_we_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1088.240 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 1088.085 ;
      LAYER met1 ;
        RECT 0.070 9.220 348.610 1088.980 ;
      LAYER met2 ;
        RECT 0.100 1095.720 1.190 1098.725 ;
        RECT 2.030 1095.720 4.410 1098.725 ;
        RECT 5.250 1095.720 8.090 1098.725 ;
        RECT 8.930 1095.720 11.770 1098.725 ;
        RECT 12.610 1095.720 15.450 1098.725 ;
        RECT 16.290 1095.720 18.670 1098.725 ;
        RECT 19.510 1095.720 22.350 1098.725 ;
        RECT 23.190 1095.720 26.030 1098.725 ;
        RECT 26.870 1095.720 29.710 1098.725 ;
        RECT 30.550 1095.720 32.930 1098.725 ;
        RECT 33.770 1095.720 36.610 1098.725 ;
        RECT 37.450 1095.720 40.290 1098.725 ;
        RECT 41.130 1095.720 43.970 1098.725 ;
        RECT 44.810 1095.720 47.190 1098.725 ;
        RECT 48.030 1095.720 50.870 1098.725 ;
        RECT 51.710 1095.720 54.550 1098.725 ;
        RECT 55.390 1095.720 58.230 1098.725 ;
        RECT 59.070 1095.720 61.910 1098.725 ;
        RECT 62.750 1095.720 65.130 1098.725 ;
        RECT 65.970 1095.720 68.810 1098.725 ;
        RECT 69.650 1095.720 72.490 1098.725 ;
        RECT 73.330 1095.720 76.170 1098.725 ;
        RECT 77.010 1095.720 79.390 1098.725 ;
        RECT 80.230 1095.720 83.070 1098.725 ;
        RECT 83.910 1095.720 86.750 1098.725 ;
        RECT 87.590 1095.720 90.430 1098.725 ;
        RECT 91.270 1095.720 93.650 1098.725 ;
        RECT 94.490 1095.720 97.330 1098.725 ;
        RECT 98.170 1095.720 101.010 1098.725 ;
        RECT 101.850 1095.720 104.690 1098.725 ;
        RECT 105.530 1095.720 107.910 1098.725 ;
        RECT 108.750 1095.720 111.590 1098.725 ;
        RECT 112.430 1095.720 115.270 1098.725 ;
        RECT 116.110 1095.720 118.950 1098.725 ;
        RECT 119.790 1095.720 122.630 1098.725 ;
        RECT 123.470 1095.720 125.850 1098.725 ;
        RECT 126.690 1095.720 129.530 1098.725 ;
        RECT 130.370 1095.720 133.210 1098.725 ;
        RECT 134.050 1095.720 136.890 1098.725 ;
        RECT 137.730 1095.720 140.110 1098.725 ;
        RECT 140.950 1095.720 143.790 1098.725 ;
        RECT 144.630 1095.720 147.470 1098.725 ;
        RECT 148.310 1095.720 151.150 1098.725 ;
        RECT 151.990 1095.720 154.370 1098.725 ;
        RECT 155.210 1095.720 158.050 1098.725 ;
        RECT 158.890 1095.720 161.730 1098.725 ;
        RECT 162.570 1095.720 165.410 1098.725 ;
        RECT 166.250 1095.720 168.630 1098.725 ;
        RECT 169.470 1095.720 172.310 1098.725 ;
        RECT 173.150 1095.720 175.990 1098.725 ;
        RECT 176.830 1095.720 179.670 1098.725 ;
        RECT 180.510 1095.720 183.350 1098.725 ;
        RECT 184.190 1095.720 186.570 1098.725 ;
        RECT 187.410 1095.720 190.250 1098.725 ;
        RECT 191.090 1095.720 193.930 1098.725 ;
        RECT 194.770 1095.720 197.610 1098.725 ;
        RECT 198.450 1095.720 200.830 1098.725 ;
        RECT 201.670 1095.720 204.510 1098.725 ;
        RECT 205.350 1095.720 208.190 1098.725 ;
        RECT 209.030 1095.720 211.870 1098.725 ;
        RECT 212.710 1095.720 215.090 1098.725 ;
        RECT 215.930 1095.720 218.770 1098.725 ;
        RECT 219.610 1095.720 222.450 1098.725 ;
        RECT 223.290 1095.720 226.130 1098.725 ;
        RECT 226.970 1095.720 229.350 1098.725 ;
        RECT 230.190 1095.720 233.030 1098.725 ;
        RECT 233.870 1095.720 236.710 1098.725 ;
        RECT 237.550 1095.720 240.390 1098.725 ;
        RECT 241.230 1095.720 244.070 1098.725 ;
        RECT 244.910 1095.720 247.290 1098.725 ;
        RECT 248.130 1095.720 250.970 1098.725 ;
        RECT 251.810 1095.720 254.650 1098.725 ;
        RECT 255.490 1095.720 258.330 1098.725 ;
        RECT 259.170 1095.720 261.550 1098.725 ;
        RECT 262.390 1095.720 265.230 1098.725 ;
        RECT 266.070 1095.720 268.910 1098.725 ;
        RECT 269.750 1095.720 272.590 1098.725 ;
        RECT 273.430 1095.720 275.810 1098.725 ;
        RECT 276.650 1095.720 279.490 1098.725 ;
        RECT 280.330 1095.720 283.170 1098.725 ;
        RECT 284.010 1095.720 286.850 1098.725 ;
        RECT 287.690 1095.720 290.070 1098.725 ;
        RECT 290.910 1095.720 293.750 1098.725 ;
        RECT 294.590 1095.720 297.430 1098.725 ;
        RECT 298.270 1095.720 301.110 1098.725 ;
        RECT 301.950 1095.720 304.790 1098.725 ;
        RECT 305.630 1095.720 308.010 1098.725 ;
        RECT 308.850 1095.720 311.690 1098.725 ;
        RECT 312.530 1095.720 315.370 1098.725 ;
        RECT 316.210 1095.720 319.050 1098.725 ;
        RECT 319.890 1095.720 322.270 1098.725 ;
        RECT 323.110 1095.720 325.950 1098.725 ;
        RECT 326.790 1095.720 329.630 1098.725 ;
        RECT 330.470 1095.720 333.310 1098.725 ;
        RECT 334.150 1095.720 336.530 1098.725 ;
        RECT 337.370 1095.720 340.210 1098.725 ;
        RECT 341.050 1095.720 343.890 1098.725 ;
        RECT 344.730 1095.720 347.570 1098.725 ;
        RECT 348.410 1095.720 348.580 1098.725 ;
        RECT 0.100 4.280 348.580 1095.720 ;
        RECT 0.100 1.515 1.190 4.280 ;
        RECT 2.030 1.515 3.950 4.280 ;
        RECT 4.790 1.515 6.710 4.280 ;
        RECT 7.550 1.515 9.930 4.280 ;
        RECT 10.770 1.515 12.690 4.280 ;
        RECT 13.530 1.515 15.450 4.280 ;
        RECT 16.290 1.515 18.670 4.280 ;
        RECT 19.510 1.515 21.430 4.280 ;
        RECT 22.270 1.515 24.190 4.280 ;
        RECT 25.030 1.515 27.410 4.280 ;
        RECT 28.250 1.515 30.170 4.280 ;
        RECT 31.010 1.515 32.930 4.280 ;
        RECT 33.770 1.515 36.150 4.280 ;
        RECT 36.990 1.515 38.910 4.280 ;
        RECT 39.750 1.515 41.670 4.280 ;
        RECT 42.510 1.515 44.890 4.280 ;
        RECT 45.730 1.515 47.650 4.280 ;
        RECT 48.490 1.515 50.410 4.280 ;
        RECT 51.250 1.515 53.630 4.280 ;
        RECT 54.470 1.515 56.390 4.280 ;
        RECT 57.230 1.515 59.150 4.280 ;
        RECT 59.990 1.515 62.370 4.280 ;
        RECT 63.210 1.515 65.130 4.280 ;
        RECT 65.970 1.515 67.890 4.280 ;
        RECT 68.730 1.515 71.110 4.280 ;
        RECT 71.950 1.515 73.870 4.280 ;
        RECT 74.710 1.515 76.630 4.280 ;
        RECT 77.470 1.515 79.850 4.280 ;
        RECT 80.690 1.515 82.610 4.280 ;
        RECT 83.450 1.515 85.370 4.280 ;
        RECT 86.210 1.515 88.590 4.280 ;
        RECT 89.430 1.515 91.350 4.280 ;
        RECT 92.190 1.515 94.110 4.280 ;
        RECT 94.950 1.515 97.330 4.280 ;
        RECT 98.170 1.515 100.090 4.280 ;
        RECT 100.930 1.515 102.850 4.280 ;
        RECT 103.690 1.515 106.070 4.280 ;
        RECT 106.910 1.515 108.830 4.280 ;
        RECT 109.670 1.515 111.590 4.280 ;
        RECT 112.430 1.515 114.810 4.280 ;
        RECT 115.650 1.515 117.570 4.280 ;
        RECT 118.410 1.515 120.790 4.280 ;
        RECT 121.630 1.515 123.550 4.280 ;
        RECT 124.390 1.515 126.310 4.280 ;
        RECT 127.150 1.515 129.530 4.280 ;
        RECT 130.370 1.515 132.290 4.280 ;
        RECT 133.130 1.515 135.050 4.280 ;
        RECT 135.890 1.515 138.270 4.280 ;
        RECT 139.110 1.515 141.030 4.280 ;
        RECT 141.870 1.515 143.790 4.280 ;
        RECT 144.630 1.515 147.010 4.280 ;
        RECT 147.850 1.515 149.770 4.280 ;
        RECT 150.610 1.515 152.530 4.280 ;
        RECT 153.370 1.515 155.750 4.280 ;
        RECT 156.590 1.515 158.510 4.280 ;
        RECT 159.350 1.515 161.270 4.280 ;
        RECT 162.110 1.515 164.490 4.280 ;
        RECT 165.330 1.515 167.250 4.280 ;
        RECT 168.090 1.515 170.010 4.280 ;
        RECT 170.850 1.515 173.230 4.280 ;
        RECT 174.070 1.515 175.990 4.280 ;
        RECT 176.830 1.515 178.750 4.280 ;
        RECT 179.590 1.515 181.970 4.280 ;
        RECT 182.810 1.515 184.730 4.280 ;
        RECT 185.570 1.515 187.490 4.280 ;
        RECT 188.330 1.515 190.710 4.280 ;
        RECT 191.550 1.515 193.470 4.280 ;
        RECT 194.310 1.515 196.230 4.280 ;
        RECT 197.070 1.515 199.450 4.280 ;
        RECT 200.290 1.515 202.210 4.280 ;
        RECT 203.050 1.515 204.970 4.280 ;
        RECT 205.810 1.515 208.190 4.280 ;
        RECT 209.030 1.515 210.950 4.280 ;
        RECT 211.790 1.515 213.710 4.280 ;
        RECT 214.550 1.515 216.930 4.280 ;
        RECT 217.770 1.515 219.690 4.280 ;
        RECT 220.530 1.515 222.450 4.280 ;
        RECT 223.290 1.515 225.670 4.280 ;
        RECT 226.510 1.515 228.430 4.280 ;
        RECT 229.270 1.515 231.190 4.280 ;
        RECT 232.030 1.515 234.410 4.280 ;
        RECT 235.250 1.515 237.170 4.280 ;
        RECT 238.010 1.515 240.390 4.280 ;
        RECT 241.230 1.515 243.150 4.280 ;
        RECT 243.990 1.515 245.910 4.280 ;
        RECT 246.750 1.515 249.130 4.280 ;
        RECT 249.970 1.515 251.890 4.280 ;
        RECT 252.730 1.515 254.650 4.280 ;
        RECT 255.490 1.515 257.870 4.280 ;
        RECT 258.710 1.515 260.630 4.280 ;
        RECT 261.470 1.515 263.390 4.280 ;
        RECT 264.230 1.515 266.610 4.280 ;
        RECT 267.450 1.515 269.370 4.280 ;
        RECT 270.210 1.515 272.130 4.280 ;
        RECT 272.970 1.515 275.350 4.280 ;
        RECT 276.190 1.515 278.110 4.280 ;
        RECT 278.950 1.515 280.870 4.280 ;
        RECT 281.710 1.515 284.090 4.280 ;
        RECT 284.930 1.515 286.850 4.280 ;
        RECT 287.690 1.515 289.610 4.280 ;
        RECT 290.450 1.515 292.830 4.280 ;
        RECT 293.670 1.515 295.590 4.280 ;
        RECT 296.430 1.515 298.350 4.280 ;
        RECT 299.190 1.515 301.570 4.280 ;
        RECT 302.410 1.515 304.330 4.280 ;
        RECT 305.170 1.515 307.090 4.280 ;
        RECT 307.930 1.515 310.310 4.280 ;
        RECT 311.150 1.515 313.070 4.280 ;
        RECT 313.910 1.515 315.830 4.280 ;
        RECT 316.670 1.515 319.050 4.280 ;
        RECT 319.890 1.515 321.810 4.280 ;
        RECT 322.650 1.515 324.570 4.280 ;
        RECT 325.410 1.515 327.790 4.280 ;
        RECT 328.630 1.515 330.550 4.280 ;
        RECT 331.390 1.515 333.310 4.280 ;
        RECT 334.150 1.515 336.530 4.280 ;
        RECT 337.370 1.515 339.290 4.280 ;
        RECT 340.130 1.515 342.050 4.280 ;
        RECT 342.890 1.515 345.270 4.280 ;
        RECT 346.110 1.515 348.030 4.280 ;
      LAYER met3 ;
        RECT 4.400 1097.880 346.000 1098.705 ;
        RECT 4.400 1097.840 345.600 1097.880 ;
        RECT 4.000 1096.520 345.600 1097.840 ;
        RECT 4.400 1096.480 345.600 1096.520 ;
        RECT 4.400 1095.120 346.000 1096.480 ;
        RECT 4.000 1093.800 346.000 1095.120 ;
        RECT 4.400 1092.440 346.000 1093.800 ;
        RECT 4.400 1092.400 345.600 1092.440 ;
        RECT 4.000 1091.080 345.600 1092.400 ;
        RECT 4.400 1091.040 345.600 1091.080 ;
        RECT 4.400 1089.680 346.000 1091.040 ;
        RECT 4.000 1088.360 346.000 1089.680 ;
        RECT 4.400 1087.000 346.000 1088.360 ;
        RECT 4.400 1086.960 345.600 1087.000 ;
        RECT 4.000 1085.640 345.600 1086.960 ;
        RECT 4.400 1085.600 345.600 1085.640 ;
        RECT 4.400 1084.240 346.000 1085.600 ;
        RECT 4.000 1082.920 346.000 1084.240 ;
        RECT 4.400 1081.520 346.000 1082.920 ;
        RECT 4.000 1080.880 346.000 1081.520 ;
        RECT 4.000 1080.200 345.600 1080.880 ;
        RECT 4.400 1079.480 345.600 1080.200 ;
        RECT 4.400 1078.800 346.000 1079.480 ;
        RECT 4.000 1077.480 346.000 1078.800 ;
        RECT 4.400 1076.080 346.000 1077.480 ;
        RECT 4.000 1075.440 346.000 1076.080 ;
        RECT 4.000 1074.760 345.600 1075.440 ;
        RECT 4.400 1074.040 345.600 1074.760 ;
        RECT 4.400 1073.360 346.000 1074.040 ;
        RECT 4.000 1072.040 346.000 1073.360 ;
        RECT 4.400 1070.640 346.000 1072.040 ;
        RECT 4.000 1070.000 346.000 1070.640 ;
        RECT 4.000 1069.320 345.600 1070.000 ;
        RECT 4.400 1068.600 345.600 1069.320 ;
        RECT 4.400 1067.920 346.000 1068.600 ;
        RECT 4.000 1066.600 346.000 1067.920 ;
        RECT 4.400 1065.200 346.000 1066.600 ;
        RECT 4.000 1064.560 346.000 1065.200 ;
        RECT 4.000 1063.880 345.600 1064.560 ;
        RECT 4.400 1063.160 345.600 1063.880 ;
        RECT 4.400 1062.480 346.000 1063.160 ;
        RECT 4.000 1061.160 346.000 1062.480 ;
        RECT 4.400 1059.760 346.000 1061.160 ;
        RECT 4.000 1058.440 346.000 1059.760 ;
        RECT 4.400 1057.040 345.600 1058.440 ;
        RECT 4.000 1055.720 346.000 1057.040 ;
        RECT 4.400 1054.320 346.000 1055.720 ;
        RECT 4.000 1053.000 346.000 1054.320 ;
        RECT 4.400 1051.600 345.600 1053.000 ;
        RECT 4.000 1050.280 346.000 1051.600 ;
        RECT 4.400 1048.880 346.000 1050.280 ;
        RECT 4.000 1047.560 346.000 1048.880 ;
        RECT 4.400 1046.160 345.600 1047.560 ;
        RECT 4.000 1044.840 346.000 1046.160 ;
        RECT 4.400 1043.440 346.000 1044.840 ;
        RECT 4.000 1042.120 346.000 1043.440 ;
        RECT 4.400 1040.720 345.600 1042.120 ;
        RECT 4.000 1038.720 346.000 1040.720 ;
        RECT 4.400 1037.320 346.000 1038.720 ;
        RECT 4.000 1036.000 346.000 1037.320 ;
        RECT 4.400 1034.600 345.600 1036.000 ;
        RECT 4.000 1033.280 346.000 1034.600 ;
        RECT 4.400 1031.880 346.000 1033.280 ;
        RECT 4.000 1030.560 346.000 1031.880 ;
        RECT 4.400 1029.160 345.600 1030.560 ;
        RECT 4.000 1027.840 346.000 1029.160 ;
        RECT 4.400 1026.440 346.000 1027.840 ;
        RECT 4.000 1025.120 346.000 1026.440 ;
        RECT 4.400 1023.720 345.600 1025.120 ;
        RECT 4.000 1022.400 346.000 1023.720 ;
        RECT 4.400 1021.000 346.000 1022.400 ;
        RECT 4.000 1019.680 346.000 1021.000 ;
        RECT 4.400 1018.280 345.600 1019.680 ;
        RECT 4.000 1016.960 346.000 1018.280 ;
        RECT 4.400 1015.560 346.000 1016.960 ;
        RECT 4.000 1014.240 346.000 1015.560 ;
        RECT 4.400 1013.560 346.000 1014.240 ;
        RECT 4.400 1012.840 345.600 1013.560 ;
        RECT 4.000 1012.160 345.600 1012.840 ;
        RECT 4.000 1011.520 346.000 1012.160 ;
        RECT 4.400 1010.120 346.000 1011.520 ;
        RECT 4.000 1008.800 346.000 1010.120 ;
        RECT 4.400 1008.120 346.000 1008.800 ;
        RECT 4.400 1007.400 345.600 1008.120 ;
        RECT 4.000 1006.720 345.600 1007.400 ;
        RECT 4.000 1006.080 346.000 1006.720 ;
        RECT 4.400 1004.680 346.000 1006.080 ;
        RECT 4.000 1003.360 346.000 1004.680 ;
        RECT 4.400 1002.680 346.000 1003.360 ;
        RECT 4.400 1001.960 345.600 1002.680 ;
        RECT 4.000 1001.280 345.600 1001.960 ;
        RECT 4.000 1000.640 346.000 1001.280 ;
        RECT 4.400 999.240 346.000 1000.640 ;
        RECT 4.000 997.920 346.000 999.240 ;
        RECT 4.400 997.240 346.000 997.920 ;
        RECT 4.400 996.520 345.600 997.240 ;
        RECT 4.000 995.840 345.600 996.520 ;
        RECT 4.000 995.200 346.000 995.840 ;
        RECT 4.400 993.800 346.000 995.200 ;
        RECT 4.000 992.480 346.000 993.800 ;
        RECT 4.400 991.120 346.000 992.480 ;
        RECT 4.400 991.080 345.600 991.120 ;
        RECT 4.000 989.760 345.600 991.080 ;
        RECT 4.400 989.720 345.600 989.760 ;
        RECT 4.400 988.360 346.000 989.720 ;
        RECT 4.000 987.040 346.000 988.360 ;
        RECT 4.400 985.680 346.000 987.040 ;
        RECT 4.400 985.640 345.600 985.680 ;
        RECT 4.000 984.320 345.600 985.640 ;
        RECT 4.400 984.280 345.600 984.320 ;
        RECT 4.400 982.920 346.000 984.280 ;
        RECT 4.000 981.600 346.000 982.920 ;
        RECT 4.400 980.240 346.000 981.600 ;
        RECT 4.400 980.200 345.600 980.240 ;
        RECT 4.000 978.840 345.600 980.200 ;
        RECT 4.000 978.200 346.000 978.840 ;
        RECT 4.400 976.800 346.000 978.200 ;
        RECT 4.000 975.480 346.000 976.800 ;
        RECT 4.400 974.800 346.000 975.480 ;
        RECT 4.400 974.080 345.600 974.800 ;
        RECT 4.000 973.400 345.600 974.080 ;
        RECT 4.000 972.760 346.000 973.400 ;
        RECT 4.400 971.360 346.000 972.760 ;
        RECT 4.000 970.040 346.000 971.360 ;
        RECT 4.400 968.680 346.000 970.040 ;
        RECT 4.400 968.640 345.600 968.680 ;
        RECT 4.000 967.320 345.600 968.640 ;
        RECT 4.400 967.280 345.600 967.320 ;
        RECT 4.400 965.920 346.000 967.280 ;
        RECT 4.000 964.600 346.000 965.920 ;
        RECT 4.400 963.240 346.000 964.600 ;
        RECT 4.400 963.200 345.600 963.240 ;
        RECT 4.000 961.880 345.600 963.200 ;
        RECT 4.400 961.840 345.600 961.880 ;
        RECT 4.400 960.480 346.000 961.840 ;
        RECT 4.000 959.160 346.000 960.480 ;
        RECT 4.400 957.800 346.000 959.160 ;
        RECT 4.400 957.760 345.600 957.800 ;
        RECT 4.000 956.440 345.600 957.760 ;
        RECT 4.400 956.400 345.600 956.440 ;
        RECT 4.400 955.040 346.000 956.400 ;
        RECT 4.000 953.720 346.000 955.040 ;
        RECT 4.400 952.360 346.000 953.720 ;
        RECT 4.400 952.320 345.600 952.360 ;
        RECT 4.000 951.000 345.600 952.320 ;
        RECT 4.400 950.960 345.600 951.000 ;
        RECT 4.400 949.600 346.000 950.960 ;
        RECT 4.000 948.280 346.000 949.600 ;
        RECT 4.400 946.880 346.000 948.280 ;
        RECT 4.000 946.240 346.000 946.880 ;
        RECT 4.000 945.560 345.600 946.240 ;
        RECT 4.400 944.840 345.600 945.560 ;
        RECT 4.400 944.160 346.000 944.840 ;
        RECT 4.000 942.840 346.000 944.160 ;
        RECT 4.400 941.440 346.000 942.840 ;
        RECT 4.000 940.800 346.000 941.440 ;
        RECT 4.000 940.120 345.600 940.800 ;
        RECT 4.400 939.400 345.600 940.120 ;
        RECT 4.400 938.720 346.000 939.400 ;
        RECT 4.000 937.400 346.000 938.720 ;
        RECT 4.400 936.000 346.000 937.400 ;
        RECT 4.000 935.360 346.000 936.000 ;
        RECT 4.000 934.680 345.600 935.360 ;
        RECT 4.400 933.960 345.600 934.680 ;
        RECT 4.400 933.280 346.000 933.960 ;
        RECT 4.000 931.960 346.000 933.280 ;
        RECT 4.400 930.560 346.000 931.960 ;
        RECT 4.000 929.920 346.000 930.560 ;
        RECT 4.000 929.240 345.600 929.920 ;
        RECT 4.400 928.520 345.600 929.240 ;
        RECT 4.400 927.840 346.000 928.520 ;
        RECT 4.000 926.520 346.000 927.840 ;
        RECT 4.400 925.120 346.000 926.520 ;
        RECT 4.000 923.800 346.000 925.120 ;
        RECT 4.400 922.400 345.600 923.800 ;
        RECT 4.000 921.080 346.000 922.400 ;
        RECT 4.400 919.680 346.000 921.080 ;
        RECT 4.000 918.360 346.000 919.680 ;
        RECT 4.000 917.680 345.600 918.360 ;
        RECT 4.400 916.960 345.600 917.680 ;
        RECT 4.400 916.280 346.000 916.960 ;
        RECT 4.000 914.960 346.000 916.280 ;
        RECT 4.400 913.560 346.000 914.960 ;
        RECT 4.000 912.920 346.000 913.560 ;
        RECT 4.000 912.240 345.600 912.920 ;
        RECT 4.400 911.520 345.600 912.240 ;
        RECT 4.400 910.840 346.000 911.520 ;
        RECT 4.000 909.520 346.000 910.840 ;
        RECT 4.400 908.120 346.000 909.520 ;
        RECT 4.000 907.480 346.000 908.120 ;
        RECT 4.000 906.800 345.600 907.480 ;
        RECT 4.400 906.080 345.600 906.800 ;
        RECT 4.400 905.400 346.000 906.080 ;
        RECT 4.000 904.080 346.000 905.400 ;
        RECT 4.400 902.680 346.000 904.080 ;
        RECT 4.000 901.360 346.000 902.680 ;
        RECT 4.400 899.960 345.600 901.360 ;
        RECT 4.000 898.640 346.000 899.960 ;
        RECT 4.400 897.240 346.000 898.640 ;
        RECT 4.000 895.920 346.000 897.240 ;
        RECT 4.400 894.520 345.600 895.920 ;
        RECT 4.000 893.200 346.000 894.520 ;
        RECT 4.400 891.800 346.000 893.200 ;
        RECT 4.000 890.480 346.000 891.800 ;
        RECT 4.400 889.080 345.600 890.480 ;
        RECT 4.000 887.760 346.000 889.080 ;
        RECT 4.400 886.360 346.000 887.760 ;
        RECT 4.000 885.040 346.000 886.360 ;
        RECT 4.400 883.640 345.600 885.040 ;
        RECT 4.000 882.320 346.000 883.640 ;
        RECT 4.400 880.920 346.000 882.320 ;
        RECT 4.000 879.600 346.000 880.920 ;
        RECT 4.400 878.920 346.000 879.600 ;
        RECT 4.400 878.200 345.600 878.920 ;
        RECT 4.000 877.520 345.600 878.200 ;
        RECT 4.000 876.880 346.000 877.520 ;
        RECT 4.400 875.480 346.000 876.880 ;
        RECT 4.000 874.160 346.000 875.480 ;
        RECT 4.400 873.480 346.000 874.160 ;
        RECT 4.400 872.760 345.600 873.480 ;
        RECT 4.000 872.080 345.600 872.760 ;
        RECT 4.000 871.440 346.000 872.080 ;
        RECT 4.400 870.040 346.000 871.440 ;
        RECT 4.000 868.720 346.000 870.040 ;
        RECT 4.400 868.040 346.000 868.720 ;
        RECT 4.400 867.320 345.600 868.040 ;
        RECT 4.000 866.640 345.600 867.320 ;
        RECT 4.000 866.000 346.000 866.640 ;
        RECT 4.400 864.600 346.000 866.000 ;
        RECT 4.000 863.280 346.000 864.600 ;
        RECT 4.400 862.600 346.000 863.280 ;
        RECT 4.400 861.880 345.600 862.600 ;
        RECT 4.000 861.200 345.600 861.880 ;
        RECT 4.000 860.560 346.000 861.200 ;
        RECT 4.400 859.160 346.000 860.560 ;
        RECT 4.000 857.160 346.000 859.160 ;
        RECT 4.400 856.480 346.000 857.160 ;
        RECT 4.400 855.760 345.600 856.480 ;
        RECT 4.000 855.080 345.600 855.760 ;
        RECT 4.000 854.440 346.000 855.080 ;
        RECT 4.400 853.040 346.000 854.440 ;
        RECT 4.000 851.720 346.000 853.040 ;
        RECT 4.400 851.040 346.000 851.720 ;
        RECT 4.400 850.320 345.600 851.040 ;
        RECT 4.000 849.640 345.600 850.320 ;
        RECT 4.000 849.000 346.000 849.640 ;
        RECT 4.400 847.600 346.000 849.000 ;
        RECT 4.000 846.280 346.000 847.600 ;
        RECT 4.400 845.600 346.000 846.280 ;
        RECT 4.400 844.880 345.600 845.600 ;
        RECT 4.000 844.200 345.600 844.880 ;
        RECT 4.000 843.560 346.000 844.200 ;
        RECT 4.400 842.160 346.000 843.560 ;
        RECT 4.000 840.840 346.000 842.160 ;
        RECT 4.400 840.160 346.000 840.840 ;
        RECT 4.400 839.440 345.600 840.160 ;
        RECT 4.000 838.760 345.600 839.440 ;
        RECT 4.000 838.120 346.000 838.760 ;
        RECT 4.400 836.720 346.000 838.120 ;
        RECT 4.000 835.400 346.000 836.720 ;
        RECT 4.400 834.040 346.000 835.400 ;
        RECT 4.400 834.000 345.600 834.040 ;
        RECT 4.000 832.680 345.600 834.000 ;
        RECT 4.400 832.640 345.600 832.680 ;
        RECT 4.400 831.280 346.000 832.640 ;
        RECT 4.000 829.960 346.000 831.280 ;
        RECT 4.400 828.600 346.000 829.960 ;
        RECT 4.400 828.560 345.600 828.600 ;
        RECT 4.000 827.240 345.600 828.560 ;
        RECT 4.400 827.200 345.600 827.240 ;
        RECT 4.400 825.840 346.000 827.200 ;
        RECT 4.000 824.520 346.000 825.840 ;
        RECT 4.400 823.160 346.000 824.520 ;
        RECT 4.400 823.120 345.600 823.160 ;
        RECT 4.000 821.800 345.600 823.120 ;
        RECT 4.400 821.760 345.600 821.800 ;
        RECT 4.400 820.400 346.000 821.760 ;
        RECT 4.000 819.080 346.000 820.400 ;
        RECT 4.400 817.680 346.000 819.080 ;
        RECT 4.000 817.040 346.000 817.680 ;
        RECT 4.000 816.360 345.600 817.040 ;
        RECT 4.400 815.640 345.600 816.360 ;
        RECT 4.400 814.960 346.000 815.640 ;
        RECT 4.000 813.640 346.000 814.960 ;
        RECT 4.400 812.240 346.000 813.640 ;
        RECT 4.000 811.600 346.000 812.240 ;
        RECT 4.000 810.920 345.600 811.600 ;
        RECT 4.400 810.200 345.600 810.920 ;
        RECT 4.400 809.520 346.000 810.200 ;
        RECT 4.000 808.200 346.000 809.520 ;
        RECT 4.400 806.800 346.000 808.200 ;
        RECT 4.000 806.160 346.000 806.800 ;
        RECT 4.000 805.480 345.600 806.160 ;
        RECT 4.400 804.760 345.600 805.480 ;
        RECT 4.400 804.080 346.000 804.760 ;
        RECT 4.000 802.760 346.000 804.080 ;
        RECT 4.400 801.360 346.000 802.760 ;
        RECT 4.000 800.720 346.000 801.360 ;
        RECT 4.000 800.040 345.600 800.720 ;
        RECT 4.400 799.320 345.600 800.040 ;
        RECT 4.400 798.640 346.000 799.320 ;
        RECT 4.000 797.320 346.000 798.640 ;
        RECT 4.400 795.920 346.000 797.320 ;
        RECT 4.000 794.600 346.000 795.920 ;
        RECT 4.000 793.920 345.600 794.600 ;
        RECT 4.400 793.200 345.600 793.920 ;
        RECT 4.400 792.520 346.000 793.200 ;
        RECT 4.000 791.200 346.000 792.520 ;
        RECT 4.400 789.800 346.000 791.200 ;
        RECT 4.000 789.160 346.000 789.800 ;
        RECT 4.000 788.480 345.600 789.160 ;
        RECT 4.400 787.760 345.600 788.480 ;
        RECT 4.400 787.080 346.000 787.760 ;
        RECT 4.000 785.760 346.000 787.080 ;
        RECT 4.400 784.360 346.000 785.760 ;
        RECT 4.000 783.720 346.000 784.360 ;
        RECT 4.000 783.040 345.600 783.720 ;
        RECT 4.400 782.320 345.600 783.040 ;
        RECT 4.400 781.640 346.000 782.320 ;
        RECT 4.000 780.320 346.000 781.640 ;
        RECT 4.400 778.920 346.000 780.320 ;
        RECT 4.000 778.280 346.000 778.920 ;
        RECT 4.000 777.600 345.600 778.280 ;
        RECT 4.400 776.880 345.600 777.600 ;
        RECT 4.400 776.200 346.000 776.880 ;
        RECT 4.000 774.880 346.000 776.200 ;
        RECT 4.400 773.480 346.000 774.880 ;
        RECT 4.000 772.160 346.000 773.480 ;
        RECT 4.400 770.760 345.600 772.160 ;
        RECT 4.000 769.440 346.000 770.760 ;
        RECT 4.400 768.040 346.000 769.440 ;
        RECT 4.000 766.720 346.000 768.040 ;
        RECT 4.400 765.320 345.600 766.720 ;
        RECT 4.000 764.000 346.000 765.320 ;
        RECT 4.400 762.600 346.000 764.000 ;
        RECT 4.000 761.280 346.000 762.600 ;
        RECT 4.400 759.880 345.600 761.280 ;
        RECT 4.000 758.560 346.000 759.880 ;
        RECT 4.400 757.160 346.000 758.560 ;
        RECT 4.000 755.840 346.000 757.160 ;
        RECT 4.400 754.440 345.600 755.840 ;
        RECT 4.000 753.120 346.000 754.440 ;
        RECT 4.400 751.720 346.000 753.120 ;
        RECT 4.000 750.400 346.000 751.720 ;
        RECT 4.400 749.720 346.000 750.400 ;
        RECT 4.400 749.000 345.600 749.720 ;
        RECT 4.000 748.320 345.600 749.000 ;
        RECT 4.000 747.680 346.000 748.320 ;
        RECT 4.400 746.280 346.000 747.680 ;
        RECT 4.000 744.960 346.000 746.280 ;
        RECT 4.400 744.280 346.000 744.960 ;
        RECT 4.400 743.560 345.600 744.280 ;
        RECT 4.000 742.880 345.600 743.560 ;
        RECT 4.000 742.240 346.000 742.880 ;
        RECT 4.400 740.840 346.000 742.240 ;
        RECT 4.000 739.520 346.000 740.840 ;
        RECT 4.400 738.840 346.000 739.520 ;
        RECT 4.400 738.120 345.600 738.840 ;
        RECT 4.000 737.440 345.600 738.120 ;
        RECT 4.000 736.800 346.000 737.440 ;
        RECT 4.400 735.400 346.000 736.800 ;
        RECT 4.000 733.400 346.000 735.400 ;
        RECT 4.400 732.000 345.600 733.400 ;
        RECT 4.000 730.680 346.000 732.000 ;
        RECT 4.400 729.280 346.000 730.680 ;
        RECT 4.000 727.960 346.000 729.280 ;
        RECT 4.400 727.280 346.000 727.960 ;
        RECT 4.400 726.560 345.600 727.280 ;
        RECT 4.000 725.880 345.600 726.560 ;
        RECT 4.000 725.240 346.000 725.880 ;
        RECT 4.400 723.840 346.000 725.240 ;
        RECT 4.000 722.520 346.000 723.840 ;
        RECT 4.400 721.840 346.000 722.520 ;
        RECT 4.400 721.120 345.600 721.840 ;
        RECT 4.000 720.440 345.600 721.120 ;
        RECT 4.000 719.800 346.000 720.440 ;
        RECT 4.400 718.400 346.000 719.800 ;
        RECT 4.000 717.080 346.000 718.400 ;
        RECT 4.400 716.400 346.000 717.080 ;
        RECT 4.400 715.680 345.600 716.400 ;
        RECT 4.000 715.000 345.600 715.680 ;
        RECT 4.000 714.360 346.000 715.000 ;
        RECT 4.400 712.960 346.000 714.360 ;
        RECT 4.000 711.640 346.000 712.960 ;
        RECT 4.400 710.960 346.000 711.640 ;
        RECT 4.400 710.240 345.600 710.960 ;
        RECT 4.000 709.560 345.600 710.240 ;
        RECT 4.000 708.920 346.000 709.560 ;
        RECT 4.400 707.520 346.000 708.920 ;
        RECT 4.000 706.200 346.000 707.520 ;
        RECT 4.400 704.840 346.000 706.200 ;
        RECT 4.400 704.800 345.600 704.840 ;
        RECT 4.000 703.480 345.600 704.800 ;
        RECT 4.400 703.440 345.600 703.480 ;
        RECT 4.400 702.080 346.000 703.440 ;
        RECT 4.000 700.760 346.000 702.080 ;
        RECT 4.400 699.400 346.000 700.760 ;
        RECT 4.400 699.360 345.600 699.400 ;
        RECT 4.000 698.040 345.600 699.360 ;
        RECT 4.400 698.000 345.600 698.040 ;
        RECT 4.400 696.640 346.000 698.000 ;
        RECT 4.000 695.320 346.000 696.640 ;
        RECT 4.400 693.960 346.000 695.320 ;
        RECT 4.400 693.920 345.600 693.960 ;
        RECT 4.000 692.600 345.600 693.920 ;
        RECT 4.400 692.560 345.600 692.600 ;
        RECT 4.400 691.200 346.000 692.560 ;
        RECT 4.000 689.880 346.000 691.200 ;
        RECT 4.400 688.520 346.000 689.880 ;
        RECT 4.400 688.480 345.600 688.520 ;
        RECT 4.000 687.160 345.600 688.480 ;
        RECT 4.400 687.120 345.600 687.160 ;
        RECT 4.400 685.760 346.000 687.120 ;
        RECT 4.000 684.440 346.000 685.760 ;
        RECT 4.400 683.040 346.000 684.440 ;
        RECT 4.000 682.400 346.000 683.040 ;
        RECT 4.000 681.720 345.600 682.400 ;
        RECT 4.400 681.000 345.600 681.720 ;
        RECT 4.400 680.320 346.000 681.000 ;
        RECT 4.000 679.000 346.000 680.320 ;
        RECT 4.400 677.600 346.000 679.000 ;
        RECT 4.000 676.960 346.000 677.600 ;
        RECT 4.000 676.280 345.600 676.960 ;
        RECT 4.400 675.560 345.600 676.280 ;
        RECT 4.400 674.880 346.000 675.560 ;
        RECT 4.000 672.880 346.000 674.880 ;
        RECT 4.400 671.520 346.000 672.880 ;
        RECT 4.400 671.480 345.600 671.520 ;
        RECT 4.000 670.160 345.600 671.480 ;
        RECT 4.400 670.120 345.600 670.160 ;
        RECT 4.400 668.760 346.000 670.120 ;
        RECT 4.000 667.440 346.000 668.760 ;
        RECT 4.400 666.080 346.000 667.440 ;
        RECT 4.400 666.040 345.600 666.080 ;
        RECT 4.000 664.720 345.600 666.040 ;
        RECT 4.400 664.680 345.600 664.720 ;
        RECT 4.400 663.320 346.000 664.680 ;
        RECT 4.000 662.000 346.000 663.320 ;
        RECT 4.400 660.600 346.000 662.000 ;
        RECT 4.000 659.960 346.000 660.600 ;
        RECT 4.000 659.280 345.600 659.960 ;
        RECT 4.400 658.560 345.600 659.280 ;
        RECT 4.400 657.880 346.000 658.560 ;
        RECT 4.000 656.560 346.000 657.880 ;
        RECT 4.400 655.160 346.000 656.560 ;
        RECT 4.000 654.520 346.000 655.160 ;
        RECT 4.000 653.840 345.600 654.520 ;
        RECT 4.400 653.120 345.600 653.840 ;
        RECT 4.400 652.440 346.000 653.120 ;
        RECT 4.000 651.120 346.000 652.440 ;
        RECT 4.400 649.720 346.000 651.120 ;
        RECT 4.000 649.080 346.000 649.720 ;
        RECT 4.000 648.400 345.600 649.080 ;
        RECT 4.400 647.680 345.600 648.400 ;
        RECT 4.400 647.000 346.000 647.680 ;
        RECT 4.000 645.680 346.000 647.000 ;
        RECT 4.400 644.280 346.000 645.680 ;
        RECT 4.000 643.640 346.000 644.280 ;
        RECT 4.000 642.960 345.600 643.640 ;
        RECT 4.400 642.240 345.600 642.960 ;
        RECT 4.400 641.560 346.000 642.240 ;
        RECT 4.000 640.240 346.000 641.560 ;
        RECT 4.400 638.840 346.000 640.240 ;
        RECT 4.000 637.520 346.000 638.840 ;
        RECT 4.400 636.120 345.600 637.520 ;
        RECT 4.000 634.800 346.000 636.120 ;
        RECT 4.400 633.400 346.000 634.800 ;
        RECT 4.000 632.080 346.000 633.400 ;
        RECT 4.400 630.680 345.600 632.080 ;
        RECT 4.000 629.360 346.000 630.680 ;
        RECT 4.400 627.960 346.000 629.360 ;
        RECT 4.000 626.640 346.000 627.960 ;
        RECT 4.400 625.240 345.600 626.640 ;
        RECT 4.000 623.920 346.000 625.240 ;
        RECT 4.400 622.520 346.000 623.920 ;
        RECT 4.000 621.200 346.000 622.520 ;
        RECT 4.400 619.800 345.600 621.200 ;
        RECT 4.000 618.480 346.000 619.800 ;
        RECT 4.400 617.080 346.000 618.480 ;
        RECT 4.000 615.760 346.000 617.080 ;
        RECT 4.400 615.080 346.000 615.760 ;
        RECT 4.400 614.360 345.600 615.080 ;
        RECT 4.000 613.680 345.600 614.360 ;
        RECT 4.000 612.360 346.000 613.680 ;
        RECT 4.400 610.960 346.000 612.360 ;
        RECT 4.000 609.640 346.000 610.960 ;
        RECT 4.400 608.240 345.600 609.640 ;
        RECT 4.000 606.920 346.000 608.240 ;
        RECT 4.400 605.520 346.000 606.920 ;
        RECT 4.000 604.200 346.000 605.520 ;
        RECT 4.400 602.800 345.600 604.200 ;
        RECT 4.000 601.480 346.000 602.800 ;
        RECT 4.400 600.080 346.000 601.480 ;
        RECT 4.000 598.760 346.000 600.080 ;
        RECT 4.400 597.360 345.600 598.760 ;
        RECT 4.000 596.040 346.000 597.360 ;
        RECT 4.400 594.640 346.000 596.040 ;
        RECT 4.000 593.320 346.000 594.640 ;
        RECT 4.400 592.640 346.000 593.320 ;
        RECT 4.400 591.920 345.600 592.640 ;
        RECT 4.000 591.240 345.600 591.920 ;
        RECT 4.000 590.600 346.000 591.240 ;
        RECT 4.400 589.200 346.000 590.600 ;
        RECT 4.000 587.880 346.000 589.200 ;
        RECT 4.400 587.200 346.000 587.880 ;
        RECT 4.400 586.480 345.600 587.200 ;
        RECT 4.000 585.800 345.600 586.480 ;
        RECT 4.000 585.160 346.000 585.800 ;
        RECT 4.400 583.760 346.000 585.160 ;
        RECT 4.000 582.440 346.000 583.760 ;
        RECT 4.400 581.760 346.000 582.440 ;
        RECT 4.400 581.040 345.600 581.760 ;
        RECT 4.000 580.360 345.600 581.040 ;
        RECT 4.000 579.720 346.000 580.360 ;
        RECT 4.400 578.320 346.000 579.720 ;
        RECT 4.000 577.000 346.000 578.320 ;
        RECT 4.400 576.320 346.000 577.000 ;
        RECT 4.400 575.600 345.600 576.320 ;
        RECT 4.000 574.920 345.600 575.600 ;
        RECT 4.000 574.280 346.000 574.920 ;
        RECT 4.400 572.880 346.000 574.280 ;
        RECT 4.000 571.560 346.000 572.880 ;
        RECT 4.400 570.200 346.000 571.560 ;
        RECT 4.400 570.160 345.600 570.200 ;
        RECT 4.000 568.840 345.600 570.160 ;
        RECT 4.400 568.800 345.600 568.840 ;
        RECT 4.400 567.440 346.000 568.800 ;
        RECT 4.000 566.120 346.000 567.440 ;
        RECT 4.400 564.760 346.000 566.120 ;
        RECT 4.400 564.720 345.600 564.760 ;
        RECT 4.000 563.400 345.600 564.720 ;
        RECT 4.400 563.360 345.600 563.400 ;
        RECT 4.400 562.000 346.000 563.360 ;
        RECT 4.000 560.680 346.000 562.000 ;
        RECT 4.400 559.320 346.000 560.680 ;
        RECT 4.400 559.280 345.600 559.320 ;
        RECT 4.000 557.960 345.600 559.280 ;
        RECT 4.400 557.920 345.600 557.960 ;
        RECT 4.400 556.560 346.000 557.920 ;
        RECT 4.000 555.240 346.000 556.560 ;
        RECT 4.400 553.880 346.000 555.240 ;
        RECT 4.400 553.840 345.600 553.880 ;
        RECT 4.000 552.520 345.600 553.840 ;
        RECT 4.400 552.480 345.600 552.520 ;
        RECT 4.400 551.120 346.000 552.480 ;
        RECT 4.000 549.120 346.000 551.120 ;
        RECT 4.400 547.760 346.000 549.120 ;
        RECT 4.400 547.720 345.600 547.760 ;
        RECT 4.000 546.400 345.600 547.720 ;
        RECT 4.400 546.360 345.600 546.400 ;
        RECT 4.400 545.000 346.000 546.360 ;
        RECT 4.000 543.680 346.000 545.000 ;
        RECT 4.400 542.320 346.000 543.680 ;
        RECT 4.400 542.280 345.600 542.320 ;
        RECT 4.000 540.960 345.600 542.280 ;
        RECT 4.400 540.920 345.600 540.960 ;
        RECT 4.400 539.560 346.000 540.920 ;
        RECT 4.000 538.240 346.000 539.560 ;
        RECT 4.400 536.880 346.000 538.240 ;
        RECT 4.400 536.840 345.600 536.880 ;
        RECT 4.000 535.520 345.600 536.840 ;
        RECT 4.400 535.480 345.600 535.520 ;
        RECT 4.400 534.120 346.000 535.480 ;
        RECT 4.000 532.800 346.000 534.120 ;
        RECT 4.400 531.400 346.000 532.800 ;
        RECT 4.000 530.760 346.000 531.400 ;
        RECT 4.000 530.080 345.600 530.760 ;
        RECT 4.400 529.360 345.600 530.080 ;
        RECT 4.400 528.680 346.000 529.360 ;
        RECT 4.000 527.360 346.000 528.680 ;
        RECT 4.400 525.960 346.000 527.360 ;
        RECT 4.000 525.320 346.000 525.960 ;
        RECT 4.000 524.640 345.600 525.320 ;
        RECT 4.400 523.920 345.600 524.640 ;
        RECT 4.400 523.240 346.000 523.920 ;
        RECT 4.000 521.920 346.000 523.240 ;
        RECT 4.400 520.520 346.000 521.920 ;
        RECT 4.000 519.880 346.000 520.520 ;
        RECT 4.000 519.200 345.600 519.880 ;
        RECT 4.400 518.480 345.600 519.200 ;
        RECT 4.400 517.800 346.000 518.480 ;
        RECT 4.000 516.480 346.000 517.800 ;
        RECT 4.400 515.080 346.000 516.480 ;
        RECT 4.000 514.440 346.000 515.080 ;
        RECT 4.000 513.760 345.600 514.440 ;
        RECT 4.400 513.040 345.600 513.760 ;
        RECT 4.400 512.360 346.000 513.040 ;
        RECT 4.000 511.040 346.000 512.360 ;
        RECT 4.400 509.640 346.000 511.040 ;
        RECT 4.000 508.320 346.000 509.640 ;
        RECT 4.400 506.920 345.600 508.320 ;
        RECT 4.000 505.600 346.000 506.920 ;
        RECT 4.400 504.200 346.000 505.600 ;
        RECT 4.000 502.880 346.000 504.200 ;
        RECT 4.400 501.480 345.600 502.880 ;
        RECT 4.000 500.160 346.000 501.480 ;
        RECT 4.400 498.760 346.000 500.160 ;
        RECT 4.000 497.440 346.000 498.760 ;
        RECT 4.400 496.040 345.600 497.440 ;
        RECT 4.000 494.720 346.000 496.040 ;
        RECT 4.400 493.320 346.000 494.720 ;
        RECT 4.000 492.000 346.000 493.320 ;
        RECT 4.400 490.600 345.600 492.000 ;
        RECT 4.000 488.600 346.000 490.600 ;
        RECT 4.400 487.200 346.000 488.600 ;
        RECT 4.000 485.880 346.000 487.200 ;
        RECT 4.400 484.480 345.600 485.880 ;
        RECT 4.000 483.160 346.000 484.480 ;
        RECT 4.400 481.760 346.000 483.160 ;
        RECT 4.000 480.440 346.000 481.760 ;
        RECT 4.400 479.040 345.600 480.440 ;
        RECT 4.000 477.720 346.000 479.040 ;
        RECT 4.400 476.320 346.000 477.720 ;
        RECT 4.000 475.000 346.000 476.320 ;
        RECT 4.400 473.600 345.600 475.000 ;
        RECT 4.000 472.280 346.000 473.600 ;
        RECT 4.400 470.880 346.000 472.280 ;
        RECT 4.000 469.560 346.000 470.880 ;
        RECT 4.400 468.160 345.600 469.560 ;
        RECT 4.000 466.840 346.000 468.160 ;
        RECT 4.400 465.440 346.000 466.840 ;
        RECT 4.000 464.120 346.000 465.440 ;
        RECT 4.400 463.440 346.000 464.120 ;
        RECT 4.400 462.720 345.600 463.440 ;
        RECT 4.000 462.040 345.600 462.720 ;
        RECT 4.000 461.400 346.000 462.040 ;
        RECT 4.400 460.000 346.000 461.400 ;
        RECT 4.000 458.680 346.000 460.000 ;
        RECT 4.400 458.000 346.000 458.680 ;
        RECT 4.400 457.280 345.600 458.000 ;
        RECT 4.000 456.600 345.600 457.280 ;
        RECT 4.000 455.960 346.000 456.600 ;
        RECT 4.400 454.560 346.000 455.960 ;
        RECT 4.000 453.240 346.000 454.560 ;
        RECT 4.400 452.560 346.000 453.240 ;
        RECT 4.400 451.840 345.600 452.560 ;
        RECT 4.000 451.160 345.600 451.840 ;
        RECT 4.000 450.520 346.000 451.160 ;
        RECT 4.400 449.120 346.000 450.520 ;
        RECT 4.000 447.800 346.000 449.120 ;
        RECT 4.400 447.120 346.000 447.800 ;
        RECT 4.400 446.400 345.600 447.120 ;
        RECT 4.000 445.720 345.600 446.400 ;
        RECT 4.000 445.080 346.000 445.720 ;
        RECT 4.400 443.680 346.000 445.080 ;
        RECT 4.000 442.360 346.000 443.680 ;
        RECT 4.400 441.000 346.000 442.360 ;
        RECT 4.400 440.960 345.600 441.000 ;
        RECT 4.000 439.640 345.600 440.960 ;
        RECT 4.400 439.600 345.600 439.640 ;
        RECT 4.400 438.240 346.000 439.600 ;
        RECT 4.000 436.920 346.000 438.240 ;
        RECT 4.400 435.560 346.000 436.920 ;
        RECT 4.400 435.520 345.600 435.560 ;
        RECT 4.000 434.200 345.600 435.520 ;
        RECT 4.400 434.160 345.600 434.200 ;
        RECT 4.400 432.800 346.000 434.160 ;
        RECT 4.000 431.480 346.000 432.800 ;
        RECT 4.400 430.120 346.000 431.480 ;
        RECT 4.400 430.080 345.600 430.120 ;
        RECT 4.000 428.720 345.600 430.080 ;
        RECT 4.000 428.080 346.000 428.720 ;
        RECT 4.400 426.680 346.000 428.080 ;
        RECT 4.000 425.360 346.000 426.680 ;
        RECT 4.400 424.680 346.000 425.360 ;
        RECT 4.400 423.960 345.600 424.680 ;
        RECT 4.000 423.280 345.600 423.960 ;
        RECT 4.000 422.640 346.000 423.280 ;
        RECT 4.400 421.240 346.000 422.640 ;
        RECT 4.000 419.920 346.000 421.240 ;
        RECT 4.400 418.560 346.000 419.920 ;
        RECT 4.400 418.520 345.600 418.560 ;
        RECT 4.000 417.200 345.600 418.520 ;
        RECT 4.400 417.160 345.600 417.200 ;
        RECT 4.400 415.800 346.000 417.160 ;
        RECT 4.000 414.480 346.000 415.800 ;
        RECT 4.400 413.120 346.000 414.480 ;
        RECT 4.400 413.080 345.600 413.120 ;
        RECT 4.000 411.760 345.600 413.080 ;
        RECT 4.400 411.720 345.600 411.760 ;
        RECT 4.400 410.360 346.000 411.720 ;
        RECT 4.000 409.040 346.000 410.360 ;
        RECT 4.400 407.680 346.000 409.040 ;
        RECT 4.400 407.640 345.600 407.680 ;
        RECT 4.000 406.320 345.600 407.640 ;
        RECT 4.400 406.280 345.600 406.320 ;
        RECT 4.400 404.920 346.000 406.280 ;
        RECT 4.000 403.600 346.000 404.920 ;
        RECT 4.400 402.240 346.000 403.600 ;
        RECT 4.400 402.200 345.600 402.240 ;
        RECT 4.000 400.880 345.600 402.200 ;
        RECT 4.400 400.840 345.600 400.880 ;
        RECT 4.400 399.480 346.000 400.840 ;
        RECT 4.000 398.160 346.000 399.480 ;
        RECT 4.400 396.760 346.000 398.160 ;
        RECT 4.000 396.120 346.000 396.760 ;
        RECT 4.000 395.440 345.600 396.120 ;
        RECT 4.400 394.720 345.600 395.440 ;
        RECT 4.400 394.040 346.000 394.720 ;
        RECT 4.000 392.720 346.000 394.040 ;
        RECT 4.400 391.320 346.000 392.720 ;
        RECT 4.000 390.680 346.000 391.320 ;
        RECT 4.000 390.000 345.600 390.680 ;
        RECT 4.400 389.280 345.600 390.000 ;
        RECT 4.400 388.600 346.000 389.280 ;
        RECT 4.000 387.280 346.000 388.600 ;
        RECT 4.400 385.880 346.000 387.280 ;
        RECT 4.000 385.240 346.000 385.880 ;
        RECT 4.000 384.560 345.600 385.240 ;
        RECT 4.400 383.840 345.600 384.560 ;
        RECT 4.400 383.160 346.000 383.840 ;
        RECT 4.000 381.840 346.000 383.160 ;
        RECT 4.400 380.440 346.000 381.840 ;
        RECT 4.000 379.800 346.000 380.440 ;
        RECT 4.000 379.120 345.600 379.800 ;
        RECT 4.400 378.400 345.600 379.120 ;
        RECT 4.400 377.720 346.000 378.400 ;
        RECT 4.000 376.400 346.000 377.720 ;
        RECT 4.400 375.000 346.000 376.400 ;
        RECT 4.000 373.680 346.000 375.000 ;
        RECT 4.400 372.280 345.600 373.680 ;
        RECT 4.000 370.960 346.000 372.280 ;
        RECT 4.400 369.560 346.000 370.960 ;
        RECT 4.000 368.240 346.000 369.560 ;
        RECT 4.000 367.560 345.600 368.240 ;
        RECT 4.400 366.840 345.600 367.560 ;
        RECT 4.400 366.160 346.000 366.840 ;
        RECT 4.000 364.840 346.000 366.160 ;
        RECT 4.400 363.440 346.000 364.840 ;
        RECT 4.000 362.800 346.000 363.440 ;
        RECT 4.000 362.120 345.600 362.800 ;
        RECT 4.400 361.400 345.600 362.120 ;
        RECT 4.400 360.720 346.000 361.400 ;
        RECT 4.000 359.400 346.000 360.720 ;
        RECT 4.400 358.000 346.000 359.400 ;
        RECT 4.000 357.360 346.000 358.000 ;
        RECT 4.000 356.680 345.600 357.360 ;
        RECT 4.400 355.960 345.600 356.680 ;
        RECT 4.400 355.280 346.000 355.960 ;
        RECT 4.000 353.960 346.000 355.280 ;
        RECT 4.400 352.560 346.000 353.960 ;
        RECT 4.000 351.240 346.000 352.560 ;
        RECT 4.400 349.840 345.600 351.240 ;
        RECT 4.000 348.520 346.000 349.840 ;
        RECT 4.400 347.120 346.000 348.520 ;
        RECT 4.000 345.800 346.000 347.120 ;
        RECT 4.400 344.400 345.600 345.800 ;
        RECT 4.000 343.080 346.000 344.400 ;
        RECT 4.400 341.680 346.000 343.080 ;
        RECT 4.000 340.360 346.000 341.680 ;
        RECT 4.400 338.960 345.600 340.360 ;
        RECT 4.000 337.640 346.000 338.960 ;
        RECT 4.400 336.240 346.000 337.640 ;
        RECT 4.000 334.920 346.000 336.240 ;
        RECT 4.400 333.520 345.600 334.920 ;
        RECT 4.000 332.200 346.000 333.520 ;
        RECT 4.400 330.800 346.000 332.200 ;
        RECT 4.000 329.480 346.000 330.800 ;
        RECT 4.400 328.800 346.000 329.480 ;
        RECT 4.400 328.080 345.600 328.800 ;
        RECT 4.000 327.400 345.600 328.080 ;
        RECT 4.000 326.760 346.000 327.400 ;
        RECT 4.400 325.360 346.000 326.760 ;
        RECT 4.000 324.040 346.000 325.360 ;
        RECT 4.400 323.360 346.000 324.040 ;
        RECT 4.400 322.640 345.600 323.360 ;
        RECT 4.000 321.960 345.600 322.640 ;
        RECT 4.000 321.320 346.000 321.960 ;
        RECT 4.400 319.920 346.000 321.320 ;
        RECT 4.000 318.600 346.000 319.920 ;
        RECT 4.400 317.920 346.000 318.600 ;
        RECT 4.400 317.200 345.600 317.920 ;
        RECT 4.000 316.520 345.600 317.200 ;
        RECT 4.000 315.880 346.000 316.520 ;
        RECT 4.400 314.480 346.000 315.880 ;
        RECT 4.000 313.160 346.000 314.480 ;
        RECT 4.400 312.480 346.000 313.160 ;
        RECT 4.400 311.760 345.600 312.480 ;
        RECT 4.000 311.080 345.600 311.760 ;
        RECT 4.000 310.440 346.000 311.080 ;
        RECT 4.400 309.040 346.000 310.440 ;
        RECT 4.000 307.040 346.000 309.040 ;
        RECT 4.400 306.360 346.000 307.040 ;
        RECT 4.400 305.640 345.600 306.360 ;
        RECT 4.000 304.960 345.600 305.640 ;
        RECT 4.000 304.320 346.000 304.960 ;
        RECT 4.400 302.920 346.000 304.320 ;
        RECT 4.000 301.600 346.000 302.920 ;
        RECT 4.400 300.920 346.000 301.600 ;
        RECT 4.400 300.200 345.600 300.920 ;
        RECT 4.000 299.520 345.600 300.200 ;
        RECT 4.000 298.880 346.000 299.520 ;
        RECT 4.400 297.480 346.000 298.880 ;
        RECT 4.000 296.160 346.000 297.480 ;
        RECT 4.400 295.480 346.000 296.160 ;
        RECT 4.400 294.760 345.600 295.480 ;
        RECT 4.000 294.080 345.600 294.760 ;
        RECT 4.000 293.440 346.000 294.080 ;
        RECT 4.400 292.040 346.000 293.440 ;
        RECT 4.000 290.720 346.000 292.040 ;
        RECT 4.400 290.040 346.000 290.720 ;
        RECT 4.400 289.320 345.600 290.040 ;
        RECT 4.000 288.640 345.600 289.320 ;
        RECT 4.000 288.000 346.000 288.640 ;
        RECT 4.400 286.600 346.000 288.000 ;
        RECT 4.000 285.280 346.000 286.600 ;
        RECT 4.400 283.920 346.000 285.280 ;
        RECT 4.400 283.880 345.600 283.920 ;
        RECT 4.000 282.560 345.600 283.880 ;
        RECT 4.400 282.520 345.600 282.560 ;
        RECT 4.400 281.160 346.000 282.520 ;
        RECT 4.000 279.840 346.000 281.160 ;
        RECT 4.400 278.480 346.000 279.840 ;
        RECT 4.400 278.440 345.600 278.480 ;
        RECT 4.000 277.120 345.600 278.440 ;
        RECT 4.400 277.080 345.600 277.120 ;
        RECT 4.400 275.720 346.000 277.080 ;
        RECT 4.000 274.400 346.000 275.720 ;
        RECT 4.400 273.040 346.000 274.400 ;
        RECT 4.400 273.000 345.600 273.040 ;
        RECT 4.000 271.680 345.600 273.000 ;
        RECT 4.400 271.640 345.600 271.680 ;
        RECT 4.400 270.280 346.000 271.640 ;
        RECT 4.000 268.960 346.000 270.280 ;
        RECT 4.400 267.560 346.000 268.960 ;
        RECT 4.000 266.920 346.000 267.560 ;
        RECT 4.000 266.240 345.600 266.920 ;
        RECT 4.400 265.520 345.600 266.240 ;
        RECT 4.400 264.840 346.000 265.520 ;
        RECT 4.000 263.520 346.000 264.840 ;
        RECT 4.400 262.120 346.000 263.520 ;
        RECT 4.000 261.480 346.000 262.120 ;
        RECT 4.000 260.800 345.600 261.480 ;
        RECT 4.400 260.080 345.600 260.800 ;
        RECT 4.400 259.400 346.000 260.080 ;
        RECT 4.000 258.080 346.000 259.400 ;
        RECT 4.400 256.680 346.000 258.080 ;
        RECT 4.000 256.040 346.000 256.680 ;
        RECT 4.000 255.360 345.600 256.040 ;
        RECT 4.400 254.640 345.600 255.360 ;
        RECT 4.400 253.960 346.000 254.640 ;
        RECT 4.000 252.640 346.000 253.960 ;
        RECT 4.400 251.240 346.000 252.640 ;
        RECT 4.000 250.600 346.000 251.240 ;
        RECT 4.000 249.920 345.600 250.600 ;
        RECT 4.400 249.200 345.600 249.920 ;
        RECT 4.400 248.520 346.000 249.200 ;
        RECT 4.000 247.200 346.000 248.520 ;
        RECT 4.400 245.800 346.000 247.200 ;
        RECT 4.000 244.480 346.000 245.800 ;
        RECT 4.000 243.800 345.600 244.480 ;
        RECT 4.400 243.080 345.600 243.800 ;
        RECT 4.400 242.400 346.000 243.080 ;
        RECT 4.000 241.080 346.000 242.400 ;
        RECT 4.400 239.680 346.000 241.080 ;
        RECT 4.000 239.040 346.000 239.680 ;
        RECT 4.000 238.360 345.600 239.040 ;
        RECT 4.400 237.640 345.600 238.360 ;
        RECT 4.400 236.960 346.000 237.640 ;
        RECT 4.000 235.640 346.000 236.960 ;
        RECT 4.400 234.240 346.000 235.640 ;
        RECT 4.000 233.600 346.000 234.240 ;
        RECT 4.000 232.920 345.600 233.600 ;
        RECT 4.400 232.200 345.600 232.920 ;
        RECT 4.400 231.520 346.000 232.200 ;
        RECT 4.000 230.200 346.000 231.520 ;
        RECT 4.400 228.800 346.000 230.200 ;
        RECT 4.000 228.160 346.000 228.800 ;
        RECT 4.000 227.480 345.600 228.160 ;
        RECT 4.400 226.760 345.600 227.480 ;
        RECT 4.400 226.080 346.000 226.760 ;
        RECT 4.000 224.760 346.000 226.080 ;
        RECT 4.400 223.360 346.000 224.760 ;
        RECT 4.000 222.040 346.000 223.360 ;
        RECT 4.400 220.640 345.600 222.040 ;
        RECT 4.000 219.320 346.000 220.640 ;
        RECT 4.400 217.920 346.000 219.320 ;
        RECT 4.000 216.600 346.000 217.920 ;
        RECT 4.400 215.200 345.600 216.600 ;
        RECT 4.000 213.880 346.000 215.200 ;
        RECT 4.400 212.480 346.000 213.880 ;
        RECT 4.000 211.160 346.000 212.480 ;
        RECT 4.400 209.760 345.600 211.160 ;
        RECT 4.000 208.440 346.000 209.760 ;
        RECT 4.400 207.040 346.000 208.440 ;
        RECT 4.000 205.720 346.000 207.040 ;
        RECT 4.400 204.320 345.600 205.720 ;
        RECT 4.000 203.000 346.000 204.320 ;
        RECT 4.400 201.600 346.000 203.000 ;
        RECT 4.000 200.280 346.000 201.600 ;
        RECT 4.400 199.600 346.000 200.280 ;
        RECT 4.400 198.880 345.600 199.600 ;
        RECT 4.000 198.200 345.600 198.880 ;
        RECT 4.000 197.560 346.000 198.200 ;
        RECT 4.400 196.160 346.000 197.560 ;
        RECT 4.000 194.840 346.000 196.160 ;
        RECT 4.400 194.160 346.000 194.840 ;
        RECT 4.400 193.440 345.600 194.160 ;
        RECT 4.000 192.760 345.600 193.440 ;
        RECT 4.000 192.120 346.000 192.760 ;
        RECT 4.400 190.720 346.000 192.120 ;
        RECT 4.000 189.400 346.000 190.720 ;
        RECT 4.400 188.720 346.000 189.400 ;
        RECT 4.400 188.000 345.600 188.720 ;
        RECT 4.000 187.320 345.600 188.000 ;
        RECT 4.000 186.680 346.000 187.320 ;
        RECT 4.400 185.280 346.000 186.680 ;
        RECT 4.000 183.280 346.000 185.280 ;
        RECT 4.400 181.880 345.600 183.280 ;
        RECT 4.000 180.560 346.000 181.880 ;
        RECT 4.400 179.160 346.000 180.560 ;
        RECT 4.000 177.840 346.000 179.160 ;
        RECT 4.400 177.160 346.000 177.840 ;
        RECT 4.400 176.440 345.600 177.160 ;
        RECT 4.000 175.760 345.600 176.440 ;
        RECT 4.000 175.120 346.000 175.760 ;
        RECT 4.400 173.720 346.000 175.120 ;
        RECT 4.000 172.400 346.000 173.720 ;
        RECT 4.400 171.720 346.000 172.400 ;
        RECT 4.400 171.000 345.600 171.720 ;
        RECT 4.000 170.320 345.600 171.000 ;
        RECT 4.000 169.680 346.000 170.320 ;
        RECT 4.400 168.280 346.000 169.680 ;
        RECT 4.000 166.960 346.000 168.280 ;
        RECT 4.400 166.280 346.000 166.960 ;
        RECT 4.400 165.560 345.600 166.280 ;
        RECT 4.000 164.880 345.600 165.560 ;
        RECT 4.000 164.240 346.000 164.880 ;
        RECT 4.400 162.840 346.000 164.240 ;
        RECT 4.000 161.520 346.000 162.840 ;
        RECT 4.400 160.840 346.000 161.520 ;
        RECT 4.400 160.120 345.600 160.840 ;
        RECT 4.000 159.440 345.600 160.120 ;
        RECT 4.000 158.800 346.000 159.440 ;
        RECT 4.400 157.400 346.000 158.800 ;
        RECT 4.000 156.080 346.000 157.400 ;
        RECT 4.400 154.720 346.000 156.080 ;
        RECT 4.400 154.680 345.600 154.720 ;
        RECT 4.000 153.360 345.600 154.680 ;
        RECT 4.400 153.320 345.600 153.360 ;
        RECT 4.400 151.960 346.000 153.320 ;
        RECT 4.000 150.640 346.000 151.960 ;
        RECT 4.400 149.280 346.000 150.640 ;
        RECT 4.400 149.240 345.600 149.280 ;
        RECT 4.000 147.920 345.600 149.240 ;
        RECT 4.400 147.880 345.600 147.920 ;
        RECT 4.400 146.520 346.000 147.880 ;
        RECT 4.000 145.200 346.000 146.520 ;
        RECT 4.400 143.840 346.000 145.200 ;
        RECT 4.400 143.800 345.600 143.840 ;
        RECT 4.000 142.480 345.600 143.800 ;
        RECT 4.400 142.440 345.600 142.480 ;
        RECT 4.400 141.080 346.000 142.440 ;
        RECT 4.000 139.760 346.000 141.080 ;
        RECT 4.400 138.400 346.000 139.760 ;
        RECT 4.400 138.360 345.600 138.400 ;
        RECT 4.000 137.040 345.600 138.360 ;
        RECT 4.400 137.000 345.600 137.040 ;
        RECT 4.400 135.640 346.000 137.000 ;
        RECT 4.000 134.320 346.000 135.640 ;
        RECT 4.400 132.920 346.000 134.320 ;
        RECT 4.000 132.280 346.000 132.920 ;
        RECT 4.000 131.600 345.600 132.280 ;
        RECT 4.400 130.880 345.600 131.600 ;
        RECT 4.400 130.200 346.000 130.880 ;
        RECT 4.000 128.880 346.000 130.200 ;
        RECT 4.400 127.480 346.000 128.880 ;
        RECT 4.000 126.840 346.000 127.480 ;
        RECT 4.000 126.160 345.600 126.840 ;
        RECT 4.400 125.440 345.600 126.160 ;
        RECT 4.400 124.760 346.000 125.440 ;
        RECT 4.000 122.760 346.000 124.760 ;
        RECT 4.400 121.400 346.000 122.760 ;
        RECT 4.400 121.360 345.600 121.400 ;
        RECT 4.000 120.040 345.600 121.360 ;
        RECT 4.400 120.000 345.600 120.040 ;
        RECT 4.400 118.640 346.000 120.000 ;
        RECT 4.000 117.320 346.000 118.640 ;
        RECT 4.400 115.960 346.000 117.320 ;
        RECT 4.400 115.920 345.600 115.960 ;
        RECT 4.000 114.600 345.600 115.920 ;
        RECT 4.400 114.560 345.600 114.600 ;
        RECT 4.400 113.200 346.000 114.560 ;
        RECT 4.000 111.880 346.000 113.200 ;
        RECT 4.400 110.480 346.000 111.880 ;
        RECT 4.000 109.840 346.000 110.480 ;
        RECT 4.000 109.160 345.600 109.840 ;
        RECT 4.400 108.440 345.600 109.160 ;
        RECT 4.400 107.760 346.000 108.440 ;
        RECT 4.000 106.440 346.000 107.760 ;
        RECT 4.400 105.040 346.000 106.440 ;
        RECT 4.000 104.400 346.000 105.040 ;
        RECT 4.000 103.720 345.600 104.400 ;
        RECT 4.400 103.000 345.600 103.720 ;
        RECT 4.400 102.320 346.000 103.000 ;
        RECT 4.000 101.000 346.000 102.320 ;
        RECT 4.400 99.600 346.000 101.000 ;
        RECT 4.000 98.960 346.000 99.600 ;
        RECT 4.000 98.280 345.600 98.960 ;
        RECT 4.400 97.560 345.600 98.280 ;
        RECT 4.400 96.880 346.000 97.560 ;
        RECT 4.000 95.560 346.000 96.880 ;
        RECT 4.400 94.160 346.000 95.560 ;
        RECT 4.000 93.520 346.000 94.160 ;
        RECT 4.000 92.840 345.600 93.520 ;
        RECT 4.400 92.120 345.600 92.840 ;
        RECT 4.400 91.440 346.000 92.120 ;
        RECT 4.000 90.120 346.000 91.440 ;
        RECT 4.400 88.720 346.000 90.120 ;
        RECT 4.000 87.400 346.000 88.720 ;
        RECT 4.400 86.000 345.600 87.400 ;
        RECT 4.000 84.680 346.000 86.000 ;
        RECT 4.400 83.280 346.000 84.680 ;
        RECT 4.000 81.960 346.000 83.280 ;
        RECT 4.400 80.560 345.600 81.960 ;
        RECT 4.000 79.240 346.000 80.560 ;
        RECT 4.400 77.840 346.000 79.240 ;
        RECT 4.000 76.520 346.000 77.840 ;
        RECT 4.400 75.120 345.600 76.520 ;
        RECT 4.000 73.800 346.000 75.120 ;
        RECT 4.400 72.400 346.000 73.800 ;
        RECT 4.000 71.080 346.000 72.400 ;
        RECT 4.400 69.680 345.600 71.080 ;
        RECT 4.000 68.360 346.000 69.680 ;
        RECT 4.400 66.960 346.000 68.360 ;
        RECT 4.000 65.640 346.000 66.960 ;
        RECT 4.400 64.960 346.000 65.640 ;
        RECT 4.400 64.240 345.600 64.960 ;
        RECT 4.000 63.560 345.600 64.240 ;
        RECT 4.000 62.240 346.000 63.560 ;
        RECT 4.400 60.840 346.000 62.240 ;
        RECT 4.000 59.520 346.000 60.840 ;
        RECT 4.400 58.120 345.600 59.520 ;
        RECT 4.000 56.800 346.000 58.120 ;
        RECT 4.400 55.400 346.000 56.800 ;
        RECT 4.000 54.080 346.000 55.400 ;
        RECT 4.400 52.680 345.600 54.080 ;
        RECT 4.000 51.360 346.000 52.680 ;
        RECT 4.400 49.960 346.000 51.360 ;
        RECT 4.000 48.640 346.000 49.960 ;
        RECT 4.400 47.240 345.600 48.640 ;
        RECT 4.000 45.920 346.000 47.240 ;
        RECT 4.400 44.520 346.000 45.920 ;
        RECT 4.000 43.200 346.000 44.520 ;
        RECT 4.400 42.520 346.000 43.200 ;
        RECT 4.400 41.800 345.600 42.520 ;
        RECT 4.000 41.120 345.600 41.800 ;
        RECT 4.000 40.480 346.000 41.120 ;
        RECT 4.400 39.080 346.000 40.480 ;
        RECT 4.000 37.760 346.000 39.080 ;
        RECT 4.400 37.080 346.000 37.760 ;
        RECT 4.400 36.360 345.600 37.080 ;
        RECT 4.000 35.680 345.600 36.360 ;
        RECT 4.000 35.040 346.000 35.680 ;
        RECT 4.400 33.640 346.000 35.040 ;
        RECT 4.000 32.320 346.000 33.640 ;
        RECT 4.400 31.640 346.000 32.320 ;
        RECT 4.400 30.920 345.600 31.640 ;
        RECT 4.000 30.240 345.600 30.920 ;
        RECT 4.000 29.600 346.000 30.240 ;
        RECT 4.400 28.200 346.000 29.600 ;
        RECT 4.000 26.880 346.000 28.200 ;
        RECT 4.400 26.200 346.000 26.880 ;
        RECT 4.400 25.480 345.600 26.200 ;
        RECT 4.000 24.800 345.600 25.480 ;
        RECT 4.000 24.160 346.000 24.800 ;
        RECT 4.400 22.760 346.000 24.160 ;
        RECT 4.000 21.440 346.000 22.760 ;
        RECT 4.400 20.080 346.000 21.440 ;
        RECT 4.400 20.040 345.600 20.080 ;
        RECT 4.000 18.720 345.600 20.040 ;
        RECT 4.400 18.680 345.600 18.720 ;
        RECT 4.400 17.320 346.000 18.680 ;
        RECT 4.000 16.000 346.000 17.320 ;
        RECT 4.400 14.640 346.000 16.000 ;
        RECT 4.400 14.600 345.600 14.640 ;
        RECT 4.000 13.280 345.600 14.600 ;
        RECT 4.400 13.240 345.600 13.280 ;
        RECT 4.400 11.880 346.000 13.240 ;
        RECT 4.000 10.560 346.000 11.880 ;
        RECT 4.400 9.200 346.000 10.560 ;
        RECT 4.400 9.160 345.600 9.200 ;
        RECT 4.000 7.840 345.600 9.160 ;
        RECT 4.400 7.800 345.600 7.840 ;
        RECT 4.400 6.440 346.000 7.800 ;
        RECT 4.000 5.120 346.000 6.440 ;
        RECT 4.400 3.760 346.000 5.120 ;
        RECT 4.400 3.720 345.600 3.760 ;
        RECT 4.000 2.400 345.600 3.720 ;
        RECT 4.400 2.360 345.600 2.400 ;
        RECT 4.400 1.535 346.000 2.360 ;
      LAYER met4 ;
        RECT 4.895 19.895 20.640 1087.145 ;
        RECT 23.040 19.895 97.440 1087.145 ;
        RECT 99.840 19.895 174.240 1087.145 ;
        RECT 176.640 19.895 251.040 1087.145 ;
        RECT 253.440 19.895 295.945 1087.145 ;
  END
END WishboneInterconnect
END LIBRARY

