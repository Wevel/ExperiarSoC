VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Art
  CLASS BLOCK ;
  FOREIGN Art ;
  ORIGIN -0.200 0.000 ;
  SIZE 302.920 BY 750.000 ;
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.20000 0.00000 1.80000 750.00000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 298.20000 0.00000 299.80000 750.00000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.000 30.000 105.000 70.000 ;
        RECT 5.000 5.000 25.000 25.000 ;
      LAYER met1 ;
        RECT 85.000 60.000 105.000 70.120 ;
        RECT 65.000 50.000 105.000 60.000 ;
        RECT 45.000 40.000 105.000 50.000 ;
        RECT 25.000 30.120 105.000 40.000 ;
        RECT 25.000 30.000 85.000 30.120 ;
        RECT 25.000 5.000 45.000 25.000 ;
      LAYER met2 ;
        RECT 45.000 60.000 65.000 70.000 ;
        RECT 25.000 50.000 45.000 60.000 ;
        RECT 85.000 50.000 105.000 60.000 ;
        RECT 5.000 40.000 25.000 50.000 ;
        RECT 65.000 40.000 105.000 50.000 ;
        RECT 45.000 30.000 105.000 40.000 ;
        RECT 45.000 5.000 65.000 25.000 ;
      LAYER met3 ;
        RECT 25.000 60.000 45.000 70.000 ;
        RECT 5.000 50.000 25.000 60.000 ;
        RECT 85.000 40.000 105.000 50.000 ;
        RECT 65.000 30.000 105.000 40.000 ;
        RECT 65.000 5.000 85.000 25.000 ;
      LAYER met4 ;
        RECT 0.200 0.000 1.800 750.000 ;
        RECT 69.830 739.290 75.830 741.290 ;
        RECT 69.830 737.290 71.830 739.290 ;
        RECT 67.830 735.290 71.830 737.290 ;
        RECT 73.830 737.290 75.830 739.290 ;
        RECT 219.830 739.290 225.830 741.290 ;
        RECT 219.830 737.290 221.830 739.290 ;
        RECT 73.830 735.290 77.830 737.290 ;
        RECT 67.830 731.290 69.830 735.290 ;
        RECT 65.830 729.290 69.830 731.290 ;
        RECT 75.830 731.290 77.830 735.290 ;
        RECT 217.830 735.290 221.830 737.290 ;
        RECT 223.830 737.290 225.830 739.290 ;
        RECT 223.830 735.290 227.830 737.290 ;
        RECT 217.830 731.290 219.830 735.290 ;
        RECT 75.830 729.290 79.830 731.290 ;
        RECT 65.830 725.290 67.830 729.290 ;
        RECT 63.830 723.290 67.830 725.290 ;
        RECT 69.830 723.290 73.830 727.290 ;
        RECT 77.830 725.290 79.830 729.290 ;
        RECT 215.830 729.290 219.830 731.290 ;
        RECT 225.830 731.290 227.830 735.290 ;
        RECT 225.830 729.290 229.830 731.290 ;
        RECT 215.830 725.290 217.830 729.290 ;
        RECT 77.830 723.290 81.830 725.290 ;
        RECT 63.830 719.290 65.830 723.290 ;
        RECT 61.830 717.290 65.830 719.290 ;
        RECT 67.830 721.290 73.830 723.290 ;
        RECT 79.830 721.290 81.830 723.290 ;
        RECT 213.830 723.290 217.830 725.290 ;
        RECT 219.830 723.290 223.830 727.290 ;
        RECT 227.830 725.290 229.830 729.290 ;
        RECT 227.830 723.290 231.830 725.290 ;
        RECT 67.830 719.290 75.830 721.290 ;
        RECT 79.830 719.290 83.830 721.290 ;
        RECT 213.830 719.290 215.830 723.290 ;
        RECT 67.830 717.290 77.830 719.290 ;
        RECT 61.830 715.290 63.830 717.290 ;
        RECT 59.830 713.290 63.830 715.290 ;
        RECT 65.830 713.290 73.830 717.290 ;
        RECT 59.830 709.290 61.830 713.290 ;
        RECT 57.830 707.290 61.830 709.290 ;
        RECT 63.830 709.290 73.830 713.290 ;
        RECT 75.830 713.290 79.830 717.290 ;
        RECT 81.830 715.290 83.830 719.290 ;
        RECT 211.830 717.290 215.830 719.290 ;
        RECT 217.830 721.290 223.830 723.290 ;
        RECT 229.830 721.290 231.830 723.290 ;
        RECT 217.830 719.290 225.830 721.290 ;
        RECT 229.830 719.290 233.830 721.290 ;
        RECT 217.830 717.290 227.830 719.290 ;
        RECT 211.830 715.290 213.830 717.290 ;
        RECT 81.830 713.290 85.830 715.290 ;
        RECT 75.830 709.290 81.830 713.290 ;
        RECT 63.830 707.290 75.830 709.290 ;
        RECT 57.830 705.290 59.830 707.290 ;
        RECT 51.830 703.290 59.830 705.290 ;
        RECT 61.830 703.290 75.830 707.290 ;
        RECT 77.830 707.290 81.830 709.290 ;
        RECT 83.830 709.290 85.830 713.290 ;
        RECT 209.830 713.290 213.830 715.290 ;
        RECT 215.830 713.290 223.830 717.290 ;
        RECT 209.830 709.290 211.830 713.290 ;
        RECT 83.830 707.290 87.830 709.290 ;
        RECT 77.830 705.290 83.830 707.290 ;
        RECT 77.830 703.290 79.830 705.290 ;
        RECT 85.830 703.290 87.830 707.290 ;
        RECT 207.830 707.290 211.830 709.290 ;
        RECT 213.830 709.290 223.830 713.290 ;
        RECT 225.830 713.290 229.830 717.290 ;
        RECT 231.830 715.290 233.830 719.290 ;
        RECT 231.830 713.290 235.830 715.290 ;
        RECT 225.830 709.290 231.830 713.290 ;
        RECT 213.830 707.290 225.830 709.290 ;
        RECT 207.830 705.290 209.830 707.290 ;
        RECT 201.830 703.290 209.830 705.290 ;
        RECT 211.830 703.290 225.830 707.290 ;
        RECT 227.830 707.290 231.830 709.290 ;
        RECT 233.830 709.290 235.830 713.290 ;
        RECT 233.830 707.290 237.830 709.290 ;
        RECT 227.830 705.290 233.830 707.290 ;
        RECT 227.830 703.290 229.830 705.290 ;
        RECT 235.830 703.290 237.830 707.290 ;
        RECT 41.830 701.290 53.830 703.290 ;
        RECT 61.830 701.290 77.830 703.290 ;
        RECT 79.830 701.290 83.830 703.290 ;
        RECT 85.830 701.290 95.830 703.290 ;
        RECT 191.830 701.290 203.830 703.290 ;
        RECT 211.830 701.290 227.830 703.290 ;
        RECT 229.830 701.290 233.830 703.290 ;
        RECT 235.830 701.290 245.830 703.290 ;
        RECT 35.830 699.290 43.830 701.290 ;
        RECT 53.830 699.290 57.830 701.290 ;
        RECT 35.830 695.290 37.830 699.290 ;
        RECT 43.830 697.290 57.830 699.290 ;
        RECT 59.830 697.290 85.830 701.290 ;
        RECT 93.830 699.290 103.830 701.290 ;
        RECT 185.830 699.290 193.830 701.290 ;
        RECT 203.830 699.290 207.830 701.290 ;
        RECT 87.830 697.290 89.830 699.290 ;
        RECT 101.830 697.290 111.830 699.290 ;
        RECT 43.830 695.290 59.830 697.290 ;
        RECT 69.830 695.290 81.830 697.290 ;
        RECT 85.830 695.290 93.830 697.290 ;
        RECT 109.830 695.290 115.830 697.290 ;
        RECT 35.830 693.290 43.830 695.290 ;
        RECT 53.830 693.290 69.830 695.290 ;
        RECT 81.830 693.290 99.830 695.290 ;
        RECT 113.830 693.290 115.830 695.290 ;
        RECT 185.830 695.290 187.830 699.290 ;
        RECT 193.830 697.290 207.830 699.290 ;
        RECT 209.830 697.290 235.830 701.290 ;
        RECT 243.830 699.290 253.830 701.290 ;
        RECT 237.830 697.290 239.830 699.290 ;
        RECT 251.830 697.290 261.830 699.290 ;
        RECT 193.830 695.290 209.830 697.290 ;
        RECT 219.830 695.290 231.830 697.290 ;
        RECT 235.830 695.290 243.830 697.290 ;
        RECT 259.830 695.290 265.830 697.290 ;
        RECT 185.830 693.290 193.830 695.290 ;
        RECT 203.830 693.290 219.830 695.290 ;
        RECT 231.830 693.290 249.830 695.290 ;
        RECT 263.830 693.290 265.830 695.290 ;
        RECT 41.830 691.290 53.830 693.290 ;
        RECT 63.830 691.290 103.830 693.290 ;
        RECT 111.830 691.290 115.830 693.290 ;
        RECT 191.830 691.290 203.830 693.290 ;
        RECT 213.830 691.290 253.830 693.290 ;
        RECT 261.830 691.290 265.830 693.290 ;
        RECT 51.830 689.290 63.830 691.290 ;
        RECT 73.830 689.290 101.830 691.290 ;
        RECT 109.830 689.290 113.830 691.290 ;
        RECT 201.830 689.290 213.830 691.290 ;
        RECT 223.830 689.290 251.830 691.290 ;
        RECT 259.830 689.290 263.830 691.290 ;
        RECT 53.830 687.290 55.830 689.290 ;
        RECT 51.830 685.290 55.830 687.290 ;
        RECT 57.830 687.290 73.830 689.290 ;
        RECT 83.830 687.290 93.830 689.290 ;
        RECT 101.830 687.290 111.830 689.290 ;
        RECT 203.830 687.290 205.830 689.290 ;
        RECT 57.830 685.290 83.830 687.290 ;
        RECT 93.830 685.290 103.830 687.290 ;
        RECT 201.830 685.290 205.830 687.290 ;
        RECT 207.830 687.290 223.830 689.290 ;
        RECT 233.830 687.290 243.830 689.290 ;
        RECT 251.830 687.290 261.830 689.290 ;
        RECT 207.830 685.290 233.830 687.290 ;
        RECT 243.830 685.290 253.830 687.290 ;
        RECT 51.830 679.290 53.830 685.290 ;
        RECT 55.830 683.290 73.830 685.290 ;
        RECT 83.830 683.290 95.830 685.290 ;
        RECT 55.830 681.290 71.830 683.290 ;
        RECT 57.830 679.290 71.830 681.290 ;
        RECT 73.830 681.290 77.830 683.290 ;
        RECT 81.830 681.290 83.830 683.290 ;
        RECT 87.830 681.290 89.830 683.290 ;
        RECT 93.830 681.290 95.830 683.290 ;
        RECT 103.830 681.290 109.830 683.290 ;
        RECT 73.830 679.290 75.830 681.290 ;
        RECT 87.830 679.290 95.830 681.290 ;
        RECT 101.830 679.290 105.830 681.290 ;
        RECT 107.830 679.290 109.830 681.290 ;
        RECT 201.830 679.290 203.830 685.290 ;
        RECT 205.830 683.290 223.830 685.290 ;
        RECT 233.830 683.290 245.830 685.290 ;
        RECT 205.830 681.290 221.830 683.290 ;
        RECT 207.830 679.290 221.830 681.290 ;
        RECT 223.830 681.290 227.830 683.290 ;
        RECT 231.830 681.290 233.830 683.290 ;
        RECT 237.830 681.290 239.830 683.290 ;
        RECT 243.830 681.290 245.830 683.290 ;
        RECT 253.830 681.290 259.830 683.290 ;
        RECT 223.830 679.290 225.830 681.290 ;
        RECT 237.830 679.290 245.830 681.290 ;
        RECT 251.830 679.290 255.830 681.290 ;
        RECT 257.830 679.290 259.830 681.290 ;
        RECT 49.830 677.290 55.830 679.290 ;
        RECT 47.830 675.290 51.830 677.290 ;
        RECT 53.830 675.290 59.830 677.290 ;
        RECT 61.830 675.290 71.830 679.290 ;
        RECT 75.830 677.290 77.830 679.290 ;
        RECT 87.830 677.290 91.830 679.290 ;
        RECT 97.830 677.290 103.830 679.290 ;
        RECT 105.830 677.290 109.830 679.290 ;
        RECT 199.830 677.290 205.830 679.290 ;
        RECT 85.830 675.290 91.830 677.290 ;
        RECT 93.830 675.290 99.830 677.290 ;
        RECT 45.830 673.290 49.830 675.290 ;
        RECT 51.830 673.290 61.830 675.290 ;
        RECT 65.830 673.290 73.830 675.290 ;
        RECT 79.830 673.290 95.830 675.290 ;
        RECT 99.830 673.290 103.830 675.290 ;
        RECT 45.830 667.290 47.830 673.290 ;
        RECT 43.830 665.290 47.830 667.290 ;
        RECT 49.830 671.290 63.830 673.290 ;
        RECT 67.830 671.290 73.830 673.290 ;
        RECT 83.830 671.290 91.830 673.290 ;
        RECT 95.830 671.290 105.830 673.290 ;
        RECT 107.830 671.290 109.830 677.290 ;
        RECT 197.830 675.290 201.830 677.290 ;
        RECT 203.830 675.290 209.830 677.290 ;
        RECT 211.830 675.290 221.830 679.290 ;
        RECT 225.830 677.290 227.830 679.290 ;
        RECT 237.830 677.290 241.830 679.290 ;
        RECT 247.830 677.290 253.830 679.290 ;
        RECT 255.830 677.290 259.830 679.290 ;
        RECT 235.830 675.290 241.830 677.290 ;
        RECT 243.830 675.290 249.830 677.290 ;
        RECT 49.830 669.290 67.830 671.290 ;
        RECT 69.830 669.290 73.830 671.290 ;
        RECT 81.830 669.290 87.830 671.290 ;
        RECT 91.830 669.290 101.830 671.290 ;
        RECT 105.830 669.290 109.830 671.290 ;
        RECT 195.830 673.290 199.830 675.290 ;
        RECT 201.830 673.290 211.830 675.290 ;
        RECT 215.830 673.290 223.830 675.290 ;
        RECT 229.830 673.290 245.830 675.290 ;
        RECT 249.830 673.290 253.830 675.290 ;
        RECT 49.830 667.290 69.830 669.290 ;
        RECT 77.830 667.290 83.830 669.290 ;
        RECT 87.830 667.290 99.830 669.290 ;
        RECT 49.830 665.290 89.830 667.290 ;
        RECT 97.830 665.290 99.830 667.290 ;
        RECT 101.830 667.290 107.830 669.290 ;
        RECT 195.830 667.290 197.830 673.290 ;
        RECT 101.830 665.290 103.830 667.290 ;
        RECT 43.830 645.290 45.830 665.290 ;
        RECT 47.830 663.290 63.830 665.290 ;
        RECT 65.830 663.290 67.830 665.290 ;
        RECT 71.830 663.290 83.830 665.290 ;
        RECT 47.830 661.290 61.830 663.290 ;
        RECT 63.830 661.290 65.830 663.290 ;
        RECT 67.830 661.290 71.830 663.290 ;
        RECT 77.830 661.290 81.830 663.290 ;
        RECT 83.830 661.290 85.830 663.290 ;
        RECT 99.830 661.290 103.830 665.290 ;
        RECT 47.830 659.290 63.830 661.290 ;
        RECT 65.830 659.290 67.830 661.290 ;
        RECT 47.830 657.290 61.830 659.290 ;
        RECT 63.830 657.290 67.830 659.290 ;
        RECT 71.830 659.290 81.830 661.290 ;
        RECT 85.830 659.290 103.830 661.290 ;
        RECT 193.830 665.290 197.830 667.290 ;
        RECT 199.830 671.290 213.830 673.290 ;
        RECT 217.830 671.290 223.830 673.290 ;
        RECT 233.830 671.290 241.830 673.290 ;
        RECT 245.830 671.290 255.830 673.290 ;
        RECT 257.830 671.290 259.830 677.290 ;
        RECT 199.830 669.290 217.830 671.290 ;
        RECT 219.830 669.290 223.830 671.290 ;
        RECT 231.830 669.290 237.830 671.290 ;
        RECT 241.830 669.290 251.830 671.290 ;
        RECT 255.830 669.290 259.830 671.290 ;
        RECT 199.830 667.290 219.830 669.290 ;
        RECT 227.830 667.290 233.830 669.290 ;
        RECT 237.830 667.290 249.830 669.290 ;
        RECT 199.830 665.290 239.830 667.290 ;
        RECT 247.830 665.290 249.830 667.290 ;
        RECT 251.830 667.290 257.830 669.290 ;
        RECT 251.830 665.290 253.830 667.290 ;
        RECT 71.830 657.290 73.830 659.290 ;
        RECT 79.830 657.290 83.830 659.290 ;
        RECT 87.830 657.290 89.830 659.290 ;
        RECT 101.830 657.290 105.830 659.290 ;
        RECT 47.830 655.290 63.830 657.290 ;
        RECT 65.830 655.290 67.830 657.290 ;
        RECT 73.830 655.290 77.830 657.290 ;
        RECT 47.830 653.290 65.830 655.290 ;
        RECT 67.830 653.290 69.830 655.290 ;
        RECT 75.830 653.290 77.830 655.290 ;
        RECT 79.830 655.290 81.830 657.290 ;
        RECT 79.830 653.290 83.830 655.290 ;
        RECT 85.830 653.290 87.830 657.290 ;
        RECT 103.830 655.290 107.830 657.290 ;
        RECT 99.830 653.290 103.830 655.290 ;
        RECT 47.830 651.290 63.830 653.290 ;
        RECT 69.830 651.290 71.830 653.290 ;
        RECT 77.830 651.290 85.830 653.290 ;
        RECT 87.830 651.290 91.830 653.290 ;
        RECT 95.830 651.290 101.830 653.290 ;
        RECT 105.830 651.290 107.830 655.290 ;
        RECT 47.830 649.290 65.830 651.290 ;
        RECT 71.830 649.290 73.830 651.290 ;
        RECT 81.830 649.290 87.830 651.290 ;
        RECT 91.830 649.290 95.830 651.290 ;
        RECT 101.830 649.290 107.830 651.290 ;
        RECT 47.830 647.290 63.830 649.290 ;
        RECT 73.830 647.290 75.830 649.290 ;
        RECT 83.830 647.290 91.830 649.290 ;
        RECT 95.830 647.290 103.830 649.290 ;
        RECT 47.830 645.290 61.830 647.290 ;
        RECT 63.830 645.290 65.830 647.290 ;
        RECT 75.830 645.290 79.830 647.290 ;
        RECT 89.830 645.290 97.830 647.290 ;
        RECT 193.830 645.290 195.830 665.290 ;
        RECT 197.830 663.290 213.830 665.290 ;
        RECT 215.830 663.290 217.830 665.290 ;
        RECT 221.830 663.290 233.830 665.290 ;
        RECT 197.830 661.290 211.830 663.290 ;
        RECT 213.830 661.290 215.830 663.290 ;
        RECT 217.830 661.290 221.830 663.290 ;
        RECT 227.830 661.290 231.830 663.290 ;
        RECT 233.830 661.290 235.830 663.290 ;
        RECT 249.830 661.290 253.830 665.290 ;
        RECT 197.830 659.290 213.830 661.290 ;
        RECT 215.830 659.290 217.830 661.290 ;
        RECT 197.830 657.290 211.830 659.290 ;
        RECT 213.830 657.290 217.830 659.290 ;
        RECT 221.830 659.290 231.830 661.290 ;
        RECT 235.830 659.290 253.830 661.290 ;
        RECT 221.830 657.290 223.830 659.290 ;
        RECT 229.830 657.290 233.830 659.290 ;
        RECT 237.830 657.290 239.830 659.290 ;
        RECT 251.830 657.290 255.830 659.290 ;
        RECT 197.830 655.290 213.830 657.290 ;
        RECT 215.830 655.290 217.830 657.290 ;
        RECT 223.830 655.290 227.830 657.290 ;
        RECT 197.830 653.290 215.830 655.290 ;
        RECT 217.830 653.290 219.830 655.290 ;
        RECT 225.830 653.290 227.830 655.290 ;
        RECT 229.830 655.290 231.830 657.290 ;
        RECT 229.830 653.290 233.830 655.290 ;
        RECT 235.830 653.290 237.830 657.290 ;
        RECT 253.830 655.290 257.830 657.290 ;
        RECT 249.830 653.290 253.830 655.290 ;
        RECT 197.830 651.290 213.830 653.290 ;
        RECT 219.830 651.290 221.830 653.290 ;
        RECT 227.830 651.290 235.830 653.290 ;
        RECT 237.830 651.290 241.830 653.290 ;
        RECT 245.830 651.290 251.830 653.290 ;
        RECT 255.830 651.290 257.830 655.290 ;
        RECT 197.830 649.290 215.830 651.290 ;
        RECT 221.830 649.290 223.830 651.290 ;
        RECT 231.830 649.290 237.830 651.290 ;
        RECT 241.830 649.290 245.830 651.290 ;
        RECT 251.830 649.290 257.830 651.290 ;
        RECT 197.830 647.290 213.830 649.290 ;
        RECT 223.830 647.290 225.830 649.290 ;
        RECT 233.830 647.290 241.830 649.290 ;
        RECT 245.830 647.290 253.830 649.290 ;
        RECT 197.830 645.290 211.830 647.290 ;
        RECT 213.830 645.290 215.830 647.290 ;
        RECT 225.830 645.290 229.830 647.290 ;
        RECT 239.830 645.290 247.830 647.290 ;
        RECT 43.830 643.290 47.830 645.290 ;
        RECT 45.830 627.290 47.830 643.290 ;
        RECT 49.830 641.290 59.830 645.290 ;
        RECT 61.830 643.290 63.830 645.290 ;
        RECT 65.830 643.290 67.830 645.290 ;
        RECT 79.830 643.290 93.830 645.290 ;
        RECT 193.830 643.290 197.830 645.290 ;
        RECT 63.830 641.290 65.830 643.290 ;
        RECT 79.830 641.290 89.830 643.290 ;
        RECT 49.830 639.290 63.830 641.290 ;
        RECT 65.830 639.290 67.830 641.290 ;
        RECT 81.830 639.290 89.830 641.290 ;
        RECT 49.830 637.290 61.830 639.290 ;
        RECT 63.830 637.290 65.830 639.290 ;
        RECT 49.830 635.290 63.830 637.290 ;
        RECT 65.830 635.290 67.830 637.290 ;
        RECT 81.830 635.290 91.830 639.290 ;
        RECT 49.830 633.290 65.830 635.290 ;
        RECT 49.830 631.290 63.830 633.290 ;
        RECT 65.830 631.290 67.830 633.290 ;
        RECT 83.830 631.290 91.830 635.290 ;
        RECT 49.830 629.290 65.830 631.290 ;
        RECT 49.830 627.290 63.830 629.290 ;
        RECT 65.830 627.290 67.830 629.290 ;
        RECT 85.830 627.290 91.830 631.290 ;
        RECT 45.830 625.290 49.830 627.290 ;
        RECT 51.830 625.290 65.830 627.290 ;
        RECT 83.830 625.290 85.830 627.290 ;
        RECT 89.830 625.290 91.830 627.290 ;
        RECT 195.830 627.290 197.830 643.290 ;
        RECT 199.830 641.290 209.830 645.290 ;
        RECT 211.830 643.290 213.830 645.290 ;
        RECT 215.830 643.290 217.830 645.290 ;
        RECT 229.830 643.290 243.830 645.290 ;
        RECT 213.830 641.290 215.830 643.290 ;
        RECT 229.830 641.290 239.830 643.290 ;
        RECT 199.830 639.290 213.830 641.290 ;
        RECT 215.830 639.290 217.830 641.290 ;
        RECT 231.830 639.290 239.830 641.290 ;
        RECT 199.830 637.290 211.830 639.290 ;
        RECT 213.830 637.290 215.830 639.290 ;
        RECT 199.830 635.290 213.830 637.290 ;
        RECT 215.830 635.290 217.830 637.290 ;
        RECT 231.830 635.290 241.830 639.290 ;
        RECT 199.830 633.290 215.830 635.290 ;
        RECT 199.830 631.290 213.830 633.290 ;
        RECT 215.830 631.290 217.830 633.290 ;
        RECT 233.830 631.290 241.830 635.290 ;
        RECT 199.830 629.290 215.830 631.290 ;
        RECT 199.830 627.290 213.830 629.290 ;
        RECT 215.830 627.290 217.830 629.290 ;
        RECT 235.830 627.290 241.830 631.290 ;
        RECT 195.830 625.290 199.830 627.290 ;
        RECT 201.830 625.290 215.830 627.290 ;
        RECT 233.830 625.290 235.830 627.290 ;
        RECT 239.830 625.290 241.830 627.290 ;
        RECT 47.830 623.290 49.830 625.290 ;
        RECT 55.830 623.290 63.830 625.290 ;
        RECT 65.830 623.290 67.830 625.290 ;
        RECT 69.830 623.290 71.830 625.290 ;
        RECT 73.830 623.290 75.830 625.290 ;
        RECT 77.830 623.290 79.830 625.290 ;
        RECT 81.830 623.290 83.830 625.290 ;
        RECT 85.830 623.290 91.830 625.290 ;
        RECT 197.830 623.290 199.830 625.290 ;
        RECT 205.830 623.290 213.830 625.290 ;
        RECT 215.830 623.290 217.830 625.290 ;
        RECT 219.830 623.290 221.830 625.290 ;
        RECT 223.830 623.290 225.830 625.290 ;
        RECT 227.830 623.290 229.830 625.290 ;
        RECT 231.830 623.290 233.830 625.290 ;
        RECT 235.830 623.290 241.830 625.290 ;
        RECT 47.830 621.290 55.830 623.290 ;
        RECT 63.830 621.290 65.830 623.290 ;
        RECT 67.830 621.290 69.830 623.290 ;
        RECT 71.830 621.290 73.830 623.290 ;
        RECT 75.830 621.290 77.830 623.290 ;
        RECT 79.830 621.290 89.830 623.290 ;
        RECT 197.830 621.290 205.830 623.290 ;
        RECT 213.830 621.290 215.830 623.290 ;
        RECT 217.830 621.290 219.830 623.290 ;
        RECT 221.830 621.290 223.830 623.290 ;
        RECT 225.830 621.290 227.830 623.290 ;
        RECT 229.830 621.290 239.830 623.290 ;
        RECT 53.830 619.290 71.830 621.290 ;
        RECT 73.830 619.290 87.830 621.290 ;
        RECT 203.830 619.290 221.830 621.290 ;
        RECT 223.830 619.290 237.830 621.290 ;
        RECT 69.830 617.290 75.830 619.290 ;
        RECT 219.830 617.290 225.830 619.290 ;
        RECT 69.830 589.290 75.830 591.290 ;
        RECT 69.830 587.290 71.830 589.290 ;
        RECT 67.830 585.290 71.830 587.290 ;
        RECT 73.830 587.290 75.830 589.290 ;
        RECT 219.830 589.290 225.830 591.290 ;
        RECT 219.830 587.290 221.830 589.290 ;
        RECT 73.830 585.290 77.830 587.290 ;
        RECT 67.830 581.290 69.830 585.290 ;
        RECT 65.830 579.290 69.830 581.290 ;
        RECT 75.830 581.290 77.830 585.290 ;
        RECT 217.830 585.290 221.830 587.290 ;
        RECT 223.830 587.290 225.830 589.290 ;
        RECT 223.830 585.290 227.830 587.290 ;
        RECT 217.830 581.290 219.830 585.290 ;
        RECT 75.830 579.290 79.830 581.290 ;
        RECT 65.830 575.290 67.830 579.290 ;
        RECT 63.830 573.290 67.830 575.290 ;
        RECT 69.830 573.290 73.830 577.290 ;
        RECT 77.830 575.290 79.830 579.290 ;
        RECT 215.830 579.290 219.830 581.290 ;
        RECT 225.830 581.290 227.830 585.290 ;
        RECT 225.830 579.290 229.830 581.290 ;
        RECT 215.830 575.290 217.830 579.290 ;
        RECT 77.830 573.290 81.830 575.290 ;
        RECT 63.830 569.290 65.830 573.290 ;
        RECT 61.830 567.290 65.830 569.290 ;
        RECT 67.830 571.290 73.830 573.290 ;
        RECT 79.830 571.290 81.830 573.290 ;
        RECT 213.830 573.290 217.830 575.290 ;
        RECT 219.830 573.290 223.830 577.290 ;
        RECT 227.830 575.290 229.830 579.290 ;
        RECT 227.830 573.290 231.830 575.290 ;
        RECT 67.830 569.290 75.830 571.290 ;
        RECT 79.830 569.290 83.830 571.290 ;
        RECT 213.830 569.290 215.830 573.290 ;
        RECT 67.830 567.290 77.830 569.290 ;
        RECT 61.830 565.290 63.830 567.290 ;
        RECT 59.830 563.290 63.830 565.290 ;
        RECT 65.830 563.290 73.830 567.290 ;
        RECT 59.830 559.290 61.830 563.290 ;
        RECT 57.830 557.290 61.830 559.290 ;
        RECT 63.830 559.290 73.830 563.290 ;
        RECT 75.830 563.290 79.830 567.290 ;
        RECT 81.830 565.290 83.830 569.290 ;
        RECT 211.830 567.290 215.830 569.290 ;
        RECT 217.830 571.290 223.830 573.290 ;
        RECT 229.830 571.290 231.830 573.290 ;
        RECT 217.830 569.290 225.830 571.290 ;
        RECT 229.830 569.290 233.830 571.290 ;
        RECT 217.830 567.290 227.830 569.290 ;
        RECT 211.830 565.290 213.830 567.290 ;
        RECT 81.830 563.290 85.830 565.290 ;
        RECT 75.830 559.290 81.830 563.290 ;
        RECT 63.830 557.290 75.830 559.290 ;
        RECT 57.830 555.290 59.830 557.290 ;
        RECT 51.830 553.290 59.830 555.290 ;
        RECT 61.830 553.290 75.830 557.290 ;
        RECT 77.830 557.290 81.830 559.290 ;
        RECT 83.830 559.290 85.830 563.290 ;
        RECT 209.830 563.290 213.830 565.290 ;
        RECT 215.830 563.290 223.830 567.290 ;
        RECT 209.830 559.290 211.830 563.290 ;
        RECT 83.830 557.290 87.830 559.290 ;
        RECT 77.830 555.290 83.830 557.290 ;
        RECT 77.830 553.290 79.830 555.290 ;
        RECT 85.830 553.290 87.830 557.290 ;
        RECT 207.830 557.290 211.830 559.290 ;
        RECT 213.830 559.290 223.830 563.290 ;
        RECT 225.830 563.290 229.830 567.290 ;
        RECT 231.830 565.290 233.830 569.290 ;
        RECT 231.830 563.290 235.830 565.290 ;
        RECT 225.830 559.290 231.830 563.290 ;
        RECT 213.830 557.290 225.830 559.290 ;
        RECT 207.830 555.290 209.830 557.290 ;
        RECT 201.830 553.290 209.830 555.290 ;
        RECT 211.830 553.290 225.830 557.290 ;
        RECT 227.830 557.290 231.830 559.290 ;
        RECT 233.830 559.290 235.830 563.290 ;
        RECT 233.830 557.290 237.830 559.290 ;
        RECT 227.830 555.290 233.830 557.290 ;
        RECT 227.830 553.290 229.830 555.290 ;
        RECT 235.830 553.290 237.830 557.290 ;
        RECT 41.830 551.290 53.830 553.290 ;
        RECT 61.830 551.290 77.830 553.290 ;
        RECT 79.830 551.290 83.830 553.290 ;
        RECT 85.830 551.290 95.830 553.290 ;
        RECT 191.830 551.290 203.830 553.290 ;
        RECT 211.830 551.290 227.830 553.290 ;
        RECT 229.830 551.290 233.830 553.290 ;
        RECT 235.830 551.290 245.830 553.290 ;
        RECT 35.830 549.290 43.830 551.290 ;
        RECT 53.830 549.290 57.830 551.290 ;
        RECT 35.830 545.290 37.830 549.290 ;
        RECT 43.830 547.290 57.830 549.290 ;
        RECT 59.830 547.290 85.830 551.290 ;
        RECT 93.830 549.290 103.830 551.290 ;
        RECT 185.830 549.290 193.830 551.290 ;
        RECT 203.830 549.290 207.830 551.290 ;
        RECT 87.830 547.290 89.830 549.290 ;
        RECT 101.830 547.290 111.830 549.290 ;
        RECT 43.830 545.290 59.830 547.290 ;
        RECT 69.830 545.290 81.830 547.290 ;
        RECT 85.830 545.290 93.830 547.290 ;
        RECT 109.830 545.290 115.830 547.290 ;
        RECT 35.830 543.290 43.830 545.290 ;
        RECT 53.830 543.290 69.830 545.290 ;
        RECT 81.830 543.290 99.830 545.290 ;
        RECT 113.830 543.290 115.830 545.290 ;
        RECT 185.830 545.290 187.830 549.290 ;
        RECT 193.830 547.290 207.830 549.290 ;
        RECT 209.830 547.290 235.830 551.290 ;
        RECT 243.830 549.290 253.830 551.290 ;
        RECT 237.830 547.290 239.830 549.290 ;
        RECT 251.830 547.290 261.830 549.290 ;
        RECT 193.830 545.290 209.830 547.290 ;
        RECT 219.830 545.290 231.830 547.290 ;
        RECT 235.830 545.290 243.830 547.290 ;
        RECT 259.830 545.290 265.830 547.290 ;
        RECT 185.830 543.290 193.830 545.290 ;
        RECT 203.830 543.290 219.830 545.290 ;
        RECT 231.830 543.290 249.830 545.290 ;
        RECT 263.830 543.290 265.830 545.290 ;
        RECT 41.830 541.290 53.830 543.290 ;
        RECT 63.830 541.290 103.830 543.290 ;
        RECT 111.830 541.290 115.830 543.290 ;
        RECT 191.830 541.290 203.830 543.290 ;
        RECT 213.830 541.290 253.830 543.290 ;
        RECT 261.830 541.290 265.830 543.290 ;
        RECT 51.830 539.290 63.830 541.290 ;
        RECT 73.830 539.290 101.830 541.290 ;
        RECT 109.830 539.290 113.830 541.290 ;
        RECT 201.830 539.290 213.830 541.290 ;
        RECT 223.830 539.290 251.830 541.290 ;
        RECT 259.830 539.290 263.830 541.290 ;
        RECT 53.830 537.290 55.830 539.290 ;
        RECT 51.830 535.290 55.830 537.290 ;
        RECT 57.830 537.290 73.830 539.290 ;
        RECT 83.830 537.290 93.830 539.290 ;
        RECT 101.830 537.290 111.830 539.290 ;
        RECT 203.830 537.290 205.830 539.290 ;
        RECT 57.830 535.290 83.830 537.290 ;
        RECT 93.830 535.290 103.830 537.290 ;
        RECT 201.830 535.290 205.830 537.290 ;
        RECT 207.830 537.290 223.830 539.290 ;
        RECT 233.830 537.290 243.830 539.290 ;
        RECT 251.830 537.290 261.830 539.290 ;
        RECT 207.830 535.290 233.830 537.290 ;
        RECT 243.830 535.290 253.830 537.290 ;
        RECT 51.830 529.290 53.830 535.290 ;
        RECT 55.830 533.290 73.830 535.290 ;
        RECT 83.830 533.290 95.830 535.290 ;
        RECT 55.830 531.290 71.830 533.290 ;
        RECT 57.830 529.290 71.830 531.290 ;
        RECT 73.830 531.290 77.830 533.290 ;
        RECT 81.830 531.290 83.830 533.290 ;
        RECT 87.830 531.290 89.830 533.290 ;
        RECT 93.830 531.290 95.830 533.290 ;
        RECT 103.830 531.290 109.830 533.290 ;
        RECT 73.830 529.290 75.830 531.290 ;
        RECT 87.830 529.290 95.830 531.290 ;
        RECT 101.830 529.290 105.830 531.290 ;
        RECT 107.830 529.290 109.830 531.290 ;
        RECT 201.830 529.290 203.830 535.290 ;
        RECT 205.830 533.290 223.830 535.290 ;
        RECT 233.830 533.290 245.830 535.290 ;
        RECT 205.830 531.290 221.830 533.290 ;
        RECT 207.830 529.290 221.830 531.290 ;
        RECT 223.830 531.290 227.830 533.290 ;
        RECT 231.830 531.290 233.830 533.290 ;
        RECT 237.830 531.290 239.830 533.290 ;
        RECT 243.830 531.290 245.830 533.290 ;
        RECT 253.830 531.290 259.830 533.290 ;
        RECT 223.830 529.290 225.830 531.290 ;
        RECT 237.830 529.290 245.830 531.290 ;
        RECT 251.830 529.290 255.830 531.290 ;
        RECT 257.830 529.290 259.830 531.290 ;
        RECT 49.830 527.290 55.830 529.290 ;
        RECT 47.830 525.290 51.830 527.290 ;
        RECT 53.830 525.290 59.830 527.290 ;
        RECT 61.830 525.290 71.830 529.290 ;
        RECT 75.830 527.290 77.830 529.290 ;
        RECT 87.830 527.290 91.830 529.290 ;
        RECT 97.830 527.290 103.830 529.290 ;
        RECT 105.830 527.290 109.830 529.290 ;
        RECT 199.830 527.290 205.830 529.290 ;
        RECT 85.830 525.290 91.830 527.290 ;
        RECT 93.830 525.290 99.830 527.290 ;
        RECT 45.830 523.290 49.830 525.290 ;
        RECT 51.830 523.290 61.830 525.290 ;
        RECT 65.830 523.290 73.830 525.290 ;
        RECT 79.830 523.290 95.830 525.290 ;
        RECT 99.830 523.290 103.830 525.290 ;
        RECT 45.830 517.290 47.830 523.290 ;
        RECT 43.830 515.290 47.830 517.290 ;
        RECT 49.830 521.290 63.830 523.290 ;
        RECT 67.830 521.290 73.830 523.290 ;
        RECT 83.830 521.290 91.830 523.290 ;
        RECT 95.830 521.290 105.830 523.290 ;
        RECT 107.830 521.290 109.830 527.290 ;
        RECT 197.830 525.290 201.830 527.290 ;
        RECT 203.830 525.290 209.830 527.290 ;
        RECT 211.830 525.290 221.830 529.290 ;
        RECT 225.830 527.290 227.830 529.290 ;
        RECT 237.830 527.290 241.830 529.290 ;
        RECT 247.830 527.290 253.830 529.290 ;
        RECT 255.830 527.290 259.830 529.290 ;
        RECT 235.830 525.290 241.830 527.290 ;
        RECT 243.830 525.290 249.830 527.290 ;
        RECT 49.830 519.290 67.830 521.290 ;
        RECT 69.830 519.290 73.830 521.290 ;
        RECT 81.830 519.290 87.830 521.290 ;
        RECT 91.830 519.290 101.830 521.290 ;
        RECT 105.830 519.290 109.830 521.290 ;
        RECT 195.830 523.290 199.830 525.290 ;
        RECT 201.830 523.290 211.830 525.290 ;
        RECT 215.830 523.290 223.830 525.290 ;
        RECT 229.830 523.290 245.830 525.290 ;
        RECT 249.830 523.290 253.830 525.290 ;
        RECT 49.830 517.290 69.830 519.290 ;
        RECT 77.830 517.290 83.830 519.290 ;
        RECT 87.830 517.290 99.830 519.290 ;
        RECT 49.830 515.290 89.830 517.290 ;
        RECT 97.830 515.290 99.830 517.290 ;
        RECT 101.830 517.290 107.830 519.290 ;
        RECT 195.830 517.290 197.830 523.290 ;
        RECT 101.830 515.290 103.830 517.290 ;
        RECT 43.830 495.290 45.830 515.290 ;
        RECT 47.830 513.290 63.830 515.290 ;
        RECT 65.830 513.290 67.830 515.290 ;
        RECT 71.830 513.290 83.830 515.290 ;
        RECT 47.830 511.290 61.830 513.290 ;
        RECT 63.830 511.290 65.830 513.290 ;
        RECT 67.830 511.290 71.830 513.290 ;
        RECT 77.830 511.290 81.830 513.290 ;
        RECT 83.830 511.290 85.830 513.290 ;
        RECT 99.830 511.290 103.830 515.290 ;
        RECT 47.830 509.290 63.830 511.290 ;
        RECT 65.830 509.290 67.830 511.290 ;
        RECT 47.830 507.290 61.830 509.290 ;
        RECT 63.830 507.290 67.830 509.290 ;
        RECT 71.830 509.290 81.830 511.290 ;
        RECT 85.830 509.290 103.830 511.290 ;
        RECT 193.830 515.290 197.830 517.290 ;
        RECT 199.830 521.290 213.830 523.290 ;
        RECT 217.830 521.290 223.830 523.290 ;
        RECT 233.830 521.290 241.830 523.290 ;
        RECT 245.830 521.290 255.830 523.290 ;
        RECT 257.830 521.290 259.830 527.290 ;
        RECT 199.830 519.290 217.830 521.290 ;
        RECT 219.830 519.290 223.830 521.290 ;
        RECT 231.830 519.290 237.830 521.290 ;
        RECT 241.830 519.290 251.830 521.290 ;
        RECT 255.830 519.290 259.830 521.290 ;
        RECT 199.830 517.290 219.830 519.290 ;
        RECT 227.830 517.290 233.830 519.290 ;
        RECT 237.830 517.290 249.830 519.290 ;
        RECT 199.830 515.290 239.830 517.290 ;
        RECT 247.830 515.290 249.830 517.290 ;
        RECT 251.830 517.290 257.830 519.290 ;
        RECT 251.830 515.290 253.830 517.290 ;
        RECT 71.830 507.290 73.830 509.290 ;
        RECT 79.830 507.290 83.830 509.290 ;
        RECT 87.830 507.290 89.830 509.290 ;
        RECT 101.830 507.290 105.830 509.290 ;
        RECT 47.830 505.290 63.830 507.290 ;
        RECT 65.830 505.290 67.830 507.290 ;
        RECT 73.830 505.290 77.830 507.290 ;
        RECT 47.830 503.290 65.830 505.290 ;
        RECT 67.830 503.290 69.830 505.290 ;
        RECT 75.830 503.290 77.830 505.290 ;
        RECT 79.830 505.290 81.830 507.290 ;
        RECT 79.830 503.290 83.830 505.290 ;
        RECT 85.830 503.290 87.830 507.290 ;
        RECT 103.830 505.290 107.830 507.290 ;
        RECT 99.830 503.290 103.830 505.290 ;
        RECT 47.830 501.290 63.830 503.290 ;
        RECT 69.830 501.290 71.830 503.290 ;
        RECT 77.830 501.290 85.830 503.290 ;
        RECT 87.830 501.290 91.830 503.290 ;
        RECT 95.830 501.290 101.830 503.290 ;
        RECT 105.830 501.290 107.830 505.290 ;
        RECT 47.830 499.290 65.830 501.290 ;
        RECT 71.830 499.290 73.830 501.290 ;
        RECT 81.830 499.290 87.830 501.290 ;
        RECT 91.830 499.290 95.830 501.290 ;
        RECT 101.830 499.290 107.830 501.290 ;
        RECT 47.830 497.290 63.830 499.290 ;
        RECT 73.830 497.290 75.830 499.290 ;
        RECT 83.830 497.290 91.830 499.290 ;
        RECT 95.830 497.290 103.830 499.290 ;
        RECT 47.830 495.290 61.830 497.290 ;
        RECT 63.830 495.290 65.830 497.290 ;
        RECT 75.830 495.290 79.830 497.290 ;
        RECT 89.830 495.290 97.830 497.290 ;
        RECT 193.830 495.290 195.830 515.290 ;
        RECT 197.830 513.290 213.830 515.290 ;
        RECT 215.830 513.290 217.830 515.290 ;
        RECT 221.830 513.290 233.830 515.290 ;
        RECT 197.830 511.290 211.830 513.290 ;
        RECT 213.830 511.290 215.830 513.290 ;
        RECT 217.830 511.290 221.830 513.290 ;
        RECT 227.830 511.290 231.830 513.290 ;
        RECT 233.830 511.290 235.830 513.290 ;
        RECT 249.830 511.290 253.830 515.290 ;
        RECT 197.830 509.290 213.830 511.290 ;
        RECT 215.830 509.290 217.830 511.290 ;
        RECT 197.830 507.290 211.830 509.290 ;
        RECT 213.830 507.290 217.830 509.290 ;
        RECT 221.830 509.290 231.830 511.290 ;
        RECT 235.830 509.290 253.830 511.290 ;
        RECT 221.830 507.290 223.830 509.290 ;
        RECT 229.830 507.290 233.830 509.290 ;
        RECT 237.830 507.290 239.830 509.290 ;
        RECT 251.830 507.290 255.830 509.290 ;
        RECT 197.830 505.290 213.830 507.290 ;
        RECT 215.830 505.290 217.830 507.290 ;
        RECT 223.830 505.290 227.830 507.290 ;
        RECT 197.830 503.290 215.830 505.290 ;
        RECT 217.830 503.290 219.830 505.290 ;
        RECT 225.830 503.290 227.830 505.290 ;
        RECT 229.830 505.290 231.830 507.290 ;
        RECT 229.830 503.290 233.830 505.290 ;
        RECT 235.830 503.290 237.830 507.290 ;
        RECT 253.830 505.290 257.830 507.290 ;
        RECT 249.830 503.290 253.830 505.290 ;
        RECT 197.830 501.290 213.830 503.290 ;
        RECT 219.830 501.290 221.830 503.290 ;
        RECT 227.830 501.290 235.830 503.290 ;
        RECT 237.830 501.290 241.830 503.290 ;
        RECT 245.830 501.290 251.830 503.290 ;
        RECT 255.830 501.290 257.830 505.290 ;
        RECT 197.830 499.290 215.830 501.290 ;
        RECT 221.830 499.290 223.830 501.290 ;
        RECT 231.830 499.290 237.830 501.290 ;
        RECT 241.830 499.290 245.830 501.290 ;
        RECT 251.830 499.290 257.830 501.290 ;
        RECT 197.830 497.290 213.830 499.290 ;
        RECT 223.830 497.290 225.830 499.290 ;
        RECT 233.830 497.290 241.830 499.290 ;
        RECT 245.830 497.290 253.830 499.290 ;
        RECT 197.830 495.290 211.830 497.290 ;
        RECT 213.830 495.290 215.830 497.290 ;
        RECT 225.830 495.290 229.830 497.290 ;
        RECT 239.830 495.290 247.830 497.290 ;
        RECT 43.830 493.290 47.830 495.290 ;
        RECT 45.830 477.290 47.830 493.290 ;
        RECT 49.830 491.290 59.830 495.290 ;
        RECT 61.830 493.290 63.830 495.290 ;
        RECT 65.830 493.290 67.830 495.290 ;
        RECT 79.830 493.290 93.830 495.290 ;
        RECT 193.830 493.290 197.830 495.290 ;
        RECT 63.830 491.290 65.830 493.290 ;
        RECT 79.830 491.290 89.830 493.290 ;
        RECT 49.830 489.290 63.830 491.290 ;
        RECT 65.830 489.290 67.830 491.290 ;
        RECT 81.830 489.290 89.830 491.290 ;
        RECT 49.830 487.290 61.830 489.290 ;
        RECT 63.830 487.290 65.830 489.290 ;
        RECT 49.830 485.290 63.830 487.290 ;
        RECT 65.830 485.290 67.830 487.290 ;
        RECT 81.830 485.290 91.830 489.290 ;
        RECT 49.830 483.290 65.830 485.290 ;
        RECT 49.830 481.290 63.830 483.290 ;
        RECT 65.830 481.290 67.830 483.290 ;
        RECT 83.830 481.290 91.830 485.290 ;
        RECT 49.830 479.290 65.830 481.290 ;
        RECT 49.830 477.290 63.830 479.290 ;
        RECT 65.830 477.290 67.830 479.290 ;
        RECT 85.830 477.290 91.830 481.290 ;
        RECT 45.830 475.290 49.830 477.290 ;
        RECT 51.830 475.290 65.830 477.290 ;
        RECT 83.830 475.290 85.830 477.290 ;
        RECT 89.830 475.290 91.830 477.290 ;
        RECT 195.830 477.290 197.830 493.290 ;
        RECT 199.830 491.290 209.830 495.290 ;
        RECT 211.830 493.290 213.830 495.290 ;
        RECT 215.830 493.290 217.830 495.290 ;
        RECT 229.830 493.290 243.830 495.290 ;
        RECT 213.830 491.290 215.830 493.290 ;
        RECT 229.830 491.290 239.830 493.290 ;
        RECT 199.830 489.290 213.830 491.290 ;
        RECT 215.830 489.290 217.830 491.290 ;
        RECT 231.830 489.290 239.830 491.290 ;
        RECT 199.830 487.290 211.830 489.290 ;
        RECT 213.830 487.290 215.830 489.290 ;
        RECT 199.830 485.290 213.830 487.290 ;
        RECT 215.830 485.290 217.830 487.290 ;
        RECT 231.830 485.290 241.830 489.290 ;
        RECT 199.830 483.290 215.830 485.290 ;
        RECT 199.830 481.290 213.830 483.290 ;
        RECT 215.830 481.290 217.830 483.290 ;
        RECT 233.830 481.290 241.830 485.290 ;
        RECT 199.830 479.290 215.830 481.290 ;
        RECT 199.830 477.290 213.830 479.290 ;
        RECT 215.830 477.290 217.830 479.290 ;
        RECT 235.830 477.290 241.830 481.290 ;
        RECT 195.830 475.290 199.830 477.290 ;
        RECT 201.830 475.290 215.830 477.290 ;
        RECT 233.830 475.290 235.830 477.290 ;
        RECT 239.830 475.290 241.830 477.290 ;
        RECT 47.830 473.290 49.830 475.290 ;
        RECT 55.830 473.290 63.830 475.290 ;
        RECT 65.830 473.290 67.830 475.290 ;
        RECT 69.830 473.290 71.830 475.290 ;
        RECT 73.830 473.290 75.830 475.290 ;
        RECT 77.830 473.290 79.830 475.290 ;
        RECT 81.830 473.290 83.830 475.290 ;
        RECT 85.830 473.290 91.830 475.290 ;
        RECT 197.830 473.290 199.830 475.290 ;
        RECT 205.830 473.290 213.830 475.290 ;
        RECT 215.830 473.290 217.830 475.290 ;
        RECT 219.830 473.290 221.830 475.290 ;
        RECT 223.830 473.290 225.830 475.290 ;
        RECT 227.830 473.290 229.830 475.290 ;
        RECT 231.830 473.290 233.830 475.290 ;
        RECT 235.830 473.290 241.830 475.290 ;
        RECT 47.830 471.290 55.830 473.290 ;
        RECT 63.830 471.290 65.830 473.290 ;
        RECT 67.830 471.290 69.830 473.290 ;
        RECT 71.830 471.290 73.830 473.290 ;
        RECT 75.830 471.290 77.830 473.290 ;
        RECT 79.830 471.290 89.830 473.290 ;
        RECT 197.830 471.290 205.830 473.290 ;
        RECT 213.830 471.290 215.830 473.290 ;
        RECT 217.830 471.290 219.830 473.290 ;
        RECT 221.830 471.290 223.830 473.290 ;
        RECT 225.830 471.290 227.830 473.290 ;
        RECT 229.830 471.290 239.830 473.290 ;
        RECT 53.830 469.290 71.830 471.290 ;
        RECT 73.830 469.290 87.830 471.290 ;
        RECT 203.830 469.290 221.830 471.290 ;
        RECT 223.830 469.290 237.830 471.290 ;
        RECT 69.830 467.290 75.830 469.290 ;
        RECT 219.830 467.290 225.830 469.290 ;
        RECT 69.830 439.290 75.830 441.290 ;
        RECT 69.830 437.290 71.830 439.290 ;
        RECT 67.830 435.290 71.830 437.290 ;
        RECT 73.830 437.290 75.830 439.290 ;
        RECT 219.830 439.290 225.830 441.290 ;
        RECT 219.830 437.290 221.830 439.290 ;
        RECT 73.830 435.290 77.830 437.290 ;
        RECT 67.830 431.290 69.830 435.290 ;
        RECT 65.830 429.290 69.830 431.290 ;
        RECT 75.830 431.290 77.830 435.290 ;
        RECT 217.830 435.290 221.830 437.290 ;
        RECT 223.830 437.290 225.830 439.290 ;
        RECT 223.830 435.290 227.830 437.290 ;
        RECT 217.830 431.290 219.830 435.290 ;
        RECT 75.830 429.290 79.830 431.290 ;
        RECT 65.830 425.290 67.830 429.290 ;
        RECT 63.830 423.290 67.830 425.290 ;
        RECT 69.830 423.290 73.830 427.290 ;
        RECT 77.830 425.290 79.830 429.290 ;
        RECT 215.830 429.290 219.830 431.290 ;
        RECT 225.830 431.290 227.830 435.290 ;
        RECT 225.830 429.290 229.830 431.290 ;
        RECT 215.830 425.290 217.830 429.290 ;
        RECT 77.830 423.290 81.830 425.290 ;
        RECT 63.830 419.290 65.830 423.290 ;
        RECT 61.830 417.290 65.830 419.290 ;
        RECT 67.830 421.290 73.830 423.290 ;
        RECT 79.830 421.290 81.830 423.290 ;
        RECT 213.830 423.290 217.830 425.290 ;
        RECT 219.830 423.290 223.830 427.290 ;
        RECT 227.830 425.290 229.830 429.290 ;
        RECT 227.830 423.290 231.830 425.290 ;
        RECT 67.830 419.290 75.830 421.290 ;
        RECT 79.830 419.290 83.830 421.290 ;
        RECT 213.830 419.290 215.830 423.290 ;
        RECT 67.830 417.290 77.830 419.290 ;
        RECT 61.830 415.290 63.830 417.290 ;
        RECT 59.830 413.290 63.830 415.290 ;
        RECT 65.830 413.290 73.830 417.290 ;
        RECT 59.830 409.290 61.830 413.290 ;
        RECT 57.830 407.290 61.830 409.290 ;
        RECT 63.830 409.290 73.830 413.290 ;
        RECT 75.830 413.290 79.830 417.290 ;
        RECT 81.830 415.290 83.830 419.290 ;
        RECT 211.830 417.290 215.830 419.290 ;
        RECT 217.830 421.290 223.830 423.290 ;
        RECT 229.830 421.290 231.830 423.290 ;
        RECT 217.830 419.290 225.830 421.290 ;
        RECT 229.830 419.290 233.830 421.290 ;
        RECT 217.830 417.290 227.830 419.290 ;
        RECT 211.830 415.290 213.830 417.290 ;
        RECT 81.830 413.290 85.830 415.290 ;
        RECT 75.830 409.290 81.830 413.290 ;
        RECT 63.830 407.290 75.830 409.290 ;
        RECT 57.830 405.290 59.830 407.290 ;
        RECT 51.830 403.290 59.830 405.290 ;
        RECT 61.830 403.290 75.830 407.290 ;
        RECT 77.830 407.290 81.830 409.290 ;
        RECT 83.830 409.290 85.830 413.290 ;
        RECT 209.830 413.290 213.830 415.290 ;
        RECT 215.830 413.290 223.830 417.290 ;
        RECT 209.830 409.290 211.830 413.290 ;
        RECT 83.830 407.290 87.830 409.290 ;
        RECT 77.830 405.290 83.830 407.290 ;
        RECT 77.830 403.290 79.830 405.290 ;
        RECT 85.830 403.290 87.830 407.290 ;
        RECT 207.830 407.290 211.830 409.290 ;
        RECT 213.830 409.290 223.830 413.290 ;
        RECT 225.830 413.290 229.830 417.290 ;
        RECT 231.830 415.290 233.830 419.290 ;
        RECT 231.830 413.290 235.830 415.290 ;
        RECT 225.830 409.290 231.830 413.290 ;
        RECT 213.830 407.290 225.830 409.290 ;
        RECT 207.830 405.290 209.830 407.290 ;
        RECT 201.830 403.290 209.830 405.290 ;
        RECT 211.830 403.290 225.830 407.290 ;
        RECT 227.830 407.290 231.830 409.290 ;
        RECT 233.830 409.290 235.830 413.290 ;
        RECT 233.830 407.290 237.830 409.290 ;
        RECT 227.830 405.290 233.830 407.290 ;
        RECT 227.830 403.290 229.830 405.290 ;
        RECT 235.830 403.290 237.830 407.290 ;
        RECT 41.830 401.290 53.830 403.290 ;
        RECT 61.830 401.290 77.830 403.290 ;
        RECT 79.830 401.290 83.830 403.290 ;
        RECT 85.830 401.290 95.830 403.290 ;
        RECT 191.830 401.290 203.830 403.290 ;
        RECT 211.830 401.290 227.830 403.290 ;
        RECT 229.830 401.290 233.830 403.290 ;
        RECT 235.830 401.290 245.830 403.290 ;
        RECT 35.830 399.290 43.830 401.290 ;
        RECT 53.830 399.290 57.830 401.290 ;
        RECT 35.830 395.290 37.830 399.290 ;
        RECT 43.830 397.290 57.830 399.290 ;
        RECT 59.830 397.290 85.830 401.290 ;
        RECT 93.830 399.290 103.830 401.290 ;
        RECT 185.830 399.290 193.830 401.290 ;
        RECT 203.830 399.290 207.830 401.290 ;
        RECT 87.830 397.290 89.830 399.290 ;
        RECT 101.830 397.290 111.830 399.290 ;
        RECT 43.830 395.290 59.830 397.290 ;
        RECT 69.830 395.290 81.830 397.290 ;
        RECT 85.830 395.290 93.830 397.290 ;
        RECT 109.830 395.290 115.830 397.290 ;
        RECT 35.830 393.290 43.830 395.290 ;
        RECT 53.830 393.290 69.830 395.290 ;
        RECT 81.830 393.290 99.830 395.290 ;
        RECT 113.830 393.290 115.830 395.290 ;
        RECT 185.830 395.290 187.830 399.290 ;
        RECT 193.830 397.290 207.830 399.290 ;
        RECT 209.830 397.290 235.830 401.290 ;
        RECT 243.830 399.290 253.830 401.290 ;
        RECT 237.830 397.290 239.830 399.290 ;
        RECT 251.830 397.290 261.830 399.290 ;
        RECT 193.830 395.290 209.830 397.290 ;
        RECT 219.830 395.290 231.830 397.290 ;
        RECT 235.830 395.290 243.830 397.290 ;
        RECT 259.830 395.290 265.830 397.290 ;
        RECT 185.830 393.290 193.830 395.290 ;
        RECT 203.830 393.290 219.830 395.290 ;
        RECT 231.830 393.290 249.830 395.290 ;
        RECT 263.830 393.290 265.830 395.290 ;
        RECT 41.830 391.290 53.830 393.290 ;
        RECT 63.830 391.290 103.830 393.290 ;
        RECT 111.830 391.290 115.830 393.290 ;
        RECT 191.830 391.290 203.830 393.290 ;
        RECT 213.830 391.290 253.830 393.290 ;
        RECT 261.830 391.290 265.830 393.290 ;
        RECT 51.830 389.290 63.830 391.290 ;
        RECT 73.830 389.290 101.830 391.290 ;
        RECT 109.830 389.290 113.830 391.290 ;
        RECT 201.830 389.290 213.830 391.290 ;
        RECT 223.830 389.290 251.830 391.290 ;
        RECT 259.830 389.290 263.830 391.290 ;
        RECT 53.830 387.290 55.830 389.290 ;
        RECT 51.830 385.290 55.830 387.290 ;
        RECT 57.830 387.290 73.830 389.290 ;
        RECT 83.830 387.290 93.830 389.290 ;
        RECT 101.830 387.290 111.830 389.290 ;
        RECT 203.830 387.290 205.830 389.290 ;
        RECT 57.830 385.290 83.830 387.290 ;
        RECT 93.830 385.290 103.830 387.290 ;
        RECT 201.830 385.290 205.830 387.290 ;
        RECT 207.830 387.290 223.830 389.290 ;
        RECT 233.830 387.290 243.830 389.290 ;
        RECT 251.830 387.290 261.830 389.290 ;
        RECT 207.830 385.290 233.830 387.290 ;
        RECT 243.830 385.290 253.830 387.290 ;
        RECT 51.830 379.290 53.830 385.290 ;
        RECT 55.830 383.290 73.830 385.290 ;
        RECT 83.830 383.290 95.830 385.290 ;
        RECT 55.830 381.290 71.830 383.290 ;
        RECT 57.830 379.290 71.830 381.290 ;
        RECT 73.830 381.290 77.830 383.290 ;
        RECT 81.830 381.290 83.830 383.290 ;
        RECT 87.830 381.290 89.830 383.290 ;
        RECT 93.830 381.290 95.830 383.290 ;
        RECT 103.830 381.290 109.830 383.290 ;
        RECT 73.830 379.290 75.830 381.290 ;
        RECT 87.830 379.290 95.830 381.290 ;
        RECT 101.830 379.290 105.830 381.290 ;
        RECT 107.830 379.290 109.830 381.290 ;
        RECT 201.830 379.290 203.830 385.290 ;
        RECT 205.830 383.290 223.830 385.290 ;
        RECT 233.830 383.290 245.830 385.290 ;
        RECT 205.830 381.290 221.830 383.290 ;
        RECT 207.830 379.290 221.830 381.290 ;
        RECT 223.830 381.290 227.830 383.290 ;
        RECT 231.830 381.290 233.830 383.290 ;
        RECT 237.830 381.290 239.830 383.290 ;
        RECT 243.830 381.290 245.830 383.290 ;
        RECT 253.830 381.290 259.830 383.290 ;
        RECT 223.830 379.290 225.830 381.290 ;
        RECT 237.830 379.290 245.830 381.290 ;
        RECT 251.830 379.290 255.830 381.290 ;
        RECT 257.830 379.290 259.830 381.290 ;
        RECT 49.830 377.290 55.830 379.290 ;
        RECT 47.830 375.290 51.830 377.290 ;
        RECT 53.830 375.290 59.830 377.290 ;
        RECT 61.830 375.290 71.830 379.290 ;
        RECT 75.830 377.290 77.830 379.290 ;
        RECT 87.830 377.290 91.830 379.290 ;
        RECT 97.830 377.290 103.830 379.290 ;
        RECT 105.830 377.290 109.830 379.290 ;
        RECT 199.830 377.290 205.830 379.290 ;
        RECT 85.830 375.290 91.830 377.290 ;
        RECT 93.830 375.290 99.830 377.290 ;
        RECT 45.830 373.290 49.830 375.290 ;
        RECT 51.830 373.290 61.830 375.290 ;
        RECT 65.830 373.290 73.830 375.290 ;
        RECT 79.830 373.290 95.830 375.290 ;
        RECT 99.830 373.290 103.830 375.290 ;
        RECT 45.830 367.290 47.830 373.290 ;
        RECT 43.830 365.290 47.830 367.290 ;
        RECT 49.830 371.290 63.830 373.290 ;
        RECT 67.830 371.290 73.830 373.290 ;
        RECT 83.830 371.290 91.830 373.290 ;
        RECT 95.830 371.290 105.830 373.290 ;
        RECT 107.830 371.290 109.830 377.290 ;
        RECT 197.830 375.290 201.830 377.290 ;
        RECT 203.830 375.290 209.830 377.290 ;
        RECT 211.830 375.290 221.830 379.290 ;
        RECT 225.830 377.290 227.830 379.290 ;
        RECT 237.830 377.290 241.830 379.290 ;
        RECT 247.830 377.290 253.830 379.290 ;
        RECT 255.830 377.290 259.830 379.290 ;
        RECT 235.830 375.290 241.830 377.290 ;
        RECT 243.830 375.290 249.830 377.290 ;
        RECT 49.830 369.290 67.830 371.290 ;
        RECT 69.830 369.290 73.830 371.290 ;
        RECT 81.830 369.290 87.830 371.290 ;
        RECT 91.830 369.290 101.830 371.290 ;
        RECT 105.830 369.290 109.830 371.290 ;
        RECT 195.830 373.290 199.830 375.290 ;
        RECT 201.830 373.290 211.830 375.290 ;
        RECT 215.830 373.290 223.830 375.290 ;
        RECT 229.830 373.290 245.830 375.290 ;
        RECT 249.830 373.290 253.830 375.290 ;
        RECT 49.830 367.290 69.830 369.290 ;
        RECT 77.830 367.290 83.830 369.290 ;
        RECT 87.830 367.290 99.830 369.290 ;
        RECT 49.830 365.290 89.830 367.290 ;
        RECT 97.830 365.290 99.830 367.290 ;
        RECT 101.830 367.290 107.830 369.290 ;
        RECT 195.830 367.290 197.830 373.290 ;
        RECT 101.830 365.290 103.830 367.290 ;
        RECT 43.830 345.290 45.830 365.290 ;
        RECT 47.830 363.290 63.830 365.290 ;
        RECT 65.830 363.290 67.830 365.290 ;
        RECT 71.830 363.290 83.830 365.290 ;
        RECT 47.830 361.290 61.830 363.290 ;
        RECT 63.830 361.290 65.830 363.290 ;
        RECT 67.830 361.290 71.830 363.290 ;
        RECT 77.830 361.290 81.830 363.290 ;
        RECT 83.830 361.290 85.830 363.290 ;
        RECT 99.830 361.290 103.830 365.290 ;
        RECT 47.830 359.290 63.830 361.290 ;
        RECT 65.830 359.290 67.830 361.290 ;
        RECT 47.830 357.290 61.830 359.290 ;
        RECT 63.830 357.290 67.830 359.290 ;
        RECT 71.830 359.290 81.830 361.290 ;
        RECT 85.830 359.290 103.830 361.290 ;
        RECT 193.830 365.290 197.830 367.290 ;
        RECT 199.830 371.290 213.830 373.290 ;
        RECT 217.830 371.290 223.830 373.290 ;
        RECT 233.830 371.290 241.830 373.290 ;
        RECT 245.830 371.290 255.830 373.290 ;
        RECT 257.830 371.290 259.830 377.290 ;
        RECT 199.830 369.290 217.830 371.290 ;
        RECT 219.830 369.290 223.830 371.290 ;
        RECT 231.830 369.290 237.830 371.290 ;
        RECT 241.830 369.290 251.830 371.290 ;
        RECT 255.830 369.290 259.830 371.290 ;
        RECT 199.830 367.290 219.830 369.290 ;
        RECT 227.830 367.290 233.830 369.290 ;
        RECT 237.830 367.290 249.830 369.290 ;
        RECT 199.830 365.290 239.830 367.290 ;
        RECT 247.830 365.290 249.830 367.290 ;
        RECT 251.830 367.290 257.830 369.290 ;
        RECT 251.830 365.290 253.830 367.290 ;
        RECT 71.830 357.290 73.830 359.290 ;
        RECT 79.830 357.290 83.830 359.290 ;
        RECT 87.830 357.290 89.830 359.290 ;
        RECT 101.830 357.290 105.830 359.290 ;
        RECT 47.830 355.290 63.830 357.290 ;
        RECT 65.830 355.290 67.830 357.290 ;
        RECT 73.830 355.290 77.830 357.290 ;
        RECT 47.830 353.290 65.830 355.290 ;
        RECT 67.830 353.290 69.830 355.290 ;
        RECT 75.830 353.290 77.830 355.290 ;
        RECT 79.830 355.290 81.830 357.290 ;
        RECT 79.830 353.290 83.830 355.290 ;
        RECT 85.830 353.290 87.830 357.290 ;
        RECT 103.830 355.290 107.830 357.290 ;
        RECT 99.830 353.290 103.830 355.290 ;
        RECT 47.830 351.290 63.830 353.290 ;
        RECT 69.830 351.290 71.830 353.290 ;
        RECT 77.830 351.290 85.830 353.290 ;
        RECT 87.830 351.290 91.830 353.290 ;
        RECT 95.830 351.290 101.830 353.290 ;
        RECT 105.830 351.290 107.830 355.290 ;
        RECT 47.830 349.290 65.830 351.290 ;
        RECT 71.830 349.290 73.830 351.290 ;
        RECT 81.830 349.290 87.830 351.290 ;
        RECT 91.830 349.290 95.830 351.290 ;
        RECT 101.830 349.290 107.830 351.290 ;
        RECT 47.830 347.290 63.830 349.290 ;
        RECT 73.830 347.290 75.830 349.290 ;
        RECT 83.830 347.290 91.830 349.290 ;
        RECT 95.830 347.290 103.830 349.290 ;
        RECT 47.830 345.290 61.830 347.290 ;
        RECT 63.830 345.290 65.830 347.290 ;
        RECT 75.830 345.290 79.830 347.290 ;
        RECT 89.830 345.290 97.830 347.290 ;
        RECT 193.830 345.290 195.830 365.290 ;
        RECT 197.830 363.290 213.830 365.290 ;
        RECT 215.830 363.290 217.830 365.290 ;
        RECT 221.830 363.290 233.830 365.290 ;
        RECT 197.830 361.290 211.830 363.290 ;
        RECT 213.830 361.290 215.830 363.290 ;
        RECT 217.830 361.290 221.830 363.290 ;
        RECT 227.830 361.290 231.830 363.290 ;
        RECT 233.830 361.290 235.830 363.290 ;
        RECT 249.830 361.290 253.830 365.290 ;
        RECT 197.830 359.290 213.830 361.290 ;
        RECT 215.830 359.290 217.830 361.290 ;
        RECT 197.830 357.290 211.830 359.290 ;
        RECT 213.830 357.290 217.830 359.290 ;
        RECT 221.830 359.290 231.830 361.290 ;
        RECT 235.830 359.290 253.830 361.290 ;
        RECT 221.830 357.290 223.830 359.290 ;
        RECT 229.830 357.290 233.830 359.290 ;
        RECT 237.830 357.290 239.830 359.290 ;
        RECT 251.830 357.290 255.830 359.290 ;
        RECT 197.830 355.290 213.830 357.290 ;
        RECT 215.830 355.290 217.830 357.290 ;
        RECT 223.830 355.290 227.830 357.290 ;
        RECT 197.830 353.290 215.830 355.290 ;
        RECT 217.830 353.290 219.830 355.290 ;
        RECT 225.830 353.290 227.830 355.290 ;
        RECT 229.830 355.290 231.830 357.290 ;
        RECT 229.830 353.290 233.830 355.290 ;
        RECT 235.830 353.290 237.830 357.290 ;
        RECT 253.830 355.290 257.830 357.290 ;
        RECT 249.830 353.290 253.830 355.290 ;
        RECT 197.830 351.290 213.830 353.290 ;
        RECT 219.830 351.290 221.830 353.290 ;
        RECT 227.830 351.290 235.830 353.290 ;
        RECT 237.830 351.290 241.830 353.290 ;
        RECT 245.830 351.290 251.830 353.290 ;
        RECT 255.830 351.290 257.830 355.290 ;
        RECT 197.830 349.290 215.830 351.290 ;
        RECT 221.830 349.290 223.830 351.290 ;
        RECT 231.830 349.290 237.830 351.290 ;
        RECT 241.830 349.290 245.830 351.290 ;
        RECT 251.830 349.290 257.830 351.290 ;
        RECT 197.830 347.290 213.830 349.290 ;
        RECT 223.830 347.290 225.830 349.290 ;
        RECT 233.830 347.290 241.830 349.290 ;
        RECT 245.830 347.290 253.830 349.290 ;
        RECT 197.830 345.290 211.830 347.290 ;
        RECT 213.830 345.290 215.830 347.290 ;
        RECT 225.830 345.290 229.830 347.290 ;
        RECT 239.830 345.290 247.830 347.290 ;
        RECT 43.830 343.290 47.830 345.290 ;
        RECT 45.830 327.290 47.830 343.290 ;
        RECT 49.830 341.290 59.830 345.290 ;
        RECT 61.830 343.290 63.830 345.290 ;
        RECT 65.830 343.290 67.830 345.290 ;
        RECT 79.830 343.290 93.830 345.290 ;
        RECT 193.830 343.290 197.830 345.290 ;
        RECT 63.830 341.290 65.830 343.290 ;
        RECT 79.830 341.290 89.830 343.290 ;
        RECT 49.830 339.290 63.830 341.290 ;
        RECT 65.830 339.290 67.830 341.290 ;
        RECT 81.830 339.290 89.830 341.290 ;
        RECT 49.830 337.290 61.830 339.290 ;
        RECT 63.830 337.290 65.830 339.290 ;
        RECT 49.830 335.290 63.830 337.290 ;
        RECT 65.830 335.290 67.830 337.290 ;
        RECT 81.830 335.290 91.830 339.290 ;
        RECT 49.830 333.290 65.830 335.290 ;
        RECT 49.830 331.290 63.830 333.290 ;
        RECT 65.830 331.290 67.830 333.290 ;
        RECT 83.830 331.290 91.830 335.290 ;
        RECT 49.830 329.290 65.830 331.290 ;
        RECT 49.830 327.290 63.830 329.290 ;
        RECT 65.830 327.290 67.830 329.290 ;
        RECT 85.830 327.290 91.830 331.290 ;
        RECT 45.830 325.290 49.830 327.290 ;
        RECT 51.830 325.290 65.830 327.290 ;
        RECT 83.830 325.290 85.830 327.290 ;
        RECT 89.830 325.290 91.830 327.290 ;
        RECT 195.830 327.290 197.830 343.290 ;
        RECT 199.830 341.290 209.830 345.290 ;
        RECT 211.830 343.290 213.830 345.290 ;
        RECT 215.830 343.290 217.830 345.290 ;
        RECT 229.830 343.290 243.830 345.290 ;
        RECT 213.830 341.290 215.830 343.290 ;
        RECT 229.830 341.290 239.830 343.290 ;
        RECT 199.830 339.290 213.830 341.290 ;
        RECT 215.830 339.290 217.830 341.290 ;
        RECT 231.830 339.290 239.830 341.290 ;
        RECT 199.830 337.290 211.830 339.290 ;
        RECT 213.830 337.290 215.830 339.290 ;
        RECT 199.830 335.290 213.830 337.290 ;
        RECT 215.830 335.290 217.830 337.290 ;
        RECT 231.830 335.290 241.830 339.290 ;
        RECT 199.830 333.290 215.830 335.290 ;
        RECT 199.830 331.290 213.830 333.290 ;
        RECT 215.830 331.290 217.830 333.290 ;
        RECT 233.830 331.290 241.830 335.290 ;
        RECT 199.830 329.290 215.830 331.290 ;
        RECT 199.830 327.290 213.830 329.290 ;
        RECT 215.830 327.290 217.830 329.290 ;
        RECT 235.830 327.290 241.830 331.290 ;
        RECT 195.830 325.290 199.830 327.290 ;
        RECT 201.830 325.290 215.830 327.290 ;
        RECT 233.830 325.290 235.830 327.290 ;
        RECT 239.830 325.290 241.830 327.290 ;
        RECT 47.830 323.290 49.830 325.290 ;
        RECT 55.830 323.290 63.830 325.290 ;
        RECT 65.830 323.290 67.830 325.290 ;
        RECT 69.830 323.290 71.830 325.290 ;
        RECT 73.830 323.290 75.830 325.290 ;
        RECT 77.830 323.290 79.830 325.290 ;
        RECT 81.830 323.290 83.830 325.290 ;
        RECT 85.830 323.290 91.830 325.290 ;
        RECT 197.830 323.290 199.830 325.290 ;
        RECT 205.830 323.290 213.830 325.290 ;
        RECT 215.830 323.290 217.830 325.290 ;
        RECT 219.830 323.290 221.830 325.290 ;
        RECT 223.830 323.290 225.830 325.290 ;
        RECT 227.830 323.290 229.830 325.290 ;
        RECT 231.830 323.290 233.830 325.290 ;
        RECT 235.830 323.290 241.830 325.290 ;
        RECT 47.830 321.290 55.830 323.290 ;
        RECT 63.830 321.290 65.830 323.290 ;
        RECT 67.830 321.290 69.830 323.290 ;
        RECT 71.830 321.290 73.830 323.290 ;
        RECT 75.830 321.290 77.830 323.290 ;
        RECT 79.830 321.290 89.830 323.290 ;
        RECT 197.830 321.290 205.830 323.290 ;
        RECT 213.830 321.290 215.830 323.290 ;
        RECT 217.830 321.290 219.830 323.290 ;
        RECT 221.830 321.290 223.830 323.290 ;
        RECT 225.830 321.290 227.830 323.290 ;
        RECT 229.830 321.290 239.830 323.290 ;
        RECT 53.830 319.290 71.830 321.290 ;
        RECT 73.830 319.290 87.830 321.290 ;
        RECT 203.830 319.290 221.830 321.290 ;
        RECT 223.830 319.290 237.830 321.290 ;
        RECT 69.830 317.290 75.830 319.290 ;
        RECT 219.830 317.290 225.830 319.290 ;
        RECT 5.000 60.000 25.000 70.000 ;
        RECT 85.000 30.000 105.000 40.000 ;
        RECT 85.000 5.000 105.000 25.000 ;
        RECT 298.200 0.000 299.800 750.000 ;
  END
END Art
END LIBRARY

