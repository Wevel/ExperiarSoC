magic
tech sky130A
magscale 1 2
timestamp 1653395146
<< obsli1 >>
rect 1104 2159 88872 177361
<< obsm1 >>
rect 14 1300 89962 177744
<< metal2 >>
rect 1122 179200 1178 180000
rect 3422 179200 3478 180000
rect 5722 179200 5778 180000
rect 8022 179200 8078 180000
rect 10322 179200 10378 180000
rect 12622 179200 12678 180000
rect 14922 179200 14978 180000
rect 17222 179200 17278 180000
rect 19522 179200 19578 180000
rect 21822 179200 21878 180000
rect 24122 179200 24178 180000
rect 26422 179200 26478 180000
rect 28722 179200 28778 180000
rect 31114 179200 31170 180000
rect 33414 179200 33470 180000
rect 35714 179200 35770 180000
rect 38014 179200 38070 180000
rect 40314 179200 40370 180000
rect 42614 179200 42670 180000
rect 44914 179200 44970 180000
rect 47214 179200 47270 180000
rect 49514 179200 49570 180000
rect 51814 179200 51870 180000
rect 54114 179200 54170 180000
rect 56414 179200 56470 180000
rect 58714 179200 58770 180000
rect 61106 179200 61162 180000
rect 63406 179200 63462 180000
rect 65706 179200 65762 180000
rect 68006 179200 68062 180000
rect 70306 179200 70362 180000
rect 72606 179200 72662 180000
rect 74906 179200 74962 180000
rect 77206 179200 77262 180000
rect 79506 179200 79562 180000
rect 81806 179200 81862 180000
rect 84106 179200 84162 180000
rect 86406 179200 86462 180000
rect 88706 179200 88762 180000
rect 754 0 810 800
rect 2318 0 2374 800
rect 3974 0 4030 800
rect 5630 0 5686 800
rect 7286 0 7342 800
rect 8850 0 8906 800
rect 10506 0 10562 800
rect 12162 0 12218 800
rect 13818 0 13874 800
rect 15474 0 15530 800
rect 17038 0 17094 800
rect 18694 0 18750 800
rect 20350 0 20406 800
rect 22006 0 22062 800
rect 23570 0 23626 800
rect 25226 0 25282 800
rect 26882 0 26938 800
rect 28538 0 28594 800
rect 30194 0 30250 800
rect 31758 0 31814 800
rect 33414 0 33470 800
rect 35070 0 35126 800
rect 36726 0 36782 800
rect 38290 0 38346 800
rect 39946 0 40002 800
rect 41602 0 41658 800
rect 43258 0 43314 800
rect 44914 0 44970 800
rect 46478 0 46534 800
rect 48134 0 48190 800
rect 49790 0 49846 800
rect 51446 0 51502 800
rect 53102 0 53158 800
rect 54666 0 54722 800
rect 56322 0 56378 800
rect 57978 0 58034 800
rect 59634 0 59690 800
rect 61198 0 61254 800
rect 62854 0 62910 800
rect 64510 0 64566 800
rect 66166 0 66222 800
rect 67822 0 67878 800
rect 69386 0 69442 800
rect 71042 0 71098 800
rect 72698 0 72754 800
rect 74354 0 74410 800
rect 75918 0 75974 800
rect 77574 0 77630 800
rect 79230 0 79286 800
rect 80886 0 80942 800
rect 82542 0 82598 800
rect 84106 0 84162 800
rect 85762 0 85818 800
rect 87418 0 87474 800
rect 89074 0 89130 800
<< obsm2 >>
rect 18 179144 1066 179625
rect 1234 179144 3366 179625
rect 3534 179144 5666 179625
rect 5834 179144 7966 179625
rect 8134 179144 10266 179625
rect 10434 179144 12566 179625
rect 12734 179144 14866 179625
rect 15034 179144 17166 179625
rect 17334 179144 19466 179625
rect 19634 179144 21766 179625
rect 21934 179144 24066 179625
rect 24234 179144 26366 179625
rect 26534 179144 28666 179625
rect 28834 179144 31058 179625
rect 31226 179144 33358 179625
rect 33526 179144 35658 179625
rect 35826 179144 37958 179625
rect 38126 179144 40258 179625
rect 40426 179144 42558 179625
rect 42726 179144 44858 179625
rect 45026 179144 47158 179625
rect 47326 179144 49458 179625
rect 49626 179144 51758 179625
rect 51926 179144 54058 179625
rect 54226 179144 56358 179625
rect 56526 179144 58658 179625
rect 58826 179144 61050 179625
rect 61218 179144 63350 179625
rect 63518 179144 65650 179625
rect 65818 179144 67950 179625
rect 68118 179144 70250 179625
rect 70418 179144 72550 179625
rect 72718 179144 74850 179625
rect 75018 179144 77150 179625
rect 77318 179144 79450 179625
rect 79618 179144 81750 179625
rect 81918 179144 84050 179625
rect 84218 179144 86350 179625
rect 86518 179144 88650 179625
rect 88818 179144 89958 179625
rect 18 856 89958 179144
rect 18 439 698 856
rect 866 439 2262 856
rect 2430 439 3918 856
rect 4086 439 5574 856
rect 5742 439 7230 856
rect 7398 439 8794 856
rect 8962 439 10450 856
rect 10618 439 12106 856
rect 12274 439 13762 856
rect 13930 439 15418 856
rect 15586 439 16982 856
rect 17150 439 18638 856
rect 18806 439 20294 856
rect 20462 439 21950 856
rect 22118 439 23514 856
rect 23682 439 25170 856
rect 25338 439 26826 856
rect 26994 439 28482 856
rect 28650 439 30138 856
rect 30306 439 31702 856
rect 31870 439 33358 856
rect 33526 439 35014 856
rect 35182 439 36670 856
rect 36838 439 38234 856
rect 38402 439 39890 856
rect 40058 439 41546 856
rect 41714 439 43202 856
rect 43370 439 44858 856
rect 45026 439 46422 856
rect 46590 439 48078 856
rect 48246 439 49734 856
rect 49902 439 51390 856
rect 51558 439 53046 856
rect 53214 439 54610 856
rect 54778 439 56266 856
rect 56434 439 57922 856
rect 58090 439 59578 856
rect 59746 439 61142 856
rect 61310 439 62798 856
rect 62966 439 64454 856
rect 64622 439 66110 856
rect 66278 439 67766 856
rect 67934 439 69330 856
rect 69498 439 70986 856
rect 71154 439 72642 856
rect 72810 439 74298 856
rect 74466 439 75862 856
rect 76030 439 77518 856
rect 77686 439 79174 856
rect 79342 439 80830 856
rect 80998 439 82486 856
rect 82654 439 84050 856
rect 84218 439 85706 856
rect 85874 439 87362 856
rect 87530 439 89018 856
rect 89186 439 89958 856
<< metal3 >>
rect 0 179528 800 179648
rect 89200 179528 90000 179648
rect 0 178576 800 178696
rect 89200 178576 90000 178696
rect 0 177624 800 177744
rect 89200 177760 90000 177880
rect 0 176672 800 176792
rect 89200 176808 90000 176928
rect 89200 175992 90000 176112
rect 0 175720 800 175840
rect 89200 175040 90000 175160
rect 0 174768 800 174888
rect 89200 174224 90000 174344
rect 0 173816 800 173936
rect 89200 173272 90000 173392
rect 0 173000 800 173120
rect 89200 172456 90000 172576
rect 0 172048 800 172168
rect 89200 171504 90000 171624
rect 0 171096 800 171216
rect 89200 170552 90000 170672
rect 0 170144 800 170264
rect 89200 169736 90000 169856
rect 0 169192 800 169312
rect 89200 168784 90000 168904
rect 0 168240 800 168360
rect 89200 167968 90000 168088
rect 0 167288 800 167408
rect 89200 167016 90000 167136
rect 0 166472 800 166592
rect 89200 166200 90000 166320
rect 0 165520 800 165640
rect 89200 165248 90000 165368
rect 0 164568 800 164688
rect 89200 164432 90000 164552
rect 0 163616 800 163736
rect 89200 163480 90000 163600
rect 0 162664 800 162784
rect 89200 162528 90000 162648
rect 0 161712 800 161832
rect 89200 161712 90000 161832
rect 0 160760 800 160880
rect 89200 160760 90000 160880
rect 0 159944 800 160064
rect 89200 159944 90000 160064
rect 0 158992 800 159112
rect 89200 158992 90000 159112
rect 0 158040 800 158160
rect 89200 158176 90000 158296
rect 0 157088 800 157208
rect 89200 157224 90000 157344
rect 89200 156408 90000 156528
rect 0 156136 800 156256
rect 89200 155456 90000 155576
rect 0 155184 800 155304
rect 89200 154504 90000 154624
rect 0 154232 800 154352
rect 89200 153688 90000 153808
rect 0 153416 800 153536
rect 89200 152736 90000 152856
rect 0 152464 800 152584
rect 89200 151920 90000 152040
rect 0 151512 800 151632
rect 89200 150968 90000 151088
rect 0 150560 800 150680
rect 89200 150152 90000 150272
rect 0 149608 800 149728
rect 89200 149200 90000 149320
rect 0 148656 800 148776
rect 89200 148384 90000 148504
rect 0 147704 800 147824
rect 89200 147432 90000 147552
rect 0 146888 800 147008
rect 89200 146480 90000 146600
rect 0 145936 800 146056
rect 89200 145664 90000 145784
rect 0 144984 800 145104
rect 89200 144712 90000 144832
rect 0 144032 800 144152
rect 89200 143896 90000 144016
rect 0 143080 800 143200
rect 89200 142944 90000 143064
rect 0 142128 800 142248
rect 89200 142128 90000 142248
rect 0 141176 800 141296
rect 89200 141176 90000 141296
rect 0 140360 800 140480
rect 89200 140360 90000 140480
rect 0 139408 800 139528
rect 89200 139408 90000 139528
rect 0 138456 800 138576
rect 89200 138456 90000 138576
rect 0 137504 800 137624
rect 89200 137640 90000 137760
rect 0 136552 800 136672
rect 89200 136688 90000 136808
rect 89200 135872 90000 135992
rect 0 135600 800 135720
rect 89200 134920 90000 135040
rect 0 134648 800 134768
rect 89200 134104 90000 134224
rect 0 133696 800 133816
rect 89200 133152 90000 133272
rect 0 132880 800 133000
rect 89200 132336 90000 132456
rect 0 131928 800 132048
rect 89200 131384 90000 131504
rect 0 130976 800 131096
rect 89200 130432 90000 130552
rect 0 130024 800 130144
rect 89200 129616 90000 129736
rect 0 129072 800 129192
rect 89200 128664 90000 128784
rect 0 128120 800 128240
rect 89200 127848 90000 127968
rect 0 127168 800 127288
rect 89200 126896 90000 127016
rect 0 126352 800 126472
rect 89200 126080 90000 126200
rect 0 125400 800 125520
rect 89200 125128 90000 125248
rect 0 124448 800 124568
rect 89200 124312 90000 124432
rect 0 123496 800 123616
rect 89200 123360 90000 123480
rect 0 122544 800 122664
rect 89200 122408 90000 122528
rect 0 121592 800 121712
rect 89200 121592 90000 121712
rect 0 120640 800 120760
rect 89200 120640 90000 120760
rect 0 119824 800 119944
rect 89200 119824 90000 119944
rect 0 118872 800 118992
rect 89200 118872 90000 118992
rect 0 117920 800 118040
rect 89200 118056 90000 118176
rect 0 116968 800 117088
rect 89200 117104 90000 117224
rect 89200 116288 90000 116408
rect 0 116016 800 116136
rect 89200 115336 90000 115456
rect 0 115064 800 115184
rect 89200 114384 90000 114504
rect 0 114112 800 114232
rect 89200 113568 90000 113688
rect 0 113296 800 113416
rect 89200 112616 90000 112736
rect 0 112344 800 112464
rect 89200 111800 90000 111920
rect 0 111392 800 111512
rect 89200 110848 90000 110968
rect 0 110440 800 110560
rect 89200 110032 90000 110152
rect 0 109488 800 109608
rect 89200 109080 90000 109200
rect 0 108536 800 108656
rect 89200 108264 90000 108384
rect 0 107584 800 107704
rect 89200 107312 90000 107432
rect 0 106768 800 106888
rect 89200 106360 90000 106480
rect 0 105816 800 105936
rect 89200 105544 90000 105664
rect 0 104864 800 104984
rect 89200 104592 90000 104712
rect 0 103912 800 104032
rect 89200 103776 90000 103896
rect 0 102960 800 103080
rect 89200 102824 90000 102944
rect 0 102008 800 102128
rect 89200 102008 90000 102128
rect 0 101056 800 101176
rect 89200 101056 90000 101176
rect 0 100240 800 100360
rect 89200 100240 90000 100360
rect 0 99288 800 99408
rect 89200 99288 90000 99408
rect 0 98336 800 98456
rect 89200 98336 90000 98456
rect 0 97384 800 97504
rect 89200 97520 90000 97640
rect 0 96432 800 96552
rect 89200 96568 90000 96688
rect 89200 95752 90000 95872
rect 0 95480 800 95600
rect 89200 94800 90000 94920
rect 0 94528 800 94648
rect 89200 93984 90000 94104
rect 0 93712 800 93832
rect 89200 93032 90000 93152
rect 0 92760 800 92880
rect 89200 92216 90000 92336
rect 0 91808 800 91928
rect 89200 91264 90000 91384
rect 0 90856 800 90976
rect 89200 90448 90000 90568
rect 0 89904 800 90024
rect 89200 89496 90000 89616
rect 0 88952 800 89072
rect 89200 88544 90000 88664
rect 0 88000 800 88120
rect 89200 87728 90000 87848
rect 0 87048 800 87168
rect 89200 86776 90000 86896
rect 0 86232 800 86352
rect 89200 85960 90000 86080
rect 0 85280 800 85400
rect 89200 85008 90000 85128
rect 0 84328 800 84448
rect 89200 84192 90000 84312
rect 0 83376 800 83496
rect 89200 83240 90000 83360
rect 0 82424 800 82544
rect 89200 82424 90000 82544
rect 0 81472 800 81592
rect 89200 81472 90000 81592
rect 0 80520 800 80640
rect 89200 80520 90000 80640
rect 0 79704 800 79824
rect 89200 79704 90000 79824
rect 0 78752 800 78872
rect 89200 78752 90000 78872
rect 0 77800 800 77920
rect 89200 77936 90000 78056
rect 0 76848 800 76968
rect 89200 76984 90000 77104
rect 89200 76168 90000 76288
rect 0 75896 800 76016
rect 89200 75216 90000 75336
rect 0 74944 800 75064
rect 89200 74400 90000 74520
rect 0 73992 800 74112
rect 89200 73448 90000 73568
rect 0 73176 800 73296
rect 89200 72496 90000 72616
rect 0 72224 800 72344
rect 89200 71680 90000 71800
rect 0 71272 800 71392
rect 89200 70728 90000 70848
rect 0 70320 800 70440
rect 89200 69912 90000 70032
rect 0 69368 800 69488
rect 89200 68960 90000 69080
rect 0 68416 800 68536
rect 89200 68144 90000 68264
rect 0 67464 800 67584
rect 89200 67192 90000 67312
rect 0 66648 800 66768
rect 89200 66376 90000 66496
rect 0 65696 800 65816
rect 89200 65424 90000 65544
rect 0 64744 800 64864
rect 89200 64472 90000 64592
rect 0 63792 800 63912
rect 89200 63656 90000 63776
rect 0 62840 800 62960
rect 89200 62704 90000 62824
rect 0 61888 800 62008
rect 89200 61888 90000 62008
rect 0 60936 800 61056
rect 89200 60936 90000 61056
rect 0 60120 800 60240
rect 89200 60120 90000 60240
rect 0 59168 800 59288
rect 89200 59168 90000 59288
rect 0 58216 800 58336
rect 89200 58352 90000 58472
rect 0 57264 800 57384
rect 89200 57400 90000 57520
rect 0 56312 800 56432
rect 89200 56448 90000 56568
rect 89200 55632 90000 55752
rect 0 55360 800 55480
rect 89200 54680 90000 54800
rect 0 54408 800 54528
rect 89200 53864 90000 53984
rect 0 53592 800 53712
rect 89200 52912 90000 53032
rect 0 52640 800 52760
rect 89200 52096 90000 52216
rect 0 51688 800 51808
rect 89200 51144 90000 51264
rect 0 50736 800 50856
rect 89200 50328 90000 50448
rect 0 49784 800 49904
rect 89200 49376 90000 49496
rect 0 48832 800 48952
rect 89200 48424 90000 48544
rect 0 47880 800 48000
rect 89200 47608 90000 47728
rect 0 47064 800 47184
rect 89200 46656 90000 46776
rect 0 46112 800 46232
rect 89200 45840 90000 45960
rect 0 45160 800 45280
rect 89200 44888 90000 45008
rect 0 44208 800 44328
rect 89200 44072 90000 44192
rect 0 43256 800 43376
rect 89200 43120 90000 43240
rect 0 42304 800 42424
rect 89200 42304 90000 42424
rect 0 41352 800 41472
rect 89200 41352 90000 41472
rect 0 40400 800 40520
rect 89200 40400 90000 40520
rect 0 39584 800 39704
rect 89200 39584 90000 39704
rect 0 38632 800 38752
rect 89200 38632 90000 38752
rect 0 37680 800 37800
rect 89200 37816 90000 37936
rect 0 36728 800 36848
rect 89200 36864 90000 36984
rect 89200 36048 90000 36168
rect 0 35776 800 35896
rect 89200 35096 90000 35216
rect 0 34824 800 34944
rect 89200 34280 90000 34400
rect 0 33872 800 33992
rect 89200 33328 90000 33448
rect 0 33056 800 33176
rect 89200 32376 90000 32496
rect 0 32104 800 32224
rect 89200 31560 90000 31680
rect 0 31152 800 31272
rect 89200 30608 90000 30728
rect 0 30200 800 30320
rect 89200 29792 90000 29912
rect 0 29248 800 29368
rect 89200 28840 90000 28960
rect 0 28296 800 28416
rect 89200 28024 90000 28144
rect 0 27344 800 27464
rect 89200 27072 90000 27192
rect 0 26528 800 26648
rect 89200 26256 90000 26376
rect 0 25576 800 25696
rect 89200 25304 90000 25424
rect 0 24624 800 24744
rect 89200 24352 90000 24472
rect 0 23672 800 23792
rect 89200 23536 90000 23656
rect 0 22720 800 22840
rect 89200 22584 90000 22704
rect 0 21768 800 21888
rect 89200 21768 90000 21888
rect 0 20816 800 20936
rect 89200 20816 90000 20936
rect 0 20000 800 20120
rect 89200 20000 90000 20120
rect 0 19048 800 19168
rect 89200 19048 90000 19168
rect 0 18096 800 18216
rect 89200 18232 90000 18352
rect 0 17144 800 17264
rect 89200 17280 90000 17400
rect 0 16192 800 16312
rect 89200 16328 90000 16448
rect 89200 15512 90000 15632
rect 0 15240 800 15360
rect 89200 14560 90000 14680
rect 0 14288 800 14408
rect 89200 13744 90000 13864
rect 0 13472 800 13592
rect 89200 12792 90000 12912
rect 0 12520 800 12640
rect 89200 11976 90000 12096
rect 0 11568 800 11688
rect 89200 11024 90000 11144
rect 0 10616 800 10736
rect 89200 10208 90000 10328
rect 0 9664 800 9784
rect 89200 9256 90000 9376
rect 0 8712 800 8832
rect 89200 8304 90000 8424
rect 0 7760 800 7880
rect 89200 7488 90000 7608
rect 0 6944 800 7064
rect 89200 6536 90000 6656
rect 0 5992 800 6112
rect 89200 5720 90000 5840
rect 0 5040 800 5160
rect 89200 4768 90000 4888
rect 0 4088 800 4208
rect 89200 3952 90000 4072
rect 0 3136 800 3256
rect 89200 3000 90000 3120
rect 0 2184 800 2304
rect 89200 2184 90000 2304
rect 0 1232 800 1352
rect 89200 1232 90000 1352
rect 0 416 800 536
rect 89200 416 90000 536
<< obsm3 >>
rect 880 179448 89120 179621
rect 13 178776 89963 179448
rect 880 178496 89120 178776
rect 13 177960 89963 178496
rect 13 177824 89120 177960
rect 880 177680 89120 177824
rect 880 177544 89963 177680
rect 13 177008 89963 177544
rect 13 176872 89120 177008
rect 880 176728 89120 176872
rect 880 176592 89963 176728
rect 13 176192 89963 176592
rect 13 175920 89120 176192
rect 880 175912 89120 175920
rect 880 175640 89963 175912
rect 13 175240 89963 175640
rect 13 174968 89120 175240
rect 880 174960 89120 174968
rect 880 174688 89963 174960
rect 13 174424 89963 174688
rect 13 174144 89120 174424
rect 13 174016 89963 174144
rect 880 173736 89963 174016
rect 13 173472 89963 173736
rect 13 173200 89120 173472
rect 880 173192 89120 173200
rect 880 172920 89963 173192
rect 13 172656 89963 172920
rect 13 172376 89120 172656
rect 13 172248 89963 172376
rect 880 171968 89963 172248
rect 13 171704 89963 171968
rect 13 171424 89120 171704
rect 13 171296 89963 171424
rect 880 171016 89963 171296
rect 13 170752 89963 171016
rect 13 170472 89120 170752
rect 13 170344 89963 170472
rect 880 170064 89963 170344
rect 13 169936 89963 170064
rect 13 169656 89120 169936
rect 13 169392 89963 169656
rect 880 169112 89963 169392
rect 13 168984 89963 169112
rect 13 168704 89120 168984
rect 13 168440 89963 168704
rect 880 168168 89963 168440
rect 880 168160 89120 168168
rect 13 167888 89120 168160
rect 13 167488 89963 167888
rect 880 167216 89963 167488
rect 880 167208 89120 167216
rect 13 166936 89120 167208
rect 13 166672 89963 166936
rect 880 166400 89963 166672
rect 880 166392 89120 166400
rect 13 166120 89120 166392
rect 13 165720 89963 166120
rect 880 165448 89963 165720
rect 880 165440 89120 165448
rect 13 165168 89120 165440
rect 13 164768 89963 165168
rect 880 164632 89963 164768
rect 880 164488 89120 164632
rect 13 164352 89120 164488
rect 13 163816 89963 164352
rect 880 163680 89963 163816
rect 880 163536 89120 163680
rect 13 163400 89120 163536
rect 13 162864 89963 163400
rect 880 162728 89963 162864
rect 880 162584 89120 162728
rect 13 162448 89120 162584
rect 13 161912 89963 162448
rect 880 161632 89120 161912
rect 13 160960 89963 161632
rect 880 160680 89120 160960
rect 13 160144 89963 160680
rect 880 159864 89120 160144
rect 13 159192 89963 159864
rect 880 158912 89120 159192
rect 13 158376 89963 158912
rect 13 158240 89120 158376
rect 880 158096 89120 158240
rect 880 157960 89963 158096
rect 13 157424 89963 157960
rect 13 157288 89120 157424
rect 880 157144 89120 157288
rect 880 157008 89963 157144
rect 13 156608 89963 157008
rect 13 156336 89120 156608
rect 880 156328 89120 156336
rect 880 156056 89963 156328
rect 13 155656 89963 156056
rect 13 155384 89120 155656
rect 880 155376 89120 155384
rect 880 155104 89963 155376
rect 13 154704 89963 155104
rect 13 154432 89120 154704
rect 880 154424 89120 154432
rect 880 154152 89963 154424
rect 13 153888 89963 154152
rect 13 153616 89120 153888
rect 880 153608 89120 153616
rect 880 153336 89963 153608
rect 13 152936 89963 153336
rect 13 152664 89120 152936
rect 880 152656 89120 152664
rect 880 152384 89963 152656
rect 13 152120 89963 152384
rect 13 151840 89120 152120
rect 13 151712 89963 151840
rect 880 151432 89963 151712
rect 13 151168 89963 151432
rect 13 150888 89120 151168
rect 13 150760 89963 150888
rect 880 150480 89963 150760
rect 13 150352 89963 150480
rect 13 150072 89120 150352
rect 13 149808 89963 150072
rect 880 149528 89963 149808
rect 13 149400 89963 149528
rect 13 149120 89120 149400
rect 13 148856 89963 149120
rect 880 148584 89963 148856
rect 880 148576 89120 148584
rect 13 148304 89120 148576
rect 13 147904 89963 148304
rect 880 147632 89963 147904
rect 880 147624 89120 147632
rect 13 147352 89120 147624
rect 13 147088 89963 147352
rect 880 146808 89963 147088
rect 13 146680 89963 146808
rect 13 146400 89120 146680
rect 13 146136 89963 146400
rect 880 145864 89963 146136
rect 880 145856 89120 145864
rect 13 145584 89120 145856
rect 13 145184 89963 145584
rect 880 144912 89963 145184
rect 880 144904 89120 144912
rect 13 144632 89120 144904
rect 13 144232 89963 144632
rect 880 144096 89963 144232
rect 880 143952 89120 144096
rect 13 143816 89120 143952
rect 13 143280 89963 143816
rect 880 143144 89963 143280
rect 880 143000 89120 143144
rect 13 142864 89120 143000
rect 13 142328 89963 142864
rect 880 142048 89120 142328
rect 13 141376 89963 142048
rect 880 141096 89120 141376
rect 13 140560 89963 141096
rect 880 140280 89120 140560
rect 13 139608 89963 140280
rect 880 139328 89120 139608
rect 13 138656 89963 139328
rect 880 138376 89120 138656
rect 13 137840 89963 138376
rect 13 137704 89120 137840
rect 880 137560 89120 137704
rect 880 137424 89963 137560
rect 13 136888 89963 137424
rect 13 136752 89120 136888
rect 880 136608 89120 136752
rect 880 136472 89963 136608
rect 13 136072 89963 136472
rect 13 135800 89120 136072
rect 880 135792 89120 135800
rect 880 135520 89963 135792
rect 13 135120 89963 135520
rect 13 134848 89120 135120
rect 880 134840 89120 134848
rect 880 134568 89963 134840
rect 13 134304 89963 134568
rect 13 134024 89120 134304
rect 13 133896 89963 134024
rect 880 133616 89963 133896
rect 13 133352 89963 133616
rect 13 133080 89120 133352
rect 880 133072 89120 133080
rect 880 132800 89963 133072
rect 13 132536 89963 132800
rect 13 132256 89120 132536
rect 13 132128 89963 132256
rect 880 131848 89963 132128
rect 13 131584 89963 131848
rect 13 131304 89120 131584
rect 13 131176 89963 131304
rect 880 130896 89963 131176
rect 13 130632 89963 130896
rect 13 130352 89120 130632
rect 13 130224 89963 130352
rect 880 129944 89963 130224
rect 13 129816 89963 129944
rect 13 129536 89120 129816
rect 13 129272 89963 129536
rect 880 128992 89963 129272
rect 13 128864 89963 128992
rect 13 128584 89120 128864
rect 13 128320 89963 128584
rect 880 128048 89963 128320
rect 880 128040 89120 128048
rect 13 127768 89120 128040
rect 13 127368 89963 127768
rect 880 127096 89963 127368
rect 880 127088 89120 127096
rect 13 126816 89120 127088
rect 13 126552 89963 126816
rect 880 126280 89963 126552
rect 880 126272 89120 126280
rect 13 126000 89120 126272
rect 13 125600 89963 126000
rect 880 125328 89963 125600
rect 880 125320 89120 125328
rect 13 125048 89120 125320
rect 13 124648 89963 125048
rect 880 124512 89963 124648
rect 880 124368 89120 124512
rect 13 124232 89120 124368
rect 13 123696 89963 124232
rect 880 123560 89963 123696
rect 880 123416 89120 123560
rect 13 123280 89120 123416
rect 13 122744 89963 123280
rect 880 122608 89963 122744
rect 880 122464 89120 122608
rect 13 122328 89120 122464
rect 13 121792 89963 122328
rect 880 121512 89120 121792
rect 13 120840 89963 121512
rect 880 120560 89120 120840
rect 13 120024 89963 120560
rect 880 119744 89120 120024
rect 13 119072 89963 119744
rect 880 118792 89120 119072
rect 13 118256 89963 118792
rect 13 118120 89120 118256
rect 880 117976 89120 118120
rect 880 117840 89963 117976
rect 13 117304 89963 117840
rect 13 117168 89120 117304
rect 880 117024 89120 117168
rect 880 116888 89963 117024
rect 13 116488 89963 116888
rect 13 116216 89120 116488
rect 880 116208 89120 116216
rect 880 115936 89963 116208
rect 13 115536 89963 115936
rect 13 115264 89120 115536
rect 880 115256 89120 115264
rect 880 114984 89963 115256
rect 13 114584 89963 114984
rect 13 114312 89120 114584
rect 880 114304 89120 114312
rect 880 114032 89963 114304
rect 13 113768 89963 114032
rect 13 113496 89120 113768
rect 880 113488 89120 113496
rect 880 113216 89963 113488
rect 13 112816 89963 113216
rect 13 112544 89120 112816
rect 880 112536 89120 112544
rect 880 112264 89963 112536
rect 13 112000 89963 112264
rect 13 111720 89120 112000
rect 13 111592 89963 111720
rect 880 111312 89963 111592
rect 13 111048 89963 111312
rect 13 110768 89120 111048
rect 13 110640 89963 110768
rect 880 110360 89963 110640
rect 13 110232 89963 110360
rect 13 109952 89120 110232
rect 13 109688 89963 109952
rect 880 109408 89963 109688
rect 13 109280 89963 109408
rect 13 109000 89120 109280
rect 13 108736 89963 109000
rect 880 108464 89963 108736
rect 880 108456 89120 108464
rect 13 108184 89120 108456
rect 13 107784 89963 108184
rect 880 107512 89963 107784
rect 880 107504 89120 107512
rect 13 107232 89120 107504
rect 13 106968 89963 107232
rect 880 106688 89963 106968
rect 13 106560 89963 106688
rect 13 106280 89120 106560
rect 13 106016 89963 106280
rect 880 105744 89963 106016
rect 880 105736 89120 105744
rect 13 105464 89120 105736
rect 13 105064 89963 105464
rect 880 104792 89963 105064
rect 880 104784 89120 104792
rect 13 104512 89120 104784
rect 13 104112 89963 104512
rect 880 103976 89963 104112
rect 880 103832 89120 103976
rect 13 103696 89120 103832
rect 13 103160 89963 103696
rect 880 103024 89963 103160
rect 880 102880 89120 103024
rect 13 102744 89120 102880
rect 13 102208 89963 102744
rect 880 101928 89120 102208
rect 13 101256 89963 101928
rect 880 100976 89120 101256
rect 13 100440 89963 100976
rect 880 100160 89120 100440
rect 13 99488 89963 100160
rect 880 99208 89120 99488
rect 13 98536 89963 99208
rect 880 98256 89120 98536
rect 13 97720 89963 98256
rect 13 97584 89120 97720
rect 880 97440 89120 97584
rect 880 97304 89963 97440
rect 13 96768 89963 97304
rect 13 96632 89120 96768
rect 880 96488 89120 96632
rect 880 96352 89963 96488
rect 13 95952 89963 96352
rect 13 95680 89120 95952
rect 880 95672 89120 95680
rect 880 95400 89963 95672
rect 13 95000 89963 95400
rect 13 94728 89120 95000
rect 880 94720 89120 94728
rect 880 94448 89963 94720
rect 13 94184 89963 94448
rect 13 93912 89120 94184
rect 880 93904 89120 93912
rect 880 93632 89963 93904
rect 13 93232 89963 93632
rect 13 92960 89120 93232
rect 880 92952 89120 92960
rect 880 92680 89963 92952
rect 13 92416 89963 92680
rect 13 92136 89120 92416
rect 13 92008 89963 92136
rect 880 91728 89963 92008
rect 13 91464 89963 91728
rect 13 91184 89120 91464
rect 13 91056 89963 91184
rect 880 90776 89963 91056
rect 13 90648 89963 90776
rect 13 90368 89120 90648
rect 13 90104 89963 90368
rect 880 89824 89963 90104
rect 13 89696 89963 89824
rect 13 89416 89120 89696
rect 13 89152 89963 89416
rect 880 88872 89963 89152
rect 13 88744 89963 88872
rect 13 88464 89120 88744
rect 13 88200 89963 88464
rect 880 87928 89963 88200
rect 880 87920 89120 87928
rect 13 87648 89120 87920
rect 13 87248 89963 87648
rect 880 86976 89963 87248
rect 880 86968 89120 86976
rect 13 86696 89120 86968
rect 13 86432 89963 86696
rect 880 86160 89963 86432
rect 880 86152 89120 86160
rect 13 85880 89120 86152
rect 13 85480 89963 85880
rect 880 85208 89963 85480
rect 880 85200 89120 85208
rect 13 84928 89120 85200
rect 13 84528 89963 84928
rect 880 84392 89963 84528
rect 880 84248 89120 84392
rect 13 84112 89120 84248
rect 13 83576 89963 84112
rect 880 83440 89963 83576
rect 880 83296 89120 83440
rect 13 83160 89120 83296
rect 13 82624 89963 83160
rect 880 82344 89120 82624
rect 13 81672 89963 82344
rect 880 81392 89120 81672
rect 13 80720 89963 81392
rect 880 80440 89120 80720
rect 13 79904 89963 80440
rect 880 79624 89120 79904
rect 13 78952 89963 79624
rect 880 78672 89120 78952
rect 13 78136 89963 78672
rect 13 78000 89120 78136
rect 880 77856 89120 78000
rect 880 77720 89963 77856
rect 13 77184 89963 77720
rect 13 77048 89120 77184
rect 880 76904 89120 77048
rect 880 76768 89963 76904
rect 13 76368 89963 76768
rect 13 76096 89120 76368
rect 880 76088 89120 76096
rect 880 75816 89963 76088
rect 13 75416 89963 75816
rect 13 75144 89120 75416
rect 880 75136 89120 75144
rect 880 74864 89963 75136
rect 13 74600 89963 74864
rect 13 74320 89120 74600
rect 13 74192 89963 74320
rect 880 73912 89963 74192
rect 13 73648 89963 73912
rect 13 73376 89120 73648
rect 880 73368 89120 73376
rect 880 73096 89963 73368
rect 13 72696 89963 73096
rect 13 72424 89120 72696
rect 880 72416 89120 72424
rect 880 72144 89963 72416
rect 13 71880 89963 72144
rect 13 71600 89120 71880
rect 13 71472 89963 71600
rect 880 71192 89963 71472
rect 13 70928 89963 71192
rect 13 70648 89120 70928
rect 13 70520 89963 70648
rect 880 70240 89963 70520
rect 13 70112 89963 70240
rect 13 69832 89120 70112
rect 13 69568 89963 69832
rect 880 69288 89963 69568
rect 13 69160 89963 69288
rect 13 68880 89120 69160
rect 13 68616 89963 68880
rect 880 68344 89963 68616
rect 880 68336 89120 68344
rect 13 68064 89120 68336
rect 13 67664 89963 68064
rect 880 67392 89963 67664
rect 880 67384 89120 67392
rect 13 67112 89120 67384
rect 13 66848 89963 67112
rect 880 66576 89963 66848
rect 880 66568 89120 66576
rect 13 66296 89120 66568
rect 13 65896 89963 66296
rect 880 65624 89963 65896
rect 880 65616 89120 65624
rect 13 65344 89120 65616
rect 13 64944 89963 65344
rect 880 64672 89963 64944
rect 880 64664 89120 64672
rect 13 64392 89120 64664
rect 13 63992 89963 64392
rect 880 63856 89963 63992
rect 880 63712 89120 63856
rect 13 63576 89120 63712
rect 13 63040 89963 63576
rect 880 62904 89963 63040
rect 880 62760 89120 62904
rect 13 62624 89120 62760
rect 13 62088 89963 62624
rect 880 61808 89120 62088
rect 13 61136 89963 61808
rect 880 60856 89120 61136
rect 13 60320 89963 60856
rect 880 60040 89120 60320
rect 13 59368 89963 60040
rect 880 59088 89120 59368
rect 13 58552 89963 59088
rect 13 58416 89120 58552
rect 880 58272 89120 58416
rect 880 58136 89963 58272
rect 13 57600 89963 58136
rect 13 57464 89120 57600
rect 880 57320 89120 57464
rect 880 57184 89963 57320
rect 13 56648 89963 57184
rect 13 56512 89120 56648
rect 880 56368 89120 56512
rect 880 56232 89963 56368
rect 13 55832 89963 56232
rect 13 55560 89120 55832
rect 880 55552 89120 55560
rect 880 55280 89963 55552
rect 13 54880 89963 55280
rect 13 54608 89120 54880
rect 880 54600 89120 54608
rect 880 54328 89963 54600
rect 13 54064 89963 54328
rect 13 53792 89120 54064
rect 880 53784 89120 53792
rect 880 53512 89963 53784
rect 13 53112 89963 53512
rect 13 52840 89120 53112
rect 880 52832 89120 52840
rect 880 52560 89963 52832
rect 13 52296 89963 52560
rect 13 52016 89120 52296
rect 13 51888 89963 52016
rect 880 51608 89963 51888
rect 13 51344 89963 51608
rect 13 51064 89120 51344
rect 13 50936 89963 51064
rect 880 50656 89963 50936
rect 13 50528 89963 50656
rect 13 50248 89120 50528
rect 13 49984 89963 50248
rect 880 49704 89963 49984
rect 13 49576 89963 49704
rect 13 49296 89120 49576
rect 13 49032 89963 49296
rect 880 48752 89963 49032
rect 13 48624 89963 48752
rect 13 48344 89120 48624
rect 13 48080 89963 48344
rect 880 47808 89963 48080
rect 880 47800 89120 47808
rect 13 47528 89120 47800
rect 13 47264 89963 47528
rect 880 46984 89963 47264
rect 13 46856 89963 46984
rect 13 46576 89120 46856
rect 13 46312 89963 46576
rect 880 46040 89963 46312
rect 880 46032 89120 46040
rect 13 45760 89120 46032
rect 13 45360 89963 45760
rect 880 45088 89963 45360
rect 880 45080 89120 45088
rect 13 44808 89120 45080
rect 13 44408 89963 44808
rect 880 44272 89963 44408
rect 880 44128 89120 44272
rect 13 43992 89120 44128
rect 13 43456 89963 43992
rect 880 43320 89963 43456
rect 880 43176 89120 43320
rect 13 43040 89120 43176
rect 13 42504 89963 43040
rect 880 42224 89120 42504
rect 13 41552 89963 42224
rect 880 41272 89120 41552
rect 13 40600 89963 41272
rect 880 40320 89120 40600
rect 13 39784 89963 40320
rect 880 39504 89120 39784
rect 13 38832 89963 39504
rect 880 38552 89120 38832
rect 13 38016 89963 38552
rect 13 37880 89120 38016
rect 880 37736 89120 37880
rect 880 37600 89963 37736
rect 13 37064 89963 37600
rect 13 36928 89120 37064
rect 880 36784 89120 36928
rect 880 36648 89963 36784
rect 13 36248 89963 36648
rect 13 35976 89120 36248
rect 880 35968 89120 35976
rect 880 35696 89963 35968
rect 13 35296 89963 35696
rect 13 35024 89120 35296
rect 880 35016 89120 35024
rect 880 34744 89963 35016
rect 13 34480 89963 34744
rect 13 34200 89120 34480
rect 13 34072 89963 34200
rect 880 33792 89963 34072
rect 13 33528 89963 33792
rect 13 33256 89120 33528
rect 880 33248 89120 33256
rect 880 32976 89963 33248
rect 13 32576 89963 32976
rect 13 32304 89120 32576
rect 880 32296 89120 32304
rect 880 32024 89963 32296
rect 13 31760 89963 32024
rect 13 31480 89120 31760
rect 13 31352 89963 31480
rect 880 31072 89963 31352
rect 13 30808 89963 31072
rect 13 30528 89120 30808
rect 13 30400 89963 30528
rect 880 30120 89963 30400
rect 13 29992 89963 30120
rect 13 29712 89120 29992
rect 13 29448 89963 29712
rect 880 29168 89963 29448
rect 13 29040 89963 29168
rect 13 28760 89120 29040
rect 13 28496 89963 28760
rect 880 28224 89963 28496
rect 880 28216 89120 28224
rect 13 27944 89120 28216
rect 13 27544 89963 27944
rect 880 27272 89963 27544
rect 880 27264 89120 27272
rect 13 26992 89120 27264
rect 13 26728 89963 26992
rect 880 26456 89963 26728
rect 880 26448 89120 26456
rect 13 26176 89120 26448
rect 13 25776 89963 26176
rect 880 25504 89963 25776
rect 880 25496 89120 25504
rect 13 25224 89120 25496
rect 13 24824 89963 25224
rect 880 24552 89963 24824
rect 880 24544 89120 24552
rect 13 24272 89120 24544
rect 13 23872 89963 24272
rect 880 23736 89963 23872
rect 880 23592 89120 23736
rect 13 23456 89120 23592
rect 13 22920 89963 23456
rect 880 22784 89963 22920
rect 880 22640 89120 22784
rect 13 22504 89120 22640
rect 13 21968 89963 22504
rect 880 21688 89120 21968
rect 13 21016 89963 21688
rect 880 20736 89120 21016
rect 13 20200 89963 20736
rect 880 19920 89120 20200
rect 13 19248 89963 19920
rect 880 18968 89120 19248
rect 13 18432 89963 18968
rect 13 18296 89120 18432
rect 880 18152 89120 18296
rect 880 18016 89963 18152
rect 13 17480 89963 18016
rect 13 17344 89120 17480
rect 880 17200 89120 17344
rect 880 17064 89963 17200
rect 13 16528 89963 17064
rect 13 16392 89120 16528
rect 880 16248 89120 16392
rect 880 16112 89963 16248
rect 13 15712 89963 16112
rect 13 15440 89120 15712
rect 880 15432 89120 15440
rect 880 15160 89963 15432
rect 13 14760 89963 15160
rect 13 14488 89120 14760
rect 880 14480 89120 14488
rect 880 14208 89963 14480
rect 13 13944 89963 14208
rect 13 13672 89120 13944
rect 880 13664 89120 13672
rect 880 13392 89963 13664
rect 13 12992 89963 13392
rect 13 12720 89120 12992
rect 880 12712 89120 12720
rect 880 12440 89963 12712
rect 13 12176 89963 12440
rect 13 11896 89120 12176
rect 13 11768 89963 11896
rect 880 11488 89963 11768
rect 13 11224 89963 11488
rect 13 10944 89120 11224
rect 13 10816 89963 10944
rect 880 10536 89963 10816
rect 13 10408 89963 10536
rect 13 10128 89120 10408
rect 13 9864 89963 10128
rect 880 9584 89963 9864
rect 13 9456 89963 9584
rect 13 9176 89120 9456
rect 13 8912 89963 9176
rect 880 8632 89963 8912
rect 13 8504 89963 8632
rect 13 8224 89120 8504
rect 13 7960 89963 8224
rect 880 7688 89963 7960
rect 880 7680 89120 7688
rect 13 7408 89120 7680
rect 13 7144 89963 7408
rect 880 6864 89963 7144
rect 13 6736 89963 6864
rect 13 6456 89120 6736
rect 13 6192 89963 6456
rect 880 5920 89963 6192
rect 880 5912 89120 5920
rect 13 5640 89120 5912
rect 13 5240 89963 5640
rect 880 4968 89963 5240
rect 880 4960 89120 4968
rect 13 4688 89120 4960
rect 13 4288 89963 4688
rect 880 4152 89963 4288
rect 880 4008 89120 4152
rect 13 3872 89120 4008
rect 13 3336 89963 3872
rect 880 3200 89963 3336
rect 880 3056 89120 3200
rect 13 2920 89120 3056
rect 13 2384 89963 2920
rect 880 2104 89120 2384
rect 13 1432 89963 2104
rect 880 1152 89120 1432
rect 13 616 89963 1152
rect 880 443 89120 616
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
<< obsm4 >>
rect 59 2347 4128 174045
rect 4608 2347 19488 174045
rect 19968 2347 34848 174045
rect 35328 2347 50208 174045
rect 50688 2347 65568 174045
rect 66048 2347 80928 174045
rect 81408 2347 89917 174045
<< labels >>
rlabel metal3 s 0 11568 800 11688 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 addr1[0]
port 10 nsew signal output
rlabel metal3 s 0 113296 800 113416 6 addr1[1]
port 11 nsew signal output
rlabel metal3 s 0 114112 800 114232 6 addr1[2]
port 12 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 addr1[3]
port 13 nsew signal output
rlabel metal3 s 0 116016 800 116136 6 addr1[4]
port 14 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 addr1[5]
port 15 nsew signal output
rlabel metal3 s 0 117920 800 118040 6 addr1[6]
port 16 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 addr1[7]
port 17 nsew signal output
rlabel metal3 s 0 119824 800 119944 6 addr1[8]
port 18 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 clk0
port 19 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 clk1
port 20 nsew signal output
rlabel metal2 s 1122 179200 1178 180000 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 3422 179200 3478 180000 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 5722 179200 5778 180000 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 8022 179200 8078 180000 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 10322 179200 10378 180000 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 12622 179200 12678 180000 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 14922 179200 14978 180000 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 17222 179200 17278 180000 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 89200 2184 90000 2304 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 89200 7488 90000 7608 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 89200 37816 90000 37936 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 89200 40400 90000 40520 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 89200 43120 90000 43240 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 89200 45840 90000 45960 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 89200 48424 90000 48544 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 89200 51144 90000 51264 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 89200 53864 90000 53984 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 89200 56448 90000 56568 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 89200 59168 90000 59288 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 89200 61888 90000 62008 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 89200 11024 90000 11144 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 89200 64472 90000 64592 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 89200 67192 90000 67312 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 89200 69912 90000 70032 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 89200 72496 90000 72616 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 89200 75216 90000 75336 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 89200 77936 90000 78056 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 89200 80520 90000 80640 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 89200 83240 90000 83360 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 89200 14560 90000 14680 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 89200 18232 90000 18352 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 89200 21768 90000 21888 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 89200 24352 90000 24472 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 89200 27072 90000 27192 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 89200 29792 90000 29912 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 89200 32376 90000 32496 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 89200 35096 90000 35216 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 89200 3000 90000 3120 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 89200 8304 90000 8424 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 89200 38632 90000 38752 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 89200 41352 90000 41472 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 89200 44072 90000 44192 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 89200 46656 90000 46776 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 89200 49376 90000 49496 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 89200 52096 90000 52216 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 89200 54680 90000 54800 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 89200 57400 90000 57520 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 89200 60120 90000 60240 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 89200 62704 90000 62824 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 89200 11976 90000 12096 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 89200 65424 90000 65544 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 89200 68144 90000 68264 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 89200 70728 90000 70848 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 89200 73448 90000 73568 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 89200 76168 90000 76288 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 89200 78752 90000 78872 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 89200 81472 90000 81592 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 89200 84192 90000 84312 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 89200 85960 90000 86080 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 89200 87728 90000 87848 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 89200 15512 90000 15632 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 89200 89496 90000 89616 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 89200 91264 90000 91384 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 89200 19048 90000 19168 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 89200 22584 90000 22704 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 89200 25304 90000 25424 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 89200 28024 90000 28144 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 89200 30608 90000 30728 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 89200 33328 90000 33448 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 89200 36048 90000 36168 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 89200 9256 90000 9376 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 89200 39584 90000 39704 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 89200 42304 90000 42424 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 89200 44888 90000 45008 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 89200 47608 90000 47728 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 89200 50328 90000 50448 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 89200 52912 90000 53032 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 89200 55632 90000 55752 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 89200 58352 90000 58472 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 89200 60936 90000 61056 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 89200 63656 90000 63776 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 89200 12792 90000 12912 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 89200 66376 90000 66496 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 89200 68960 90000 69080 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 89200 71680 90000 71800 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 89200 74400 90000 74520 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 89200 76984 90000 77104 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 89200 79704 90000 79824 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 89200 82424 90000 82544 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 89200 85008 90000 85128 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 89200 86776 90000 86896 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 89200 88544 90000 88664 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 89200 16328 90000 16448 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 89200 90448 90000 90568 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 89200 92216 90000 92336 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 89200 20000 90000 20120 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 89200 23536 90000 23656 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 89200 26256 90000 26376 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 89200 28840 90000 28960 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 89200 31560 90000 31680 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 89200 34280 90000 34400 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 89200 36864 90000 36984 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 89200 3952 90000 4072 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 89200 10208 90000 10328 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 89200 13744 90000 13864 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 89200 17280 90000 17400 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 89200 20816 90000 20936 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 89200 4768 90000 4888 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 89200 5720 90000 5840 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 89200 6536 90000 6656 6 core_wb_we_o
port 130 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 csb0[0]
port 131 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 csb0[1]
port 132 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 csb1[1]
port 134 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 din0[0]
port 135 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 din0[10]
port 136 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 din0[11]
port 137 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 din0[12]
port 138 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 din0[13]
port 139 nsew signal output
rlabel metal3 s 0 33056 800 33176 6 din0[14]
port 140 nsew signal output
rlabel metal3 s 0 33872 800 33992 6 din0[15]
port 141 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 din0[16]
port 142 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 din0[17]
port 143 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 din0[18]
port 144 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 din0[19]
port 145 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 din0[1]
port 146 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 din0[20]
port 147 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 din0[21]
port 148 nsew signal output
rlabel metal3 s 0 40400 800 40520 6 din0[22]
port 149 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 din0[23]
port 150 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 din0[24]
port 151 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 din0[25]
port 152 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 din0[26]
port 153 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 din0[27]
port 154 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 din0[28]
port 155 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 din0[29]
port 156 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 din0[2]
port 157 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 din0[30]
port 158 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 din0[31]
port 159 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 din0[3]
port 160 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 din0[4]
port 161 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 din0[5]
port 162 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 din0[6]
port 163 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 din0[7]
port 164 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 din0[8]
port 165 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 din0[9]
port 166 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 dout0[0]
port 167 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 dout0[10]
port 168 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 dout0[11]
port 169 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 dout0[12]
port 170 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 dout0[13]
port 171 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 dout0[14]
port 172 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 dout0[15]
port 173 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 dout0[16]
port 174 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 dout0[17]
port 175 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 dout0[18]
port 176 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 dout0[19]
port 177 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 dout0[1]
port 178 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 dout0[20]
port 179 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 dout0[21]
port 180 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 dout0[22]
port 181 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 dout0[23]
port 182 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 dout0[24]
port 183 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 dout0[25]
port 184 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 dout0[26]
port 185 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 dout0[27]
port 186 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 dout0[28]
port 187 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 dout0[29]
port 188 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 dout0[2]
port 189 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 dout0[30]
port 190 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 dout0[31]
port 191 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 dout0[32]
port 192 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 dout0[33]
port 193 nsew signal input
rlabel metal3 s 0 81472 800 81592 6 dout0[34]
port 194 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 dout0[35]
port 195 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 dout0[36]
port 196 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 dout0[37]
port 197 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 dout0[38]
port 198 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 dout0[39]
port 199 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 dout0[3]
port 200 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 dout0[40]
port 201 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 dout0[41]
port 202 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 dout0[42]
port 203 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 dout0[43]
port 204 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 dout0[44]
port 205 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 dout0[45]
port 206 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 dout0[46]
port 207 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 dout0[47]
port 208 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 dout0[48]
port 209 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 dout0[49]
port 210 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 dout0[4]
port 211 nsew signal input
rlabel metal3 s 0 96432 800 96552 6 dout0[50]
port 212 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 dout0[51]
port 213 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 dout0[52]
port 214 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 dout0[53]
port 215 nsew signal input
rlabel metal3 s 0 100240 800 100360 6 dout0[54]
port 216 nsew signal input
rlabel metal3 s 0 101056 800 101176 6 dout0[55]
port 217 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 dout0[56]
port 218 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 dout0[57]
port 219 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 dout0[58]
port 220 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 dout0[59]
port 221 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 dout0[5]
port 222 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 dout0[60]
port 223 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 dout0[61]
port 224 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 dout0[62]
port 225 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 dout0[63]
port 226 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 dout0[6]
port 227 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 dout0[7]
port 228 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 dout0[8]
port 229 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 dout0[9]
port 230 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 dout1[0]
port 231 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 dout1[10]
port 232 nsew signal input
rlabel metal3 s 0 130976 800 131096 6 dout1[11]
port 233 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 dout1[12]
port 234 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 dout1[13]
port 235 nsew signal input
rlabel metal3 s 0 133696 800 133816 6 dout1[14]
port 236 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 dout1[15]
port 237 nsew signal input
rlabel metal3 s 0 135600 800 135720 6 dout1[16]
port 238 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 dout1[17]
port 239 nsew signal input
rlabel metal3 s 0 137504 800 137624 6 dout1[18]
port 240 nsew signal input
rlabel metal3 s 0 138456 800 138576 6 dout1[19]
port 241 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 dout1[1]
port 242 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 dout1[20]
port 243 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 dout1[21]
port 244 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 dout1[22]
port 245 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 dout1[23]
port 246 nsew signal input
rlabel metal3 s 0 143080 800 143200 6 dout1[24]
port 247 nsew signal input
rlabel metal3 s 0 144032 800 144152 6 dout1[25]
port 248 nsew signal input
rlabel metal3 s 0 144984 800 145104 6 dout1[26]
port 249 nsew signal input
rlabel metal3 s 0 145936 800 146056 6 dout1[27]
port 250 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 dout1[28]
port 251 nsew signal input
rlabel metal3 s 0 147704 800 147824 6 dout1[29]
port 252 nsew signal input
rlabel metal3 s 0 122544 800 122664 6 dout1[2]
port 253 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 dout1[30]
port 254 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 dout1[31]
port 255 nsew signal input
rlabel metal3 s 0 150560 800 150680 6 dout1[32]
port 256 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 dout1[33]
port 257 nsew signal input
rlabel metal3 s 0 152464 800 152584 6 dout1[34]
port 258 nsew signal input
rlabel metal3 s 0 153416 800 153536 6 dout1[35]
port 259 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 dout1[36]
port 260 nsew signal input
rlabel metal3 s 0 155184 800 155304 6 dout1[37]
port 261 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 dout1[38]
port 262 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 dout1[39]
port 263 nsew signal input
rlabel metal3 s 0 123496 800 123616 6 dout1[3]
port 264 nsew signal input
rlabel metal3 s 0 158040 800 158160 6 dout1[40]
port 265 nsew signal input
rlabel metal3 s 0 158992 800 159112 6 dout1[41]
port 266 nsew signal input
rlabel metal3 s 0 159944 800 160064 6 dout1[42]
port 267 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 dout1[43]
port 268 nsew signal input
rlabel metal3 s 0 161712 800 161832 6 dout1[44]
port 269 nsew signal input
rlabel metal3 s 0 162664 800 162784 6 dout1[45]
port 270 nsew signal input
rlabel metal3 s 0 163616 800 163736 6 dout1[46]
port 271 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 dout1[47]
port 272 nsew signal input
rlabel metal3 s 0 165520 800 165640 6 dout1[48]
port 273 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 dout1[49]
port 274 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 dout1[4]
port 275 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 dout1[50]
port 276 nsew signal input
rlabel metal3 s 0 168240 800 168360 6 dout1[51]
port 277 nsew signal input
rlabel metal3 s 0 169192 800 169312 6 dout1[52]
port 278 nsew signal input
rlabel metal3 s 0 170144 800 170264 6 dout1[53]
port 279 nsew signal input
rlabel metal3 s 0 171096 800 171216 6 dout1[54]
port 280 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 dout1[55]
port 281 nsew signal input
rlabel metal3 s 0 173000 800 173120 6 dout1[56]
port 282 nsew signal input
rlabel metal3 s 0 173816 800 173936 6 dout1[57]
port 283 nsew signal input
rlabel metal3 s 0 174768 800 174888 6 dout1[58]
port 284 nsew signal input
rlabel metal3 s 0 175720 800 175840 6 dout1[59]
port 285 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 dout1[5]
port 286 nsew signal input
rlabel metal3 s 0 176672 800 176792 6 dout1[60]
port 287 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 dout1[61]
port 288 nsew signal input
rlabel metal3 s 0 178576 800 178696 6 dout1[62]
port 289 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 dout1[63]
port 290 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 dout1[6]
port 291 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 dout1[7]
port 292 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 dout1[8]
port 293 nsew signal input
rlabel metal3 s 0 129072 800 129192 6 dout1[9]
port 294 nsew signal input
rlabel metal3 s 0 416 800 536 6 jtag_tck
port 295 nsew signal input
rlabel metal3 s 0 1232 800 1352 6 jtag_tdi
port 296 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 jtag_tdo
port 297 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 jtag_tms
port 298 nsew signal input
rlabel metal3 s 89200 93032 90000 93152 6 localMemory_wb_ack_o
port 299 nsew signal output
rlabel metal3 s 89200 98336 90000 98456 6 localMemory_wb_adr_i[0]
port 300 nsew signal input
rlabel metal3 s 89200 128664 90000 128784 6 localMemory_wb_adr_i[10]
port 301 nsew signal input
rlabel metal3 s 89200 131384 90000 131504 6 localMemory_wb_adr_i[11]
port 302 nsew signal input
rlabel metal3 s 89200 134104 90000 134224 6 localMemory_wb_adr_i[12]
port 303 nsew signal input
rlabel metal3 s 89200 136688 90000 136808 6 localMemory_wb_adr_i[13]
port 304 nsew signal input
rlabel metal3 s 89200 139408 90000 139528 6 localMemory_wb_adr_i[14]
port 305 nsew signal input
rlabel metal3 s 89200 142128 90000 142248 6 localMemory_wb_adr_i[15]
port 306 nsew signal input
rlabel metal3 s 89200 144712 90000 144832 6 localMemory_wb_adr_i[16]
port 307 nsew signal input
rlabel metal3 s 89200 147432 90000 147552 6 localMemory_wb_adr_i[17]
port 308 nsew signal input
rlabel metal3 s 89200 150152 90000 150272 6 localMemory_wb_adr_i[18]
port 309 nsew signal input
rlabel metal3 s 89200 152736 90000 152856 6 localMemory_wb_adr_i[19]
port 310 nsew signal input
rlabel metal3 s 89200 102008 90000 102128 6 localMemory_wb_adr_i[1]
port 311 nsew signal input
rlabel metal3 s 89200 155456 90000 155576 6 localMemory_wb_adr_i[20]
port 312 nsew signal input
rlabel metal3 s 89200 158176 90000 158296 6 localMemory_wb_adr_i[21]
port 313 nsew signal input
rlabel metal3 s 89200 160760 90000 160880 6 localMemory_wb_adr_i[22]
port 314 nsew signal input
rlabel metal3 s 89200 163480 90000 163600 6 localMemory_wb_adr_i[23]
port 315 nsew signal input
rlabel metal3 s 89200 105544 90000 105664 6 localMemory_wb_adr_i[2]
port 316 nsew signal input
rlabel metal3 s 89200 109080 90000 109200 6 localMemory_wb_adr_i[3]
port 317 nsew signal input
rlabel metal3 s 89200 112616 90000 112736 6 localMemory_wb_adr_i[4]
port 318 nsew signal input
rlabel metal3 s 89200 115336 90000 115456 6 localMemory_wb_adr_i[5]
port 319 nsew signal input
rlabel metal3 s 89200 118056 90000 118176 6 localMemory_wb_adr_i[6]
port 320 nsew signal input
rlabel metal3 s 89200 120640 90000 120760 6 localMemory_wb_adr_i[7]
port 321 nsew signal input
rlabel metal3 s 89200 123360 90000 123480 6 localMemory_wb_adr_i[8]
port 322 nsew signal input
rlabel metal3 s 89200 126080 90000 126200 6 localMemory_wb_adr_i[9]
port 323 nsew signal input
rlabel metal3 s 89200 93984 90000 94104 6 localMemory_wb_cyc_i
port 324 nsew signal input
rlabel metal3 s 89200 99288 90000 99408 6 localMemory_wb_data_i[0]
port 325 nsew signal input
rlabel metal3 s 89200 129616 90000 129736 6 localMemory_wb_data_i[10]
port 326 nsew signal input
rlabel metal3 s 89200 132336 90000 132456 6 localMemory_wb_data_i[11]
port 327 nsew signal input
rlabel metal3 s 89200 134920 90000 135040 6 localMemory_wb_data_i[12]
port 328 nsew signal input
rlabel metal3 s 89200 137640 90000 137760 6 localMemory_wb_data_i[13]
port 329 nsew signal input
rlabel metal3 s 89200 140360 90000 140480 6 localMemory_wb_data_i[14]
port 330 nsew signal input
rlabel metal3 s 89200 142944 90000 143064 6 localMemory_wb_data_i[15]
port 331 nsew signal input
rlabel metal3 s 89200 145664 90000 145784 6 localMemory_wb_data_i[16]
port 332 nsew signal input
rlabel metal3 s 89200 148384 90000 148504 6 localMemory_wb_data_i[17]
port 333 nsew signal input
rlabel metal3 s 89200 150968 90000 151088 6 localMemory_wb_data_i[18]
port 334 nsew signal input
rlabel metal3 s 89200 153688 90000 153808 6 localMemory_wb_data_i[19]
port 335 nsew signal input
rlabel metal3 s 89200 102824 90000 102944 6 localMemory_wb_data_i[1]
port 336 nsew signal input
rlabel metal3 s 89200 156408 90000 156528 6 localMemory_wb_data_i[20]
port 337 nsew signal input
rlabel metal3 s 89200 158992 90000 159112 6 localMemory_wb_data_i[21]
port 338 nsew signal input
rlabel metal3 s 89200 161712 90000 161832 6 localMemory_wb_data_i[22]
port 339 nsew signal input
rlabel metal3 s 89200 164432 90000 164552 6 localMemory_wb_data_i[23]
port 340 nsew signal input
rlabel metal3 s 89200 166200 90000 166320 6 localMemory_wb_data_i[24]
port 341 nsew signal input
rlabel metal3 s 89200 167968 90000 168088 6 localMemory_wb_data_i[25]
port 342 nsew signal input
rlabel metal3 s 89200 169736 90000 169856 6 localMemory_wb_data_i[26]
port 343 nsew signal input
rlabel metal3 s 89200 171504 90000 171624 6 localMemory_wb_data_i[27]
port 344 nsew signal input
rlabel metal3 s 89200 173272 90000 173392 6 localMemory_wb_data_i[28]
port 345 nsew signal input
rlabel metal3 s 89200 175040 90000 175160 6 localMemory_wb_data_i[29]
port 346 nsew signal input
rlabel metal3 s 89200 106360 90000 106480 6 localMemory_wb_data_i[2]
port 347 nsew signal input
rlabel metal3 s 89200 176808 90000 176928 6 localMemory_wb_data_i[30]
port 348 nsew signal input
rlabel metal3 s 89200 178576 90000 178696 6 localMemory_wb_data_i[31]
port 349 nsew signal input
rlabel metal3 s 89200 110032 90000 110152 6 localMemory_wb_data_i[3]
port 350 nsew signal input
rlabel metal3 s 89200 113568 90000 113688 6 localMemory_wb_data_i[4]
port 351 nsew signal input
rlabel metal3 s 89200 116288 90000 116408 6 localMemory_wb_data_i[5]
port 352 nsew signal input
rlabel metal3 s 89200 118872 90000 118992 6 localMemory_wb_data_i[6]
port 353 nsew signal input
rlabel metal3 s 89200 121592 90000 121712 6 localMemory_wb_data_i[7]
port 354 nsew signal input
rlabel metal3 s 89200 124312 90000 124432 6 localMemory_wb_data_i[8]
port 355 nsew signal input
rlabel metal3 s 89200 126896 90000 127016 6 localMemory_wb_data_i[9]
port 356 nsew signal input
rlabel metal3 s 89200 100240 90000 100360 6 localMemory_wb_data_o[0]
port 357 nsew signal output
rlabel metal3 s 89200 130432 90000 130552 6 localMemory_wb_data_o[10]
port 358 nsew signal output
rlabel metal3 s 89200 133152 90000 133272 6 localMemory_wb_data_o[11]
port 359 nsew signal output
rlabel metal3 s 89200 135872 90000 135992 6 localMemory_wb_data_o[12]
port 360 nsew signal output
rlabel metal3 s 89200 138456 90000 138576 6 localMemory_wb_data_o[13]
port 361 nsew signal output
rlabel metal3 s 89200 141176 90000 141296 6 localMemory_wb_data_o[14]
port 362 nsew signal output
rlabel metal3 s 89200 143896 90000 144016 6 localMemory_wb_data_o[15]
port 363 nsew signal output
rlabel metal3 s 89200 146480 90000 146600 6 localMemory_wb_data_o[16]
port 364 nsew signal output
rlabel metal3 s 89200 149200 90000 149320 6 localMemory_wb_data_o[17]
port 365 nsew signal output
rlabel metal3 s 89200 151920 90000 152040 6 localMemory_wb_data_o[18]
port 366 nsew signal output
rlabel metal3 s 89200 154504 90000 154624 6 localMemory_wb_data_o[19]
port 367 nsew signal output
rlabel metal3 s 89200 103776 90000 103896 6 localMemory_wb_data_o[1]
port 368 nsew signal output
rlabel metal3 s 89200 157224 90000 157344 6 localMemory_wb_data_o[20]
port 369 nsew signal output
rlabel metal3 s 89200 159944 90000 160064 6 localMemory_wb_data_o[21]
port 370 nsew signal output
rlabel metal3 s 89200 162528 90000 162648 6 localMemory_wb_data_o[22]
port 371 nsew signal output
rlabel metal3 s 89200 165248 90000 165368 6 localMemory_wb_data_o[23]
port 372 nsew signal output
rlabel metal3 s 89200 167016 90000 167136 6 localMemory_wb_data_o[24]
port 373 nsew signal output
rlabel metal3 s 89200 168784 90000 168904 6 localMemory_wb_data_o[25]
port 374 nsew signal output
rlabel metal3 s 89200 170552 90000 170672 6 localMemory_wb_data_o[26]
port 375 nsew signal output
rlabel metal3 s 89200 172456 90000 172576 6 localMemory_wb_data_o[27]
port 376 nsew signal output
rlabel metal3 s 89200 174224 90000 174344 6 localMemory_wb_data_o[28]
port 377 nsew signal output
rlabel metal3 s 89200 175992 90000 176112 6 localMemory_wb_data_o[29]
port 378 nsew signal output
rlabel metal3 s 89200 107312 90000 107432 6 localMemory_wb_data_o[2]
port 379 nsew signal output
rlabel metal3 s 89200 177760 90000 177880 6 localMemory_wb_data_o[30]
port 380 nsew signal output
rlabel metal3 s 89200 179528 90000 179648 6 localMemory_wb_data_o[31]
port 381 nsew signal output
rlabel metal3 s 89200 110848 90000 110968 6 localMemory_wb_data_o[3]
port 382 nsew signal output
rlabel metal3 s 89200 114384 90000 114504 6 localMemory_wb_data_o[4]
port 383 nsew signal output
rlabel metal3 s 89200 117104 90000 117224 6 localMemory_wb_data_o[5]
port 384 nsew signal output
rlabel metal3 s 89200 119824 90000 119944 6 localMemory_wb_data_o[6]
port 385 nsew signal output
rlabel metal3 s 89200 122408 90000 122528 6 localMemory_wb_data_o[7]
port 386 nsew signal output
rlabel metal3 s 89200 125128 90000 125248 6 localMemory_wb_data_o[8]
port 387 nsew signal output
rlabel metal3 s 89200 127848 90000 127968 6 localMemory_wb_data_o[9]
port 388 nsew signal output
rlabel metal3 s 89200 94800 90000 94920 6 localMemory_wb_error_o
port 389 nsew signal output
rlabel metal3 s 89200 101056 90000 101176 6 localMemory_wb_sel_i[0]
port 390 nsew signal input
rlabel metal3 s 89200 104592 90000 104712 6 localMemory_wb_sel_i[1]
port 391 nsew signal input
rlabel metal3 s 89200 108264 90000 108384 6 localMemory_wb_sel_i[2]
port 392 nsew signal input
rlabel metal3 s 89200 111800 90000 111920 6 localMemory_wb_sel_i[3]
port 393 nsew signal input
rlabel metal3 s 89200 95752 90000 95872 6 localMemory_wb_stall_o
port 394 nsew signal output
rlabel metal3 s 89200 96568 90000 96688 6 localMemory_wb_stb_i
port 395 nsew signal input
rlabel metal3 s 89200 97520 90000 97640 6 localMemory_wb_we_i
port 396 nsew signal input
rlabel metal2 s 19522 179200 19578 180000 6 manufacturerID[0]
port 397 nsew signal input
rlabel metal2 s 42614 179200 42670 180000 6 manufacturerID[10]
port 398 nsew signal input
rlabel metal2 s 21822 179200 21878 180000 6 manufacturerID[1]
port 399 nsew signal input
rlabel metal2 s 24122 179200 24178 180000 6 manufacturerID[2]
port 400 nsew signal input
rlabel metal2 s 26422 179200 26478 180000 6 manufacturerID[3]
port 401 nsew signal input
rlabel metal2 s 28722 179200 28778 180000 6 manufacturerID[4]
port 402 nsew signal input
rlabel metal2 s 31114 179200 31170 180000 6 manufacturerID[5]
port 403 nsew signal input
rlabel metal2 s 33414 179200 33470 180000 6 manufacturerID[6]
port 404 nsew signal input
rlabel metal2 s 35714 179200 35770 180000 6 manufacturerID[7]
port 405 nsew signal input
rlabel metal2 s 38014 179200 38070 180000 6 manufacturerID[8]
port 406 nsew signal input
rlabel metal2 s 40314 179200 40370 180000 6 manufacturerID[9]
port 407 nsew signal input
rlabel metal2 s 44914 179200 44970 180000 6 partID[0]
port 408 nsew signal input
rlabel metal2 s 68006 179200 68062 180000 6 partID[10]
port 409 nsew signal input
rlabel metal2 s 70306 179200 70362 180000 6 partID[11]
port 410 nsew signal input
rlabel metal2 s 72606 179200 72662 180000 6 partID[12]
port 411 nsew signal input
rlabel metal2 s 74906 179200 74962 180000 6 partID[13]
port 412 nsew signal input
rlabel metal2 s 77206 179200 77262 180000 6 partID[14]
port 413 nsew signal input
rlabel metal2 s 79506 179200 79562 180000 6 partID[15]
port 414 nsew signal input
rlabel metal2 s 47214 179200 47270 180000 6 partID[1]
port 415 nsew signal input
rlabel metal2 s 49514 179200 49570 180000 6 partID[2]
port 416 nsew signal input
rlabel metal2 s 51814 179200 51870 180000 6 partID[3]
port 417 nsew signal input
rlabel metal2 s 54114 179200 54170 180000 6 partID[4]
port 418 nsew signal input
rlabel metal2 s 56414 179200 56470 180000 6 partID[5]
port 419 nsew signal input
rlabel metal2 s 58714 179200 58770 180000 6 partID[6]
port 420 nsew signal input
rlabel metal2 s 61106 179200 61162 180000 6 partID[7]
port 421 nsew signal input
rlabel metal2 s 63406 179200 63462 180000 6 partID[8]
port 422 nsew signal input
rlabel metal2 s 65706 179200 65762 180000 6 partID[9]
port 423 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 probe_errorCode[0]
port 424 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 probe_errorCode[1]
port 425 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 probe_errorCode[2]
port 426 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 probe_errorCode[3]
port 427 nsew signal output
rlabel metal2 s 754 0 810 800 6 probe_isBranch
port 428 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 probe_isCompressed
port 429 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 probe_isLoad
port 430 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 probe_isStore
port 431 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 probe_jtagInstruction[0]
port 432 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 probe_jtagInstruction[1]
port 433 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 probe_jtagInstruction[2]
port 434 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 probe_jtagInstruction[3]
port 435 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 probe_jtagInstruction[4]
port 436 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 probe_opcode[0]
port 437 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 probe_opcode[1]
port 438 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 probe_opcode[2]
port 439 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 probe_opcode[3]
port 440 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 probe_opcode[4]
port 441 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 probe_opcode[5]
port 442 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 probe_opcode[6]
port 443 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 probe_programCounter[0]
port 444 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 probe_programCounter[10]
port 445 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 probe_programCounter[11]
port 446 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 probe_programCounter[12]
port 447 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 probe_programCounter[13]
port 448 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 probe_programCounter[14]
port 449 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 probe_programCounter[15]
port 450 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 probe_programCounter[16]
port 451 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 probe_programCounter[17]
port 452 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 probe_programCounter[18]
port 453 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 probe_programCounter[19]
port 454 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 probe_programCounter[1]
port 455 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 probe_programCounter[20]
port 456 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 probe_programCounter[21]
port 457 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 probe_programCounter[22]
port 458 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 probe_programCounter[23]
port 459 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 probe_programCounter[24]
port 460 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 probe_programCounter[25]
port 461 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 probe_programCounter[26]
port 462 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 probe_programCounter[27]
port 463 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 probe_programCounter[28]
port 464 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 probe_programCounter[29]
port 465 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 probe_programCounter[2]
port 466 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 probe_programCounter[30]
port 467 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 probe_programCounter[31]
port 468 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 probe_programCounter[3]
port 469 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 probe_programCounter[4]
port 470 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 probe_programCounter[5]
port 471 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 probe_programCounter[6]
port 472 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 probe_programCounter[7]
port 473 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 probe_programCounter[8]
port 474 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 probe_programCounter[9]
port 475 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 probe_state[0]
port 476 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 probe_state[1]
port 477 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 probe_takeBranch
port 478 nsew signal output
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 479 nsew power bidirectional
rlabel metal2 s 81806 179200 81862 180000 6 versionID[0]
port 480 nsew signal input
rlabel metal2 s 84106 179200 84162 180000 6 versionID[1]
port 481 nsew signal input
rlabel metal2 s 86406 179200 86462 180000 6 versionID[2]
port 482 nsew signal input
rlabel metal2 s 88706 179200 88762 180000 6 versionID[3]
port 483 nsew signal input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 484 nsew ground bidirectional
rlabel metal3 s 89200 416 90000 536 6 wb_clk_i
port 485 nsew signal input
rlabel metal3 s 89200 1232 90000 1352 6 wb_rst_i
port 486 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 web0
port 487 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 wmask0[0]
port 488 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 wmask0[1]
port 489 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 wmask0[2]
port 490 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 wmask0[3]
port 491 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 90000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 52602258
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/signoff/ExperiarCore.magic.gds
string GDS_START 1485086
<< end >>

