* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

.subckt CaravelHost caravel_irq[0] caravel_irq[1] caravel_irq[2] caravel_irq[3] caravel_uart_rx
+ caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0] caravel_wb_adr_o[10] caravel_wb_adr_o[11]
+ caravel_wb_adr_o[12] caravel_wb_adr_o[13] caravel_wb_adr_o[14] caravel_wb_adr_o[15]
+ caravel_wb_adr_o[16] caravel_wb_adr_o[17] caravel_wb_adr_o[18] caravel_wb_adr_o[19]
+ caravel_wb_adr_o[1] caravel_wb_adr_o[20] caravel_wb_adr_o[21] caravel_wb_adr_o[22]
+ caravel_wb_adr_o[23] caravel_wb_adr_o[24] caravel_wb_adr_o[25] caravel_wb_adr_o[26]
+ caravel_wb_adr_o[27] caravel_wb_adr_o[2] caravel_wb_adr_o[3] caravel_wb_adr_o[4]
+ caravel_wb_adr_o[5] caravel_wb_adr_o[6] caravel_wb_adr_o[7] caravel_wb_adr_o[8]
+ caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0] caravel_wb_data_i[10]
+ caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13] caravel_wb_data_i[14]
+ caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17] caravel_wb_data_i[18]
+ caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20] caravel_wb_data_i[21]
+ caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24] caravel_wb_data_i[25]
+ caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28] caravel_wb_data_i[29]
+ caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31] caravel_wb_data_i[3]
+ caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6] caravel_wb_data_i[7]
+ caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0] caravel_wb_data_o[10]
+ caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13] caravel_wb_data_o[14]
+ caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17] caravel_wb_data_o[18]
+ caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20] caravel_wb_data_o[21]
+ caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24] caravel_wb_data_o[25]
+ caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28] caravel_wb_data_o[29]
+ caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31] caravel_wb_data_o[3]
+ caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6] caravel_wb_data_o[7]
+ caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i caravel_wb_sel_o[0]
+ caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3] caravel_wb_stall_i caravel_wb_stb_o
+ caravel_wb_we_o core0Index[0] core0Index[1] core0Index[2] core0Index[3] core0Index[4]
+ core0Index[5] core0Index[6] core0Index[7] core1Index[0] core1Index[1] core1Index[2]
+ core1Index[3] core1Index[4] core1Index[5] core1Index[6] core1Index[7] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] manufacturerID[0]
+ manufacturerID[10] manufacturerID[1] manufacturerID[2] manufacturerID[3] manufacturerID[4]
+ manufacturerID[5] manufacturerID[6] manufacturerID[7] manufacturerID[8] manufacturerID[9]
+ partID[0] partID[10] partID[11] partID[12] partID[13] partID[14] partID[15] partID[1]
+ partID[2] partID[3] partID[4] partID[5] partID[6] partID[7] partID[8] partID[9]
+ probe_out[0] probe_out[10] probe_out[11] probe_out[12] probe_out[13] probe_out[14]
+ probe_out[15] probe_out[16] probe_out[17] probe_out[18] probe_out[19] probe_out[1]
+ probe_out[20] probe_out[21] probe_out[22] probe_out[23] probe_out[24] probe_out[25]
+ probe_out[26] probe_out[27] probe_out[28] probe_out[29] probe_out[2] probe_out[30]
+ probe_out[31] probe_out[32] probe_out[33] probe_out[34] probe_out[35] probe_out[36]
+ probe_out[37] probe_out[38] probe_out[39] probe_out[3] probe_out[40] probe_out[41]
+ probe_out[42] probe_out[43] probe_out[44] probe_out[45] probe_out[46] probe_out[47]
+ probe_out[48] probe_out[49] probe_out[4] probe_out[50] probe_out[51] probe_out[52]
+ probe_out[53] probe_out[54] probe_out[55] probe_out[56] probe_out[57] probe_out[58]
+ probe_out[59] probe_out[5] probe_out[60] probe_out[61] probe_out[62] probe_out[63]
+ probe_out[64] probe_out[65] probe_out[66] probe_out[67] probe_out[68] probe_out[69]
+ probe_out[6] probe_out[70] probe_out[71] probe_out[72] probe_out[73] probe_out[74]
+ probe_out[75] probe_out[76] probe_out[77] probe_out[78] probe_out[79] probe_out[7]
+ probe_out[80] probe_out[81] probe_out[82] probe_out[83] probe_out[84] probe_out[85]
+ probe_out[86] probe_out[87] probe_out[88] probe_out[89] probe_out[8] probe_out[90]
+ probe_out[91] probe_out[92] probe_out[93] probe_out[94] probe_out[95] probe_out[96]
+ probe_out[97] probe_out[9] vccd1 versionID[0] versionID[1] versionID[2] versionID[3]
+ vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_data_i[0] wbs_data_i[10]
+ wbs_data_i[11] wbs_data_i[12] wbs_data_i[13] wbs_data_i[14] wbs_data_i[15] wbs_data_i[16]
+ wbs_data_i[17] wbs_data_i[18] wbs_data_i[19] wbs_data_i[1] wbs_data_i[20] wbs_data_i[21]
+ wbs_data_i[22] wbs_data_i[23] wbs_data_i[24] wbs_data_i[25] wbs_data_i[26] wbs_data_i[27]
+ wbs_data_i[28] wbs_data_i[29] wbs_data_i[2] wbs_data_i[30] wbs_data_i[31] wbs_data_i[3]
+ wbs_data_i[4] wbs_data_i[5] wbs_data_i[6] wbs_data_i[7] wbs_data_i[8] wbs_data_i[9]
+ wbs_data_o[0] wbs_data_o[10] wbs_data_o[11] wbs_data_o[12] wbs_data_o[13] wbs_data_o[14]
+ wbs_data_o[15] wbs_data_o[16] wbs_data_o[17] wbs_data_o[18] wbs_data_o[19] wbs_data_o[1]
+ wbs_data_o[20] wbs_data_o[21] wbs_data_o[22] wbs_data_o[23] wbs_data_o[24] wbs_data_o[25]
+ wbs_data_o[26] wbs_data_o[27] wbs_data_o[28] wbs_data_o[29] wbs_data_o[2] wbs_data_o[30]
+ wbs_data_o[31] wbs_data_o[3] wbs_data_o[4] wbs_data_o[5] wbs_data_o[6] wbs_data_o[7]
+ wbs_data_o[8] wbs_data_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3155_ _3136_/X _3152_/X _3154_/X _3150_/X vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__a31o_1
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3086_ _3443_/B _3089_/A _2778_/A vssd1 vssd1 vccd1 vccd1 _3087_/B sky130_fd_sc_hd__o21ai_1
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _3652_/A _5257_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _5257_/D sky130_fd_sc_hd__mux2_1
X_2939_ _5587_/Q _5571_/Q _5453_/Q _5603_/Q _3063_/S _2867_/B vssd1 vssd1 vccd1 vccd1
+ _2939_/X sky130_fd_sc_hd__mux4_2
X_5727_ _5733_/CLK _5727_/D vssd1 vssd1 vccd1 vccd1 _5727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5658_ _5658_/CLK _5658_/D vssd1 vssd1 vccd1 vccd1 _5658_/Q sky130_fd_sc_hd__dfxtp_1
X_5589_ _5589_/CLK _5589_/D vssd1 vssd1 vccd1 vccd1 _5589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold351 hold374/X vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__buf_2
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold395 _3966_/X vssd1 vssd1 vccd1 vccd1 _5205_/D sky130_fd_sc_hd__buf_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4476__61 _4478__63/A vssd1 vssd1 vccd1 vccd1 _5118_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1040 hold1650/X vssd1 vssd1 vccd1 vccd1 hold1651/A sky130_fd_sc_hd__buf_2
Xhold1051 hold1836/X vssd1 vssd1 vccd1 vccd1 hold1837/A sky130_fd_sc_hd__buf_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1073 hold1832/X vssd1 vssd1 vccd1 vccd1 hold1833/A sky130_fd_sc_hd__buf_2
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4960__545 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5718_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _5259_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3911_ _5079_/Q _3926_/A2 _3923_/B1 _3910_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5079_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3842_ _5089_/Q _5097_/Q _5098_/Q vssd1 vssd1 vccd1 vccd1 _3850_/C sky130_fd_sc_hd__or3_2
XFILLER_146_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3773_ _3773_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__and2_1
X_5512_ _5512_/CLK _5512_/D vssd1 vssd1 vccd1 vccd1 _5512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2724_ _2790_/A0 _5503_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5503_/D sky130_fd_sc_hd__mux2_1
X_2655_ _2779_/A _3589_/A vssd1 vssd1 vccd1 vccd1 _2663_/S sky130_fd_sc_hd__or2_4
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4597__182 _4964__549/A vssd1 vssd1 vccd1 vccd1 _5271_/CLK sky130_fd_sc_hd__inv_2
Xoutput401 _3709_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__clkbuf_2
X_5443_ _5443_/CLK _5443_/D vssd1 vssd1 vccd1 vccd1 _5443_/Q sky130_fd_sc_hd__dfxtp_1
X_5374_ _5374_/CLK _5374_/D vssd1 vssd1 vccd1 vccd1 _5374_/Q sky130_fd_sc_hd__dfxtp_1
X_4325_ _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4325_/Y sky130_fd_sc_hd__nor2_1
X_2586_ _3562_/A _3388_/B vssd1 vssd1 vccd1 vccd1 _2594_/S sky130_fd_sc_hd__or2_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4256_ _5746_/Q _4039_/X _4254_/X _4255_/Y vssd1 vssd1 vccd1 vccd1 _4265_/C sky130_fd_sc_hd__o22a_1
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4187_ _4181_/B _4137_/B _4184_/Y _4187_/B1 _5540_/Q vssd1 vssd1 vccd1 vccd1 _4188_/B
+ sky130_fd_sc_hd__a32oi_4
X_3207_ _3326_/C1 _3204_/X _3206_/X vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4944__529 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5702_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3138_ _5329_/Q _3138_/B vssd1 vssd1 vccd1 vccd1 _3140_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3069_ _5393_/Q _5401_/Q _3069_/S vssd1 vssd1 vccd1 vccd1 _3069_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4838__423 _4424__9/A vssd1 vssd1 vccd1 vccd1 _5531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__buf_2
XFILLER_132_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__buf_2
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__buf_2
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout650 input134/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__buf_12
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2440_ _5678_/Q vssd1 vssd1 vccd1 vccd1 _4013_/B sky130_fd_sc_hd__inv_2
XFILLER_123_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1809 hold2540/X vssd1 vssd1 vccd1 vccd1 hold2541/A sky130_fd_sc_hd__buf_2
X_5090_ _5291_/CLK _5090_/D vssd1 vssd1 vccd1 vccd1 _5090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4631__216 _4460__45/A vssd1 vssd1 vccd1 vccd1 _5308_/CLK sky130_fd_sc_hd__inv_2
X_4110_ _5744_/Q _4110_/B vssd1 vssd1 vccd1 vccd1 _4170_/A sky130_fd_sc_hd__xor2_1
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4041_ _4253_/A _4041_/B _4041_/C vssd1 vssd1 vccd1 vccd1 _4041_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4525__110 _4477__62/A vssd1 vssd1 vccd1 vccd1 _5167_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3825_ _5024_/Q _3825_/A2 _4368_/A vssd1 vssd1 vccd1 vccd1 _3825_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3756_ _5005_/Q _3750_/B _3774_/B1 _3755_/X _3774_/C1 vssd1 vssd1 vccd1 vccd1 _3756_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2707_ _3392_/A0 _5517_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5517_/D sky130_fd_sc_hd__mux2_1
X_3687_ _5260_/Q _3688_/B vssd1 vssd1 vccd1 vccd1 _3687_/X sky130_fd_sc_hd__and2_1
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5426_ _5426_/CLK _5426_/D vssd1 vssd1 vccd1 vccd1 _5426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput242 _3644_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput231 _3667_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput253 _3654_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__clkbuf_2
Xoutput220 _3682_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__clkbuf_2
X_2638_ _5605_/Q _3600_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5605_/D sky130_fd_sc_hd__mux2_1
Xoutput264 _3635_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__clkbuf_2
X_5357_ _5357_/CLK _5357_/D vssd1 vssd1 vccd1 vccd1 _5357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2569_ _2743_/A0 _5644_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5644_/D sky130_fd_sc_hd__mux2_1
Xoutput286 _5857_/X vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_12
Xoutput275 _5847_/X vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_12
XFILLER_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4308_ _4249_/B _4308_/A2 _4308_/B1 _2444_/Y vssd1 vssd1 vccd1 vccd1 _4308_/X sky130_fd_sc_hd__o22a_1
X_5288_ _5288_/CLK _5288_/D vssd1 vssd1 vccd1 vccd1 _5288_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput297 _5867_/X vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_12
XFILLER_101_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4239_ _5342_/Q _3124_/Y _4164_/B _4238_/X _4244_/S vssd1 vssd1 vccd1 vccd1 _5563_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_114_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4446__31 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5040_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout480 _3099_/B vssd1 vssd1 vccd1 vccd1 _3041_/B1 sky130_fd_sc_hd__buf_6
Xfanout491 hold364/A vssd1 vssd1 vccd1 vccd1 hold349/A sky130_fd_sc_hd__clkbuf_8
XFILLER_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3610_ _4972_/Q _3610_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4972_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3541_ _3604_/A1 _5124_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5124_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3472_ _3508_/A _3607_/B vssd1 vssd1 vccd1 vccd1 _3480_/S sky130_fd_sc_hd__or2_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5211_ _5211_/CLK _5211_/D vssd1 vssd1 vccd1 vccd1 _5211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5142_ _5142_/CLK _5142_/D vssd1 vssd1 vccd1 vccd1 _5142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2318 hold2318/A vssd1 vssd1 vccd1 vccd1 hold2318/X sky130_fd_sc_hd__buf_2
Xhold2307 hold717/X vssd1 vssd1 vccd1 vccd1 hold2307/X sky130_fd_sc_hd__buf_2
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1606 hold44/X vssd1 vssd1 vccd1 vccd1 hold1606/X sky130_fd_sc_hd__buf_2
Xhold1617 hold1617/A vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__buf_2
Xhold2329 hold2329/A vssd1 vssd1 vccd1 vccd1 hold992/A sky130_fd_sc_hd__buf_2
Xhold1628 hold2826/X vssd1 vssd1 vccd1 vccd1 hold2203/A sky130_fd_sc_hd__buf_2
X_5073_ _5752_/CLK _5073_/D vssd1 vssd1 vccd1 vccd1 _5073_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1639 hold2804/X vssd1 vssd1 vccd1 vccd1 hold2805/A sky130_fd_sc_hd__buf_2
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4024_ _4024_/A _4247_/B _4247_/C vssd1 vssd1 vccd1 vccd1 _4026_/C sky130_fd_sc_hd__and3_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3808_ _5259_/Q hold358/X _3810_/A3 hold349/X _5008_/Q vssd1 vssd1 vccd1 vccd1 _3808_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4800__385 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5491_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3739_ _3824_/A1 _3737_/X _3738_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3739_/X sky130_fd_sc_hd__o211a_4
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5409_ _5409_/CLK _5409_/D vssd1 vssd1 vccd1 vccd1 _5409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2885 hold2885/A vssd1 vssd1 vccd1 vccd1 hold2885/X sky130_fd_sc_hd__buf_2
XFILLER_56_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_117_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4937__522/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4743__328 _4744__329/A vssd1 vssd1 vccd1 vccd1 _5434_/CLK sky130_fd_sc_hd__inv_2
X_2972_ _5173_/Q _5237_/Q _3005_/S vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5691_ _5691_/CLK _5691_/D vssd1 vssd1 vccd1 vccd1 _5691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold703 hold703/A vssd1 vssd1 vccd1 vccd1 _4204_/A sky130_fd_sc_hd__buf_2
X_3524_ _5139_/Q _3614_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5139_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4637__222 _4485__70/A vssd1 vssd1 vccd1 vccd1 _5315_/CLK sky130_fd_sc_hd__inv_2
XFILLER_143_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3455_ _3608_/A1 _5201_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5201_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold758 _3831_/Y vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__buf_2
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2126 hold2126/A vssd1 vssd1 vccd1 vccd1 hold493/A sky130_fd_sc_hd__buf_2
Xhold2104 hold463/X vssd1 vssd1 vccd1 vccd1 hold2104/X sky130_fd_sc_hd__buf_2
X_3386_ _5294_/Q _3578_/A0 _3387_/S vssd1 vssd1 vccd1 vccd1 _5294_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5125_ _5125_/CLK _5125_/D vssd1 vssd1 vccd1 vccd1 _5125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1403 hold2165/X vssd1 vssd1 vccd1 vccd1 hold2166/A sky130_fd_sc_hd__buf_2
Xhold2148 hold2148/A vssd1 vssd1 vccd1 vccd1 hold542/A sky130_fd_sc_hd__buf_2
Xhold2137 hold2137/A vssd1 vssd1 vccd1 vccd1 _3875_/B1 sky130_fd_sc_hd__buf_2
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1414 hold2069/X vssd1 vssd1 vccd1 vccd1 hold2070/A sky130_fd_sc_hd__buf_2
X_5056_ _5056_/CLK _5056_/D vssd1 vssd1 vccd1 vccd1 _5056_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1447 hold1455/X vssd1 vssd1 vccd1 vccd1 hold1456/A sky130_fd_sc_hd__buf_2
X_4007_ _5670_/Q _5669_/Q vssd1 vssd1 vccd1 vccd1 _4008_/B sky130_fd_sc_hd__and2_2
Xhold1469 hold2244/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__buf_2
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5889_ _5889_/A vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__buf_2
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__buf_2
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__buf_2
Xhold2671 hold2671/A vssd1 vssd1 vccd1 vccd1 hold2671/X sky130_fd_sc_hd__buf_2
Xhold2682 hold265/X vssd1 vssd1 vccd1 vccd1 hold2682/X sky130_fd_sc_hd__buf_2
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__buf_2
Xhold63 hold84/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__buf_2
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__buf_2
XFILLER_29_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__buf_2
Xhold1992 hold2625/X vssd1 vssd1 vccd1 vccd1 hold2626/A sky130_fd_sc_hd__buf_2
XFILLER_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_85_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4457__42/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_14_wb_clk_i _4676__261/A vssd1 vssd1 vccd1 vccd1 _4693__278/A sky130_fd_sc_hd__clkbuf_16
XFILLER_77_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 _3692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3219_/X _3220_/X _3240_/S vssd1 vssd1 vccd1 vccd1 _3240_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3171_/A _3171_/B vssd1 vssd1 vccd1 vccd1 _3171_/X sky130_fd_sc_hd__and2_1
XFILLER_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4500__85 _4508__93/A vssd1 vssd1 vccd1 vccd1 _5142_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5743_ _5743_/CLK _5743_/D vssd1 vssd1 vccd1 vccd1 _5743_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2955_ _3593_/A1 _2895_/Y _2954_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5379_/D sky130_fd_sc_hd__o211a_1
X_2886_ _5065_/Q _5041_/Q _5538_/Q _4982_/Q _2941_/S0 _3024_/S vssd1 vssd1 vccd1 vccd1
+ _2886_/X sky130_fd_sc_hd__mux4_1
X_5674_ _5677_/CLK _5674_/D vssd1 vssd1 vccd1 vccd1 _5674_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold500 hold500/A vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__buf_2
X_3507_ _5154_/Q _3543_/A0 _3507_/S vssd1 vssd1 vccd1 vccd1 _5154_/D sky130_fd_sc_hd__mux2_1
Xhold522 hold522/A vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__buf_2
X_4871__456 _4875__460/A vssd1 vssd1 vccd1 vccd1 _5592_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold555 _3894_/X vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__buf_2
Xhold577 hold577/A vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__buf_2
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3438_ _5222_/Q _3593_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5222_/D sky130_fd_sc_hd__mux2_1
Xhold599 hold599/A vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__buf_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3369_ _3543_/A0 _5310_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5310_/D sky130_fd_sc_hd__mux2_1
Xhold1200 hold1910/X vssd1 vssd1 vccd1 vccd1 hold1911/A sky130_fd_sc_hd__buf_2
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912__497 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5633_/CLK sky130_fd_sc_hd__inv_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5256_/CLK _5108_/D vssd1 vssd1 vccd1 vccd1 _5108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1211 hold1915/X vssd1 vssd1 vccd1 vccd1 hold1916/A sky130_fd_sc_hd__buf_2
XFILLER_58_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1233 hold1939/X vssd1 vssd1 vccd1 vccd1 hold1940/A sky130_fd_sc_hd__buf_2
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1255 hold2476/X vssd1 vssd1 vccd1 vccd1 hold2477/A sky130_fd_sc_hd__buf_2
XFILLER_85_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4765__350 _5106_/CLK vssd1 vssd1 vccd1 vccd1 _5456_/CLK sky130_fd_sc_hd__inv_2
X_5039_ _5039_/CLK _5039_/D vssd1 vssd1 vccd1 vccd1 _5039_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1299 hold2588/X vssd1 vssd1 vccd1 vccd1 hold1857/A sky130_fd_sc_hd__buf_2
XFILLER_122_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4806__391 _4897__482/A vssd1 vssd1 vccd1 vccd1 _5497_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput120 probe_out[86] vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput131 probe_out[96] vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput142 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _2497_/B sky130_fd_sc_hd__clkbuf_2
Xinput153 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _2494_/B sky130_fd_sc_hd__clkbuf_2
Xhold2490 hold2490/A vssd1 vssd1 vccd1 vccd1 hold2490/X sky130_fd_sc_hd__buf_2
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput164 input164/A vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__buf_4
Xinput175 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _3645_/A sky130_fd_sc_hd__clkbuf_8
Xinput186 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _3655_/A sky130_fd_sc_hd__buf_4
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput197 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__buf_6
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _3571_/A _2740_/B vssd1 vssd1 vccd1 vccd1 _2748_/S sky130_fd_sc_hd__or2_4
XFILLER_145_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2671_ _5576_/Q _3569_/A1 _2672_/S vssd1 vssd1 vccd1 vccd1 _5576_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4410_ _4410_/A1 _4401_/Y _4409_/X _4368_/A vssd1 vssd1 vccd1 vccd1 _4410_/X sky130_fd_sc_hd__o211a_1
X_5390_ _5390_/CLK _5390_/D vssd1 vssd1 vccd1 vccd1 _5390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4341_ _5688_/Q _4324_/X _4340_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5687_/D sky130_fd_sc_hd__o211a_1
XFILLER_141_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4272_ _5743_/Q _4266_/B _4042_/A _4271_/Y vssd1 vssd1 vccd1 vccd1 _4277_/B sky130_fd_sc_hd__a211o_1
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3223_ _5642_/Q _3326_/B2 _3320_/C1 _3222_/X vssd1 vssd1 vccd1 vccd1 _3223_/X sky130_fd_sc_hd__o211a_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4749__334 _5010_/CLK vssd1 vssd1 vccd1 vccd1 _5440_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3154_ _3323_/C1 _3147_/X _3153_/X vssd1 vssd1 vccd1 vccd1 _3154_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3085_ _2777_/A _3081_/B _3535_/B _3083_/X _2778_/A vssd1 vssd1 vccd1 vccd1 _5373_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3987_ _3651_/A _5256_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _5256_/D sky130_fd_sc_hd__mux2_1
X_2938_ _5142_/Q _5150_/Q _5214_/Q _5134_/Q _3036_/S _2943_/S1 vssd1 vssd1 vccd1 vccd1
+ _2938_/X sky130_fd_sc_hd__mux4_2
X_5726_ _5726_/CLK _5726_/D vssd1 vssd1 vccd1 vccd1 _5726_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2869_ _2873_/B _2870_/B vssd1 vssd1 vccd1 vccd1 _2869_/Y sky130_fd_sc_hd__nor2_1
X_5657_ _5657_/CLK _5657_/D vssd1 vssd1 vccd1 vccd1 _5657_/Q sky130_fd_sc_hd__dfxtp_1
X_5588_ _5588_/CLK _5588_/D vssd1 vssd1 vccd1 vccd1 _5588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold352 hold352/A vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__buf_2
XFILLER_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold374 hold379/X vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__buf_2
Xhold363 hold371/X vssd1 vssd1 vccd1 vccd1 hold372/A sky130_fd_sc_hd__buf_2
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1030 hold1614/X vssd1 vssd1 vccd1 vccd1 hold1615/A sky130_fd_sc_hd__buf_2
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1041 hold1858/X vssd1 vssd1 vccd1 vccd1 hold1859/A sky130_fd_sc_hd__buf_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1074 hold1834/X vssd1 vssd1 vccd1 vccd1 hold1835/A sky130_fd_sc_hd__buf_2
Xhold1052 hold1838/X vssd1 vssd1 vccd1 vccd1 hold1839/A sky130_fd_sc_hd__buf_2
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1085 hold2304/X vssd1 vssd1 vccd1 vccd1 hold2305/A sky130_fd_sc_hd__buf_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4491__76 _4504__89/A vssd1 vssd1 vccd1 vccd1 _5133_/CLK sky130_fd_sc_hd__inv_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4542__127 _4421__6/A vssd1 vssd1 vccd1 vccd1 _5184_/CLK sky130_fd_sc_hd__inv_2
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3910_ _5742_/Q _3924_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3910_/X sky130_fd_sc_hd__and3_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3841_ _3844_/A _3955_/A vssd1 vssd1 vccd1 vccd1 _3959_/B sky130_fd_sc_hd__nor2_2
X_3772_ _5013_/Q _3774_/A2 _3774_/B1 _3771_/X _3774_/C1 vssd1 vssd1 vccd1 vccd1 _3772_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5511_ _5511_/CLK _5511_/D vssd1 vssd1 vccd1 vccd1 _5511_/Q sky130_fd_sc_hd__dfxtp_1
X_2723_ _3159_/A _5504_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5504_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2654_ _5370_/Q _2776_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _3589_/A sky130_fd_sc_hd__or3_4
Xoutput402 _3712_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__clkbuf_2
X_5442_ _5442_/CLK _5442_/D vssd1 vssd1 vccd1 vccd1 _5442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5373_ _5373_/CLK _5373_/D vssd1 vssd1 vccd1 vccd1 _5373_/Q sky130_fd_sc_hd__dfxtp_4
X_2585_ _5335_/Q _5334_/Q _3346_/A vssd1 vssd1 vccd1 vccd1 _3388_/B sky130_fd_sc_hd__or3_4
XFILLER_141_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4324_ _4324_/A _4324_/B _4074_/D vssd1 vssd1 vccd1 vccd1 _4324_/X sky130_fd_sc_hd__or3b_4
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _4254_/B _4254_/C _5749_/Q vssd1 vssd1 vccd1 vccd1 _4255_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4186_ _4186_/A _4186_/B vssd1 vssd1 vccd1 vccd1 _4186_/X sky130_fd_sc_hd__or2_2
X_3206_ _3323_/C1 _3205_/X _3353_/B vssd1 vssd1 vccd1 vccd1 _3206_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3137_ _5630_/Q _5520_/Q _5289_/Q _5472_/Q _3219_/S0 _3330_/S vssd1 vssd1 vccd1 vccd1
+ _3137_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3068_ _3099_/B _3066_/X _3067_/X vssd1 vssd1 vccd1 vccd1 _3068_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4877__462 _4901__486/A vssd1 vssd1 vccd1 vccd1 _5598_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5709_ _5709_/CLK _5709_/D vssd1 vssd1 vccd1 vccd1 _5709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold160 _3971_/Y vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__buf_2
XFILLER_2_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold171 _3626_/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__buf_2
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__buf_2
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__buf_2
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout640 _3732_/B vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__buf_6
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4670__255 _5006_/CLK vssd1 vssd1 vccd1 vccd1 _5358_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_4040_ _4052_/B _4052_/C _5747_/Q vssd1 vssd1 vccd1 vccd1 _4042_/B sky130_fd_sc_hd__o21a_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4711__296 _5106_/CLK vssd1 vssd1 vccd1 vccd1 _5402_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3824_ _3824_/A1 _3930_/A split4/A _5023_/Q vssd1 vssd1 vccd1 vccd1 _3824_/X sky130_fd_sc_hd__a31o_1
X_3755_ _3755_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__and2_1
X_4605__190 _5683_/CLK vssd1 vssd1 vccd1 vccd1 _5279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3686_ _5259_/Q _3688_/B vssd1 vssd1 vccd1 vccd1 _3686_/X sky130_fd_sc_hd__and2_1
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2706_ _3391_/A0 _5518_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5518_/D sky130_fd_sc_hd__mux2_1
Xoutput210 _3673_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__clkbuf_2
X_2637_ _5606_/Q _3599_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5606_/D sky130_fd_sc_hd__mux2_1
X_5425_ _5425_/CLK _5425_/D vssd1 vssd1 vccd1 vccd1 _5425_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput221 _3683_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput243 _3645_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__clkbuf_2
Xoutput232 _3668_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput254 _3655_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__clkbuf_2
Xoutput265 _3636_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5356_ _5356_/CLK _5356_/D vssd1 vssd1 vccd1 vccd1 _5356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2568_ _3573_/A0 _5645_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5645_/D sky130_fd_sc_hd__mux2_1
Xoutput276 _5848_/X vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_12
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4307_ _4306_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5673_/D sky130_fd_sc_hd__and2b_1
X_2499_ _4353_/A _3959_/A split5/A vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__and3_4
X_5287_ _5287_/CLK _5287_/D vssd1 vssd1 vccd1 vccd1 _5287_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput287 _5858_/X vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_12
Xoutput298 _5868_/X vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_12
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4238_ _5563_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__or2_1
XFILLER_101_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4169_ _4169_/A _4169_/B _4169_/C _4169_/D vssd1 vssd1 vccd1 vccd1 _4170_/D sky130_fd_sc_hd__and4_1
XFILLER_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4461__46 _5683_/CLK vssd1 vssd1 vccd1 vccd1 _5055_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4654__239 _5726_/CLK vssd1 vssd1 vccd1 vccd1 _5340_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4424__9/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout492 hold364/X vssd1 vssd1 vccd1 vccd1 _3814_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout481 _3074_/A1 vssd1 vssd1 vccd1 vccd1 _3099_/B sky130_fd_sc_hd__buf_6
XFILLER_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout470 _3357_/B vssd1 vssd1 vccd1 vccd1 _3325_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4548__133 _4423__8/A vssd1 vssd1 vccd1 vccd1 _5190_/CLK sky130_fd_sc_hd__inv_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _3603_/A1 _5125_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5125_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3471_ _5186_/Q _3615_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5186_/D sky130_fd_sc_hd__mux2_1
X_5210_ _5210_/CLK _5210_/D vssd1 vssd1 vccd1 vccd1 _5210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold929 hold929/A vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__buf_2
XFILLER_115_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5141_ _5141_/CLK _5141_/D vssd1 vssd1 vccd1 vccd1 _5141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2308 hold2308/A vssd1 vssd1 vccd1 vccd1 hold2308/X sky130_fd_sc_hd__buf_2
Xhold2319 hold2319/A vssd1 vssd1 vccd1 vccd1 hold723/A sky130_fd_sc_hd__buf_2
Xhold1607 hold1607/A vssd1 vssd1 vccd1 vccd1 _5101_/D sky130_fd_sc_hd__buf_2
X_5072_ _5752_/CLK _5072_/D vssd1 vssd1 vccd1 vccd1 _5072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1629 hold2204/X vssd1 vssd1 vccd1 vccd1 hold2205/A sky130_fd_sc_hd__buf_2
Xhold1618 hold50/X vssd1 vssd1 vccd1 vccd1 hold1618/X sky130_fd_sc_hd__buf_2
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4023_ _5744_/Q _4023_/B vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__xnor2_1
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3807_ _5258_/Q hold277/X _3814_/A3 _3814_/B1 _5007_/Q vssd1 vssd1 vccd1 vccd1 _3807_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_107_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3738_ _4999_/Q _3750_/B vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__or2_1
X_3669_ _3669_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__and2_1
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5408_ _5408_/CLK _5408_/D vssd1 vssd1 vccd1 vccd1 _5408_/Q sky130_fd_sc_hd__dfxtp_1
X_4506__91 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5148_/CLK sky130_fd_sc_hd__inv_2
X_5339_ _5339_/CLK _5339_/D vssd1 vssd1 vccd1 vccd1 _5339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2831 _4094_/X vssd1 vssd1 vccd1 vccd1 hold2831/X sky130_fd_sc_hd__buf_2
Xhold2820 hold2820/A vssd1 vssd1 vccd1 vccd1 hold2820/X sky130_fd_sc_hd__buf_2
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2875 _4416_/X vssd1 vssd1 vccd1 vccd1 hold2875/X sky130_fd_sc_hd__buf_2
XFILLER_18_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2897 hold2903/X vssd1 vssd1 vccd1 vccd1 hold2904/A sky130_fd_sc_hd__buf_2
Xhold2886 hold2886/A vssd1 vssd1 vccd1 vccd1 hold2886/X sky130_fd_sc_hd__buf_2
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4782__367 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5473_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2971_ _5221_/Q _2873_/B _2870_/B vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__a21o_1
X_5690_ _5691_/CLK _5690_/D vssd1 vssd1 vccd1 vccd1 _5690_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3523_ _5140_/Q _3613_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5140_/D sky130_fd_sc_hd__mux2_1
X_4676__261 _4676__261/A vssd1 vssd1 vccd1 vccd1 _5365_/CLK sky130_fd_sc_hd__inv_2
Xhold704 _4192_/Y vssd1 vssd1 vccd1 vccd1 _5542_/D sky130_fd_sc_hd__buf_2
XFILLER_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3454_ _3589_/A _3607_/B vssd1 vssd1 vccd1 vccd1 _3462_/S sky130_fd_sc_hd__or2_4
XFILLER_116_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold759 hold759/A vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__buf_2
Xhold748 hold748/A vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__buf_2
XFILLER_143_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2116 _3869_/X vssd1 vssd1 vccd1 vccd1 hold2116/X sky130_fd_sc_hd__buf_2
Xhold2127 hold493/X vssd1 vssd1 vccd1 vccd1 hold2127/X sky130_fd_sc_hd__buf_2
X_3385_ _5295_/Q _3568_/A1 _3387_/S vssd1 vssd1 vccd1 vccd1 _5295_/D sky130_fd_sc_hd__mux2_1
Xhold2105 hold2105/A vssd1 vssd1 vccd1 vccd1 _4983_/D sky130_fd_sc_hd__buf_2
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5124_ _5124_/CLK _5124_/D vssd1 vssd1 vccd1 vccd1 _5124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1404 hold2167/X vssd1 vssd1 vccd1 vccd1 hold2168/A sky130_fd_sc_hd__buf_2
Xhold2138 _3875_/X vssd1 vssd1 vccd1 vccd1 hold2138/X sky130_fd_sc_hd__buf_2
XFILLER_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5055_ _5055_/CLK _5055_/D vssd1 vssd1 vccd1 vccd1 _5055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1448 hold452/X vssd1 vssd1 vccd1 vccd1 hold415/A sky130_fd_sc_hd__buf_2
Xhold1459 hold1459/A vssd1 vssd1 vccd1 vccd1 hold1459/X sky130_fd_sc_hd__buf_2
X_4006_ _5668_/Q _5667_/Q _5666_/Q _5665_/Q vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__nand4_4
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4431__16 _4469__54/A vssd1 vssd1 vccd1 vccd1 _4982_/CLK sky130_fd_sc_hd__inv_2
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5888_ _5888_/A vssd1 vssd1 vccd1 vccd1 _5888_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4917__502 _4455__40/A vssd1 vssd1 vccd1 vccd1 _5638_/CLK sky130_fd_sc_hd__inv_2
XFILLER_147_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__buf_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__buf_2
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__buf_2
XFILLER_76_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__buf_2
Xhold2683 hold2683/A vssd1 vssd1 vccd1 vccd1 hold2683/X sky130_fd_sc_hd__buf_2
Xhold64 hold86/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__buf_2
Xhold2672 hold2672/A vssd1 vssd1 vccd1 vccd1 hold2672/X sky130_fd_sc_hd__buf_2
XFILLER_91_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1960 hold2047/X vssd1 vssd1 vccd1 vccd1 hold2048/A sky130_fd_sc_hd__buf_2
Xhold2694 _3796_/X vssd1 vssd1 vccd1 vccd1 hold2694/X sky130_fd_sc_hd__buf_2
Xhold86 hold9/X vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__buf_2
XFILLER_29_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__buf_2
Xhold1993 hold2627/X vssd1 vssd1 vccd1 vccd1 hold2628/A sky130_fd_sc_hd__buf_2
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 _5319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5106_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3170_ _5714_/Q _5463_/Q _5447_/Q _5479_/Q _3330_/S _3219_/S0 vssd1 vssd1 vccd1 vccd1
+ _3171_/B sky130_fd_sc_hd__mux4_1
X_4497__82 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5139_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5742_ _5742_/CLK _5742_/D vssd1 vssd1 vccd1 vccd1 _5742_/Q sky130_fd_sc_hd__dfxtp_4
X_2954_ _2863_/A _5379_/Q _3094_/A _2953_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _2954_/X
+ sky130_fd_sc_hd__a221o_1
X_2885_ _5590_/Q _5574_/Q _5456_/Q _5606_/Q _3024_/S _2941_/S0 vssd1 vssd1 vccd1 vccd1
+ _2885_/X sky130_fd_sc_hd__mux4_2
X_5673_ _5725_/CLK _5673_/D vssd1 vssd1 vccd1 vccd1 _5673_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold501 hold501/A vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__buf_2
X_3506_ _5155_/Q _3605_/A1 _3507_/S vssd1 vssd1 vccd1 vccd1 _5155_/D sky130_fd_sc_hd__mux2_1
Xhold534 hold577/X vssd1 vssd1 vccd1 vccd1 hold578/A sky130_fd_sc_hd__buf_2
Xhold512 hold512/A vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__buf_2
XFILLER_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold556 _3895_/X vssd1 vssd1 vccd1 vccd1 _5073_/D sky130_fd_sc_hd__buf_2
Xhold578 hold578/A vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__buf_2
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold589 hold589/A vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__buf_2
X_3437_ _5223_/Q _3592_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5223_/D sky130_fd_sc_hd__mux2_1
X_3368_ _3605_/A1 _5311_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5311_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5256_/CLK _5107_/D vssd1 vssd1 vccd1 vccd1 _5107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1212 hold1917/X vssd1 vssd1 vccd1 vccd1 hold1918/A sky130_fd_sc_hd__buf_2
Xhold1234 hold1941/X vssd1 vssd1 vccd1 vccd1 hold1942/A sky130_fd_sc_hd__buf_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3299_ _5442_/Q _5458_/Q _3299_/S vssd1 vssd1 vccd1 vccd1 _3299_/X sky130_fd_sc_hd__mux2_2
X_5038_ _5038_/CLK _5038_/D vssd1 vssd1 vccd1 vccd1 _5038_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1289 hold2537/X vssd1 vssd1 vccd1 vccd1 hold2538/A sky130_fd_sc_hd__buf_2
XFILLER_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput110 probe_out[77] vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput132 probe_out[97] vssd1 vssd1 vccd1 vccd1 _5934_/A sky130_fd_sc_hd__clkbuf_2
Xinput121 probe_out[87] vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput143 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _2497_/A sky130_fd_sc_hd__clkbuf_2
Xinput154 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _2494_/A sky130_fd_sc_hd__clkbuf_2
Xhold2491 hold2491/A vssd1 vssd1 vccd1 vccd1 _5319_/D sky130_fd_sc_hd__buf_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput165 input165/A vssd1 vssd1 vccd1 vccd1 _3669_/A sky130_fd_sc_hd__buf_4
Xinput176 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__clkbuf_8
Xinput187 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__buf_4
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput198 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _3637_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1790 hold2525/X vssd1 vssd1 vccd1 vccd1 hold2526/A sky130_fd_sc_hd__buf_2
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_101_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4658__243/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2670_ _5577_/Q _3577_/A0 _2672_/S vssd1 vssd1 vccd1 vccd1 _5577_/D sky130_fd_sc_hd__mux2_1
X_4894__479 _4897__482/A vssd1 vssd1 vccd1 vccd1 _5615_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4340_ _5687_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4340_/X sky130_fd_sc_hd__or2_1
XFILLER_140_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4271_ _4271_/A _4271_/B _4271_/C _4271_/D vssd1 vssd1 vccd1 vccd1 _4271_/Y sky130_fd_sc_hd__nand4_1
XFILLER_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3222_ _5650_/Q _3132_/A _3221_/X _3325_/A vssd1 vssd1 vccd1 vccd1 _3222_/X sky130_fd_sc_hd__o22a_1
XFILLER_95_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3153_ _3316_/C1 _3146_/X _3353_/B vssd1 vssd1 vccd1 vccd1 _3153_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4788__373 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5479_/CLK sky130_fd_sc_hd__inv_2
X_3084_ _5373_/Q _3443_/B _3453_/C vssd1 vssd1 vccd1 vccd1 _3535_/B sky130_fd_sc_hd__nand3_4
XFILLER_63_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3986_ _3650_/A _5255_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _5255_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2937_ _5118_/Q _5166_/Q _5351_/Q _5230_/Q _2944_/S0 _3066_/S vssd1 vssd1 vccd1 vccd1
+ _2937_/X sky130_fd_sc_hd__mux4_1
X_5725_ _5725_/CLK _5725_/D vssd1 vssd1 vccd1 vccd1 _5725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _5656_/CLK _5656_/D vssd1 vssd1 vccd1 vccd1 _5656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2868_ _2941_/S0 _3072_/S _5366_/Q vssd1 vssd1 vccd1 vccd1 _2868_/Y sky130_fd_sc_hd__a21oi_2
X_5587_ _5587_/CLK _5587_/D vssd1 vssd1 vccd1 vccd1 _5587_/Q sky130_fd_sc_hd__dfxtp_1
X_2799_ _5440_/Q _3536_/A0 _2806_/S vssd1 vssd1 vccd1 vccd1 _5440_/D sky130_fd_sc_hd__mux2_1
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__buf_2
XFILLER_117_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold353 hold353/A vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__buf_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold364 hold364/A vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__buf_2
Xhold386 hold399/X vssd1 vssd1 vccd1 vccd1 hold400/A sky130_fd_sc_hd__buf_2
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1020 hold1606/X vssd1 vssd1 vccd1 vccd1 hold1607/A sky130_fd_sc_hd__buf_2
Xhold1031 hold1616/X vssd1 vssd1 vccd1 vccd1 hold1617/A sky130_fd_sc_hd__buf_2
Xhold1042 hold1860/X vssd1 vssd1 vccd1 vccd1 hold1861/A sky130_fd_sc_hd__buf_2
XFILLER_18_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1075 hold1864/X vssd1 vssd1 vccd1 vccd1 hold1865/A sky130_fd_sc_hd__buf_2
XFILLER_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1086 hold2308/X vssd1 vssd1 vccd1 vccd1 hold2309/A sky130_fd_sc_hd__buf_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4581__166 _4477__62/A vssd1 vssd1 vccd1 vccd1 _5231_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4467__52 _4469__54/A vssd1 vssd1 vccd1 vccd1 _5061_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4822__407 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5513_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3840_ _5530_/Q _3839_/X _4186_/A _4204_/A vssd1 vssd1 vccd1 vccd1 _5025_/D sky130_fd_sc_hd__a211o_4
X_3771_ _3771_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3771_/X sky130_fd_sc_hd__and2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5510_ _5510_/CLK _5510_/D vssd1 vssd1 vccd1 vccd1 _5510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2722_ _3562_/A _2740_/B vssd1 vssd1 vccd1 vccd1 _2730_/S sky130_fd_sc_hd__or2_4
XFILLER_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2653_ _5591_/Q _3387_/A1 _2653_/S vssd1 vssd1 vccd1 vccd1 _5591_/D sky130_fd_sc_hd__mux2_1
X_5441_ _5441_/CLK _5441_/D vssd1 vssd1 vccd1 vccd1 _5441_/Q sky130_fd_sc_hd__dfxtp_1
X_4716__301 _5261_/CLK vssd1 vssd1 vccd1 vccd1 _5407_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5372_ _5372_/CLK _5372_/D vssd1 vssd1 vccd1 vccd1 _5372_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput403 _3715_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__clkbuf_2
X_2584_ _3387_/A1 _5631_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5631_/D sky130_fd_sc_hd__mux2_4
X_4323_ _4320_/X _4322_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4254_ _5749_/Q _4254_/B _4254_/C vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__and3_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3205_ _5720_/Q _5297_/Q _5270_/Q _5704_/Q _3290_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3205_/X sky130_fd_sc_hd__mux4_1
X_4185_ _4187_/B1 _4183_/Y _4184_/Y _5539_/Q _4244_/S vssd1 vssd1 vccd1 vccd1 _5539_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3136_ _5330_/Q _3140_/A vssd1 vssd1 vccd1 vccd1 _3136_/X sky130_fd_sc_hd__xor2_4
X_3067_ _5218_/Q _2866_/A _2866_/B _5026_/Q _2945_/A vssd1 vssd1 vccd1 vccd1 _3067_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_82_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ _5381_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _5208_/D sky130_fd_sc_hd__and2_1
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5708_ _5708_/CLK _5708_/D vssd1 vssd1 vccd1 vccd1 _5708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5639_ _5639_/CLK _5639_/D vssd1 vssd1 vccd1 vccd1 _5639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__buf_2
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 _3979_/S sky130_fd_sc_hd__buf_2
XFILLER_144_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__buf_2
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__buf_2
Xhold183 _3729_/B vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__buf_2
XFILLER_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout641 _3732_/B vssd1 vssd1 vccd1 vccd1 _3774_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout630 _5112_/Q vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__buf_6
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3823_ _4357_/A _5022_/Q hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__mux2_1
XFILLER_20_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3754_ _5004_/Q _3750_/B _3752_/X _3774_/B1 _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3754_/X
+ sky130_fd_sc_hd__o221a_4
Xclkbuf_leaf_9_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5751_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3685_ _5258_/Q _3688_/B vssd1 vssd1 vccd1 vccd1 _3685_/X sky130_fd_sc_hd__and2_1
X_2705_ _3390_/A0 _5519_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5519_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2636_ _2779_/A _3526_/A vssd1 vssd1 vccd1 vccd1 _2644_/S sky130_fd_sc_hd__nor2_8
X_5424_ _5424_/CLK _5424_/D vssd1 vssd1 vccd1 vccd1 _5424_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput222 _3684_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__clkbuf_2
Xoutput244 _3646_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__clkbuf_2
Xoutput233 _3669_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput211 _3674_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950__535 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5708_/CLK sky130_fd_sc_hd__inv_2
Xoutput255 _3656_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput266 _3637_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__clkbuf_2
X_5355_ _5355_/CLK _5355_/D vssd1 vssd1 vccd1 vccd1 _5355_/Q sky130_fd_sc_hd__dfxtp_1
X_2567_ _3159_/A _5646_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5646_/D sky130_fd_sc_hd__mux2_1
Xoutput277 _5849_/X vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_12
XFILLER_114_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4306_ _4039_/X _4308_/A2 _4308_/B1 _2445_/Y vssd1 vssd1 vccd1 vccd1 _4306_/X sky130_fd_sc_hd__o22a_1
X_2498_ _3711_/B split4/A vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__and2_4
X_5286_ _5286_/CLK _5286_/D vssd1 vssd1 vccd1 vccd1 _5286_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput288 _5859_/X vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_12
Xoutput299 _5869_/X vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_12
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4237_ _5341_/Q _4360_/B _4164_/B _4236_/X _4244_/S vssd1 vssd1 vccd1 vccd1 _5562_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4122_/X _4123_/Y _4157_/B _5746_/Q _4118_/C vssd1 vssd1 vccd1 vccd1 _4170_/C
+ sky130_fd_sc_hd__o221a_1
X_3119_ _3595_/A1 _5349_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5349_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4099_ _5542_/Q _5541_/Q _5540_/Q _5539_/Q vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__and4_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4693__278 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5382_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout482 _3074_/A1 vssd1 vssd1 vccd1 vccd1 _3034_/A sky130_fd_sc_hd__buf_6
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout471 _3301_/A1 vssd1 vssd1 vccd1 vccd1 _3357_/B sky130_fd_sc_hd__buf_6
Xfanout493 _3298_/B1 vssd1 vssd1 vccd1 vccd1 _3237_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_101_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4437__22 _5111_/CLK vssd1 vssd1 vccd1 vccd1 _5031_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_79_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4463__48/A sky130_fd_sc_hd__clkbuf_16
XFILLER_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4587__172 _4435__20/A vssd1 vssd1 vccd1 vccd1 _5237_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4934__519 _5244_/CLK vssd1 vssd1 vccd1 vccd1 _5655_/CLK sky130_fd_sc_hd__inv_2
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3470_ _5187_/Q _3614_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5187_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5140_ _5140_/CLK _5140_/D vssd1 vssd1 vccd1 vccd1 _5140_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2309 hold2309/A vssd1 vssd1 vccd1 vccd1 hold2309/X sky130_fd_sc_hd__buf_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5071_ _5755_/CLK _5071_/D vssd1 vssd1 vccd1 vccd1 _5071_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1608 hold2448/X vssd1 vssd1 vccd1 vccd1 hold2449/A sky130_fd_sc_hd__buf_2
Xhold1619 hold1619/A vssd1 vssd1 vccd1 vccd1 _5100_/D sky130_fd_sc_hd__buf_2
X_4022_ _2442_/Y _4071_/B _4027_/B vssd1 vssd1 vccd1 vccd1 _4023_/B sky130_fd_sc_hd__a21bo_2
X_4828__413 _5022_/CLK vssd1 vssd1 vccd1 vccd1 _5519_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3806_ hold277/X _5257_/Q _3814_/A3 _3814_/B1 _5006_/Q vssd1 vssd1 vccd1 vccd1 _3806_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3737_ _5082_/Q input10/X _3763_/B vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3668_ _3668_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__and2_1
XFILLER_134_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5407_ _5407_/CLK _5407_/D vssd1 vssd1 vccd1 vccd1 _5407_/Q sky130_fd_sc_hd__dfxtp_1
X_3599_ _4982_/Q _3599_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4982_/D sky130_fd_sc_hd__mux2_1
X_2619_ _3453_/C _2867_/A vssd1 vssd1 vccd1 vccd1 _2861_/A sky130_fd_sc_hd__xor2_4
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5338_ _5338_/CLK _5338_/D vssd1 vssd1 vccd1 vccd1 _5338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2832 hold2832/A vssd1 vssd1 vccd1 vccd1 hold2832/X sky130_fd_sc_hd__buf_2
Xhold2821 hold2821/A vssd1 vssd1 vccd1 vccd1 hold2821/X sky130_fd_sc_hd__buf_2
XFILLER_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5269_ _5269_/CLK _5269_/D vssd1 vssd1 vccd1 vccd1 _5269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2898 hold2905/X vssd1 vssd1 vccd1 vccd1 hold2906/A sky130_fd_sc_hd__buf_2
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2887 hold2887/A vssd1 vssd1 vccd1 vccd1 hold2887/X sky130_fd_sc_hd__buf_2
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4621__206 _4964__549/A vssd1 vssd1 vccd1 vccd1 _5298_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4515__100 _5684_/CLK vssd1 vssd1 vccd1 vccd1 _5157_/CLK sky130_fd_sc_hd__inv_2
XFILLER_120_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2970_ _3041_/B1 _2968_/X _2969_/X vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3522_ _5141_/Q _3612_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5141_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold727 hold727/A vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__buf_2
X_3453_ _5373_/Q _5372_/Q _3453_/C vssd1 vssd1 vccd1 vccd1 _3607_/B sky130_fd_sc_hd__nand3b_4
Xhold738 hold758/X vssd1 vssd1 vccd1 vccd1 hold759/A sky130_fd_sc_hd__buf_2
XFILLER_131_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5123_ _5123_/CLK _5123_/D vssd1 vssd1 vccd1 vccd1 _5123_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2117 hold2117/A vssd1 vssd1 vccd1 vccd1 hold488/A sky130_fd_sc_hd__buf_2
X_3384_ _5296_/Q _3576_/A0 _3387_/S vssd1 vssd1 vccd1 vccd1 _5296_/D sky130_fd_sc_hd__mux2_1
Xhold1405 hold954/X vssd1 vssd1 vccd1 vccd1 _5384_/D sky130_fd_sc_hd__buf_2
Xhold2128 hold2128/A vssd1 vssd1 vccd1 vccd1 _3865_/B1 sky130_fd_sc_hd__buf_2
Xhold2139 hold2139/A vssd1 vssd1 vccd1 vccd1 hold522/A sky130_fd_sc_hd__buf_2
X_5054_ _5054_/CLK _5054_/D vssd1 vssd1 vccd1 vccd1 _5054_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1449 hold415/X vssd1 vssd1 vccd1 vccd1 hold453/A sky130_fd_sc_hd__buf_2
Xhold1438 hold2102/X vssd1 vssd1 vccd1 vccd1 hold2103/A sky130_fd_sc_hd__buf_2
X_4005_ _5668_/Q _5667_/Q _5666_/Q _5665_/Q vssd1 vssd1 vccd1 vccd1 _4021_/C sky130_fd_sc_hd__and4_4
XFILLER_38_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5887_ _5887_/A vssd1 vssd1 vccd1 vccd1 _5887_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956__541 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5714_/CLK sky130_fd_sc_hd__inv_2
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__buf_2
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__buf_2
XFILLER_29_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold10 hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__buf_2
XFILLER_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__buf_2
Xhold2673 hold2673/A vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__buf_2
Xhold2662 _3794_/X vssd1 vssd1 vccd1 vccd1 hold2662/X sky130_fd_sc_hd__buf_2
Xhold65 hold88/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__buf_2
Xhold54 hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__buf_2
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1950 hold803/X vssd1 vssd1 vccd1 vccd1 hold1950/X sky130_fd_sc_hd__buf_2
Xhold1961 hold2049/X vssd1 vssd1 vccd1 vccd1 _3957_/B sky130_fd_sc_hd__buf_2
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__buf_2
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__buf_2
Xhold2695 hold2695/A vssd1 vssd1 vccd1 vccd1 hold2695/X sky130_fd_sc_hd__buf_2
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__buf_2
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1994 hold2629/X vssd1 vssd1 vccd1 vccd1 hold2630/A sky130_fd_sc_hd__buf_2
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4699__284 _4731__316/A vssd1 vssd1 vccd1 vccd1 _5390_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 _5320_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_94_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4921__506/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4439__24/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _2883_/X _2950_/X _2952_/X _2948_/X vssd1 vssd1 vccd1 vccd1 _2953_/X sky130_fd_sc_hd__a31o_2
X_5741_ _5742_/CLK _5741_/D vssd1 vssd1 vccd1 vccd1 _5741_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2884_ _3043_/A _2877_/X _2881_/X _3094_/B vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__o211a_1
X_5672_ _5725_/CLK _5672_/D vssd1 vssd1 vccd1 vccd1 _5672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold502 hold502/A vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__buf_2
XFILLER_144_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3505_ _5156_/Q _3604_/A1 _3507_/S vssd1 vssd1 vccd1 vccd1 _5156_/D sky130_fd_sc_hd__mux2_1
Xhold535 hold553/X vssd1 vssd1 vccd1 vccd1 hold554/A sky130_fd_sc_hd__buf_2
XFILLER_144_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold579 hold579/A vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__buf_2
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3436_ _5224_/Q _3591_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5224_/D sky130_fd_sc_hd__mux2_1
X_3367_ _3604_/A1 _5312_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5312_/D sky130_fd_sc_hd__mux2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5106_/CLK _5106_/D vssd1 vssd1 vccd1 vccd1 _5106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1213 hold1919/X vssd1 vssd1 vccd1 vccd1 hold1920/A sky130_fd_sc_hd__buf_2
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ _5037_/CLK _5037_/D vssd1 vssd1 vccd1 vccd1 _5037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1235 hold1943/X vssd1 vssd1 vccd1 vccd1 hold1944/A sky130_fd_sc_hd__buf_2
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3298_ _5418_/Q _2482_/B _3298_/B1 _5410_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _3298_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_122_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1268 hold2498/X vssd1 vssd1 vccd1 vccd1 hold2499/A sky130_fd_sc_hd__buf_2
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4733__318 _4941__526/A vssd1 vssd1 vccd1 vccd1 _5424_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput111 probe_out[78] vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__clkbuf_2
Xinput100 probe_out[68] vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__clkbuf_2
Xinput122 probe_out[88] vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__clkbuf_2
Xinput133 probe_out[9] vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput144 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _2492_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput166 input166/A vssd1 vssd1 vccd1 vccd1 _3670_/A sky130_fd_sc_hd__buf_4
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput177 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__clkbuf_8
Xinput155 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__clkbuf_2
Xhold1780 hold2497/X vssd1 vssd1 vccd1 vccd1 hold2498/A sky130_fd_sc_hd__buf_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput199 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__clkbuf_8
Xinput188 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__buf_4
Xhold1791 hold2527/X vssd1 vssd1 vccd1 vccd1 hold2528/A sky130_fd_sc_hd__buf_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4627__212 _4459__44/A vssd1 vssd1 vccd1 vccd1 _5304_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4270_ _5742_/Q _4270_/B vssd1 vssd1 vccd1 vccd1 _4274_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3221_ _5045_/Q _5634_/Q _3284_/S vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3152_ _3316_/C1 _3142_/X _3151_/X vssd1 vssd1 vccd1 vccd1 _3152_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3083_ _5373_/Q _3087_/A vssd1 vssd1 vccd1 vccd1 _3083_/X sky130_fd_sc_hd__or2_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3985_ _3649_/A _5254_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _5254_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2936_ _3592_/A1 _2895_/Y _2935_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5380_/D sky130_fd_sc_hd__o211a_1
X_5724_ _5730_/CLK _5724_/D vssd1 vssd1 vccd1 vccd1 _5724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2867_ _2867_/A _2867_/B _3066_/S vssd1 vssd1 vccd1 vccd1 _2873_/B sky130_fd_sc_hd__and3_4
X_5655_ _5655_/CLK _5655_/D vssd1 vssd1 vccd1 vccd1 _5655_/Q sky130_fd_sc_hd__dfxtp_1
X_5586_ _5586_/CLK _5586_/D vssd1 vssd1 vccd1 vccd1 _5586_/Q sky130_fd_sc_hd__dfxtp_1
Xhold310 hold320/X vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__buf_2
X_2798_ _3598_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2806_/S sky130_fd_sc_hd__nor2_8
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 _3953_/S sky130_fd_sc_hd__buf_2
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold354 hold354/A vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__buf_2
Xhold365 _3811_/X vssd1 vssd1 vccd1 vccd1 _5011_/D sky130_fd_sc_hd__buf_2
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold387 hold403/X vssd1 vssd1 vccd1 vccd1 hold404/A sky130_fd_sc_hd__buf_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold398 hold408/X vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__buf_2
X_3419_ _3592_/A1 _5239_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5239_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4399_ _4399_/A _4399_/B _4399_/C _4399_/D vssd1 vssd1 vccd1 vccd1 _4409_/B sky130_fd_sc_hd__nor4_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1032 hold1618/X vssd1 vssd1 vccd1 vccd1 hold1619/A sky130_fd_sc_hd__buf_2
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1010 hold2434/X vssd1 vssd1 vccd1 vccd1 hold2435/A sky130_fd_sc_hd__buf_2
Xhold1021 hold2440/X vssd1 vssd1 vccd1 vccd1 hold2441/A sky130_fd_sc_hd__buf_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 hold2203/X vssd1 vssd1 vccd1 vccd1 hold2204/A sky130_fd_sc_hd__buf_2
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1043 hold1862/X vssd1 vssd1 vccd1 vccd1 hold1863/A sky130_fd_sc_hd__buf_2
Xhold1076 hold1866/X vssd1 vssd1 vccd1 vccd1 hold1867/A sky130_fd_sc_hd__buf_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4482__67 _5004_/CLK vssd1 vssd1 vccd1 vccd1 _5124_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4861__446 _4898__483/A vssd1 vssd1 vccd1 vccd1 _5582_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3770_ _5012_/Q _3774_/A2 _3774_/B1 _3769_/X _3774_/C1 vssd1 vssd1 vccd1 vccd1 _3770_/X
+ sky130_fd_sc_hd__o221a_4
X_4902__487 _5243_/CLK vssd1 vssd1 vccd1 vccd1 _5623_/CLK sky130_fd_sc_hd__inv_2
X_2721_ _3339_/A1 _5505_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5505_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5440_ _5440_/CLK _5440_/D vssd1 vssd1 vccd1 vccd1 _5440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2652_ _5592_/Q _3569_/A1 _2653_/S vssd1 vssd1 vccd1 vccd1 _5592_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5371_ _5371_/CLK _5371_/D vssd1 vssd1 vccd1 vccd1 _5371_/Q sky130_fd_sc_hd__dfxtp_2
X_4755__340 _5697_/CLK vssd1 vssd1 vccd1 vccd1 _5446_/CLK sky130_fd_sc_hd__inv_2
Xoutput404 _3718_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__clkbuf_2
X_2583_ _3578_/A0 _5632_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5632_/D sky130_fd_sc_hd__mux2_4
XFILLER_114_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ _4016_/B _4322_/B _4325_/B vssd1 vssd1 vccd1 vccd1 _4322_/X sky130_fd_sc_hd__and3b_1
XFILLER_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4253_ _4253_/A _4253_/B vssd1 vssd1 vccd1 vccd1 _4265_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3204_ _5054_/Q _5278_/Q _5525_/Q _5305_/Q _3324_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3204_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4184_ _4186_/B _4184_/B vssd1 vssd1 vccd1 vccd1 _4184_/Y sky130_fd_sc_hd__nor2_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3135_ _5330_/Q _3140_/A vssd1 vssd1 vccd1 vccd1 _3169_/B sky130_fd_sc_hd__xnor2_4
X_3066_ _5170_/Q _5234_/Q _3066_/S vssd1 vssd1 vccd1 vccd1 _3066_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3968_ _5380_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _5207_/D sky130_fd_sc_hd__and2_1
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2919_ _3099_/A _2919_/B vssd1 vssd1 vccd1 vccd1 _2919_/Y sky130_fd_sc_hd__nand2_1
X_5707_ _5707_/CLK _5707_/D vssd1 vssd1 vccd1 vccd1 _5707_/Q sky130_fd_sc_hd__dfxtp_1
X_3899_ _3844_/A _3955_/A _5074_/Q hold554/X vssd1 vssd1 vccd1 vccd1 _3899_/X sky130_fd_sc_hd__a31o_1
XFILLER_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5638_ _5638_/CLK _5638_/D vssd1 vssd1 vccd1 vccd1 _5638_/Q sky130_fd_sc_hd__dfxtp_1
X_5569_ _5569_/CLK _5569_/D vssd1 vssd1 vccd1 vccd1 _5569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__buf_2
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__buf_2
Xhold162 _3976_/X vssd1 vssd1 vccd1 vccd1 _5246_/D sky130_fd_sc_hd__buf_2
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__buf_2
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__buf_2
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__buf_2
XFILLER_144_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout620 _5319_/Q vssd1 vssd1 vccd1 vccd1 _3605_/A1 sky130_fd_sc_hd__buf_4
Xfanout631 _5111_/Q vssd1 vssd1 vccd1 vccd1 _3955_/A sky130_fd_sc_hd__buf_6
XFILLER_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout642 hold137/X vssd1 vssd1 vccd1 vccd1 _3782_/A sky130_fd_sc_hd__buf_12
XFILLER_144_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739__324 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5430_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3822_ _4356_/A _5021_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _5021_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3753_ _5087_/Q _3778_/C _3778_/B vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__a21bo_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3684_ _5257_/Q _3688_/B vssd1 vssd1 vccd1 vccd1 _3684_/X sky130_fd_sc_hd__and2_1
X_2704_ _3389_/A0 _5520_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5520_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2635_ _5370_/Q _5369_/Q _2673_/B vssd1 vssd1 vccd1 vccd1 _3598_/A sky130_fd_sc_hd__or3_4
X_5423_ _5423_/CLK _5423_/D vssd1 vssd1 vccd1 vccd1 _5423_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput223 _3685_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput212 _3675_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput234 _3670_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_145_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5354_ _5354_/CLK _5354_/D vssd1 vssd1 vccd1 vccd1 _5354_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput256 _3657_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput267 _3638_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__clkbuf_2
Xoutput245 _3647_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__clkbuf_2
X_4305_ _4304_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5672_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2566_ _3562_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _2574_/S sky130_fd_sc_hd__or2_4
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2497_ _2497_/A _2497_/B _2497_/C _2497_/D vssd1 vssd1 vccd1 vccd1 _2497_/Y sky130_fd_sc_hd__nor4_4
Xoutput278 _5850_/X vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_12
Xoutput289 _5860_/X vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_12
X_5285_ _5285_/CLK _5285_/D vssd1 vssd1 vccd1 vccd1 _5285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4532__117 _5730_/CLK vssd1 vssd1 vccd1 vccd1 _5174_/CLK sky130_fd_sc_hd__inv_2
X_4236_ _5562_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4236_/X sky130_fd_sc_hd__or2_1
XFILLER_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4167_ _4253_/A _4167_/B _4167_/C vssd1 vssd1 vccd1 vccd1 _4169_/D sky130_fd_sc_hd__nand3_1
XFILLER_110_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3118_ _3594_/A1 _5350_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5350_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4098_ _5541_/Q _5540_/Q _5539_/Q vssd1 vssd1 vccd1 vccd1 _4142_/B sky130_fd_sc_hd__nand3_4
X_3049_ _5162_/Q _5347_/Q _3066_/S vssd1 vssd1 vccd1 vccd1 _3049_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout450 _3140_/X vssd1 vssd1 vccd1 vccd1 _3333_/C1 sky130_fd_sc_hd__buf_6
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout483 _2866_/Y vssd1 vssd1 vccd1 vccd1 _3074_/A1 sky130_fd_sc_hd__buf_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout472 _3128_/Y vssd1 vssd1 vccd1 vccd1 _3301_/A1 sky130_fd_sc_hd__buf_6
XFILLER_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout461 _3355_/B vssd1 vssd1 vccd1 vccd1 _3171_/A sky130_fd_sc_hd__buf_6
Xfanout494 _3128_/B vssd1 vssd1 vccd1 vccd1 _3326_/B2 sky130_fd_sc_hd__buf_6
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4452__37 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5046_/CLK sky130_fd_sc_hd__inv_2
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_4_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5084_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold909 hold909/A vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__buf_2
XFILLER_6_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _5755_/CLK _5070_/D vssd1 vssd1 vccd1 vccd1 _5070_/Q sky130_fd_sc_hd__dfxtp_1
X_4021_ _5675_/Q _4021_/B _4021_/C _4029_/C vssd1 vssd1 vccd1 vccd1 _4071_/B sky130_fd_sc_hd__nand4_4
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1609 hold2450/X vssd1 vssd1 vccd1 vccd1 hold2451/A sky130_fd_sc_hd__buf_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4867__452 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5588_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4908__493 _5022_/CLK vssd1 vssd1 vccd1 vccd1 _5629_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3805_ hold277/X _5256_/Q _3814_/A3 _3814_/B1 _5005_/Q vssd1 vssd1 vccd1 vccd1 _3805_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3736_ _3824_/A1 _3734_/X _3735_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3736_/X sky130_fd_sc_hd__o211a_4
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3667_ _3667_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__and2_1
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5406_ _5406_/CLK _5406_/D vssd1 vssd1 vccd1 vccd1 _5406_/Q sky130_fd_sc_hd__dfxtp_1
X_3598_ _3598_/A _3598_/B vssd1 vssd1 vccd1 vccd1 _3606_/S sky130_fd_sc_hd__nor2_8
X_2618_ _2776_/A _3066_/S vssd1 vssd1 vccd1 vccd1 _2862_/A sky130_fd_sc_hd__or2_1
XFILLER_142_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2549_ _5661_/Q _3390_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _5661_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5337_ _5337_/CLK _5337_/D vssd1 vssd1 vccd1 vccd1 _5337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2800 hold2800/A vssd1 vssd1 vccd1 vccd1 hold2800/X sky130_fd_sc_hd__buf_2
X_5268_ _5268_/CLK _5268_/D vssd1 vssd1 vccd1 vccd1 _5268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2844 _4083_/X vssd1 vssd1 vccd1 vccd1 hold2844/X sky130_fd_sc_hd__buf_2
X_4219_ _5530_/Q _4186_/B _4165_/Y _5555_/Q vssd1 vssd1 vccd1 vccd1 _4221_/B sky130_fd_sc_hd__a31o_1
X_5199_ _5199_/CLK _5199_/D vssd1 vssd1 vccd1 vccd1 _5199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2899 hold2907/X vssd1 vssd1 vccd1 vccd1 hold2908/A sky130_fd_sc_hd__buf_2
XFILLER_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2888 hold2888/A vssd1 vssd1 vccd1 vccd1 hold2888/X sky130_fd_sc_hd__buf_2
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4660__245 _4433__18/A vssd1 vssd1 vccd1 vccd1 _5348_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4701__286 _5247_/CLK vssd1 vssd1 vccd1 vccd1 _5392_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3521_ _5142_/Q _3611_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5142_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold728 hold728/A vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__buf_2
Xhold717 hold717/A vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__buf_2
X_3452_ _3615_/A1 _5210_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5210_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap458 _2615_/Y vssd1 vssd1 vccd1 vccd1 _4001_/A3 sky130_fd_sc_hd__clkbuf_2
Xhold739 hold760/X vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__buf_2
XFILLER_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3383_ _5297_/Q _3566_/A1 _3387_/S vssd1 vssd1 vccd1 vccd1 _5297_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5122_ _5122_/CLK _5122_/D vssd1 vssd1 vccd1 vccd1 _5122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2118 hold488/X vssd1 vssd1 vccd1 vccd1 hold2118/X sky130_fd_sc_hd__buf_2
Xhold2129 _3865_/X vssd1 vssd1 vccd1 vccd1 hold2129/X sky130_fd_sc_hd__buf_2
XFILLER_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1428 hold2088/X vssd1 vssd1 vccd1 vccd1 hold2089/A sky130_fd_sc_hd__buf_2
Xhold1439 hold2104/X vssd1 vssd1 vccd1 vccd1 hold2105/A sky130_fd_sc_hd__buf_2
X_5053_ _5053_/CLK _5053_/D vssd1 vssd1 vccd1 vccd1 _5053_/Q sky130_fd_sc_hd__dfxtp_1
X_4004_ _5667_/Q _5666_/Q _5665_/Q vssd1 vssd1 vccd1 vccd1 _4259_/B sky130_fd_sc_hd__nand3_2
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4644__229 _4658__243/A vssd1 vssd1 vccd1 vccd1 _5330_/CLK sky130_fd_sc_hd__inv_2
X_5886_ _5886_/A vssd1 vssd1 vccd1 vccd1 _5886_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3719_ _5076_/Q input4/X _3728_/S vssd1 vssd1 vccd1 vccd1 _3719_/X sky130_fd_sc_hd__mux2_4
X_4538__123 _4418__3/A vssd1 vssd1 vccd1 vccd1 _5180_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2630 hold2630/A vssd1 vssd1 vccd1 vccd1 hold2630/X sky130_fd_sc_hd__buf_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__buf_2
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__buf_2
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__buf_2
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2641 _3795_/X vssd1 vssd1 vccd1 vccd1 hold2641/X sky130_fd_sc_hd__buf_2
Xhold2663 hold2663/A vssd1 vssd1 vccd1 vccd1 hold2663/X sky130_fd_sc_hd__buf_2
Xhold2674 hold262/X vssd1 vssd1 vccd1 vccd1 hold2674/X sky130_fd_sc_hd__buf_2
Xhold55 hold87/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__buf_2
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__buf_2
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1951 hold1951/A vssd1 vssd1 vccd1 vccd1 _4374_/B1 sky130_fd_sc_hd__buf_2
Xhold1962 _3957_/X vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__buf_2
Xhold1940 hold1940/A vssd1 vssd1 vccd1 vccd1 _4383_/B1 sky130_fd_sc_hd__buf_2
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__buf_2
Xhold2696 hold2696/A vssd1 vssd1 vccd1 vccd1 hold2696/X sky130_fd_sc_hd__buf_2
Xhold66 hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__buf_2
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__buf_2
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold77 hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__buf_2
XFILLER_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1995 hold1995/A vssd1 vssd1 vccd1 vccd1 _5743_/D sky130_fd_sc_hd__buf_2
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _5694_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _5010_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2952_ _3029_/B1 _2942_/X _2951_/X vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__a21o_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5740_ _5742_/CLK _5740_/D vssd1 vssd1 vccd1 vccd1 _5740_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2883_ _5368_/Q _2883_/B vssd1 vssd1 vccd1 vccd1 _2883_/X sky130_fd_sc_hd__xor2_4
X_5671_ _5731_/CLK _5671_/D vssd1 vssd1 vccd1 vccd1 _5671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3504_ _5157_/Q _3603_/A1 _3507_/S vssd1 vssd1 vccd1 vccd1 _5157_/D sky130_fd_sc_hd__mux2_1
Xhold503 hold503/A vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__buf_2
Xhold536 _3890_/X vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__buf_2
Xhold525 hold579/X vssd1 vssd1 vccd1 vccd1 hold580/A sky130_fd_sc_hd__buf_2
XFILLER_144_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3435_ _5225_/Q _3590_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5225_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3366_ _3603_/A1 _5313_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5313_/D sky130_fd_sc_hd__mux2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5252_/CLK _5105_/D vssd1 vssd1 vccd1 vccd1 _5105_/Q sky130_fd_sc_hd__dfxtp_1
X_4488__73 _4504__89/A vssd1 vssd1 vccd1 vccd1 _5130_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1225 hold1926/X vssd1 vssd1 vccd1 vccd1 hold1927/A sky130_fd_sc_hd__buf_2
Xhold1214 hold1921/X vssd1 vssd1 vccd1 vccd1 hold1922/A sky130_fd_sc_hd__buf_2
X_3297_ _3328_/A _3297_/B vssd1 vssd1 vccd1 vccd1 _3297_/X sky130_fd_sc_hd__or2_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5036_/CLK _5036_/D vssd1 vssd1 vccd1 vccd1 _5036_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1247 hold2281/X vssd1 vssd1 vccd1 vccd1 hold2282/A sky130_fd_sc_hd__buf_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1269 hold2502/X vssd1 vssd1 vccd1 vccd1 hold2503/A sky130_fd_sc_hd__buf_2
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5869_ _5869_/A vssd1 vssd1 vccd1 vccd1 _5869_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4772__357 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5463_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput101 probe_out[69] vssd1 vssd1 vccd1 vccd1 _5906_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput123 probe_out[89] vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__clkbuf_2
Xinput112 probe_out[79] vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput145 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _2492_/A sky130_fd_sc_hd__clkbuf_2
X_4813__398 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5504_/CLK sky130_fd_sc_hd__inv_2
Xinput134 wb_rst_i vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2471 hold2844/X vssd1 vssd1 vccd1 vccd1 hold2471/X sky130_fd_sc_hd__buf_2
Xinput167 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__buf_6
Xhold2460 hold2460/A vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__buf_2
Xinput178 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__clkbuf_8
Xinput156 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput189 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__buf_4
X_4666__251 _4477__62/A vssd1 vssd1 vccd1 vccd1 _5354_/CLK sky130_fd_sc_hd__inv_2
Xhold1781 hold2499/X vssd1 vssd1 vccd1 vccd1 hold2500/A sky130_fd_sc_hd__buf_2
Xhold1792 hold2529/X vssd1 vssd1 vccd1 vccd1 hold2530/A sky130_fd_sc_hd__buf_2
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4707__292 _5006_/CLK vssd1 vssd1 vccd1 vccd1 _5398_/CLK sky130_fd_sc_hd__inv_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_110_wb_clk_i _5743_/CLK vssd1 vssd1 vccd1 vccd1 _5543_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4676__261/A sky130_fd_sc_hd__clkbuf_8
X_3220_ _5500_/Q _5492_/Q _5484_/Q _5508_/Q _3312_/S _3130_/B vssd1 vssd1 vccd1 vccd1
+ _3220_/X sky130_fd_sc_hd__mux4_2
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3151_ _3320_/C1 _3141_/X _3334_/A1 vssd1 vssd1 vccd1 vccd1 _3151_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3082_ _3443_/B _3089_/A vssd1 vssd1 vccd1 vccd1 _3087_/A sky130_fd_sc_hd__and2_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3984_ _3648_/A _5253_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _5253_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2935_ _2863_/A _5380_/Q _3094_/A _2934_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _2935_/X
+ sky130_fd_sc_hd__a221o_1
X_5723_ _5723_/CLK _5723_/D vssd1 vssd1 vccd1 vccd1 _5723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2866_ _2866_/A _2866_/B vssd1 vssd1 vccd1 vccd1 _2866_/Y sky130_fd_sc_hd__nand2_1
X_5654_ _5654_/CLK _5654_/D vssd1 vssd1 vccd1 vccd1 _5654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold311 _3948_/X vssd1 vssd1 vccd1 vccd1 _5105_/D sky130_fd_sc_hd__buf_2
X_5585_ _5585_/CLK _5585_/D vssd1 vssd1 vccd1 vccd1 _5585_/Q sky130_fd_sc_hd__dfxtp_1
X_2797_ _5371_/Q _3443_/B _5373_/Q vssd1 vssd1 vccd1 vccd1 _2843_/B sky130_fd_sc_hd__nand3b_4
Xhold300 _3930_/Y vssd1 vssd1 vccd1 vccd1 _3931_/C sky130_fd_sc_hd__buf_2
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold322 _3950_/X vssd1 vssd1 vccd1 vccd1 _5107_/D sky130_fd_sc_hd__buf_2
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold355 hold355/A vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__buf_2
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold377 hold377/A vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__buf_2
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold388 _3965_/X vssd1 vssd1 vccd1 vccd1 _5204_/D sky130_fd_sc_hd__buf_2
X_3418_ _3591_/A1 _5240_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5240_/D sky130_fd_sc_hd__mux2_1
Xhold399 hold399/A vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__buf_2
X_4398_ _5747_/Q _4398_/A2 _4397_/X hold711/A vssd1 vssd1 vccd1 vccd1 _5747_/D sky130_fd_sc_hd__o211a_1
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1000 hold1554/X vssd1 vssd1 vccd1 vccd1 hold1555/A sky130_fd_sc_hd__buf_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ _3349_/A _3349_/B vssd1 vssd1 vccd1 vccd1 _5332_/D sky130_fd_sc_hd__nor2_1
Xhold1022 hold2444/X vssd1 vssd1 vccd1 vccd1 hold2445/A sky130_fd_sc_hd__buf_2
Xhold1011 hold2438/X vssd1 vssd1 vccd1 vccd1 hold1577/A sky130_fd_sc_hd__buf_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1066 hold2207/X vssd1 vssd1 vccd1 vccd1 hold2208/A sky130_fd_sc_hd__buf_2
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1044 hold195/X vssd1 vssd1 vccd1 vccd1 input205/A sky130_fd_sc_hd__buf_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5019_ _5019_/CLK _5019_/D vssd1 vssd1 vccd1 vccd1 _5019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1099 hold2366/X vssd1 vssd1 vccd1 vccd1 hold2367/A sky130_fd_sc_hd__buf_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2290 hold979/X vssd1 vssd1 vccd1 vccd1 hold2290/X sky130_fd_sc_hd__buf_2
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2720_ _3308_/A1 _5506_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5506_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2651_ _5593_/Q _3577_/A0 _2653_/S vssd1 vssd1 vccd1 vccd1 _5593_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5370_ _5370_/CLK _5370_/D vssd1 vssd1 vccd1 vccd1 _5370_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2582_ _3577_/A0 _5633_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5633_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4321_ _5664_/Q _4078_/A _5663_/Q vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__a21o_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4252_ _5741_/Q _4270_/B _4251_/X vssd1 vssd1 vccd1 vccd1 _4268_/B sky130_fd_sc_hd__o21ba_1
XFILLER_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3203_ _3316_/C1 _3200_/X _3202_/X vssd1 vssd1 vccd1 vccd1 _3203_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _5539_/Q _4186_/A vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__nor2_1
X_4418__3 _4418__3/A vssd1 vssd1 vccd1 vccd1 _4969_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4458__43 _5564_/CLK vssd1 vssd1 vccd1 vccd1 _5052_/CLK sky130_fd_sc_hd__inv_2
X_3134_ _5329_/Q _3138_/B vssd1 vssd1 vccd1 vccd1 _3140_/A sky130_fd_sc_hd__and2_4
X_3065_ _3099_/B _3063_/X _3064_/X vssd1 vssd1 vccd1 vccd1 _3065_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _5379_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _5206_/D sky130_fd_sc_hd__and2_1
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2918_ _5143_/Q _5151_/Q _5215_/Q _5135_/Q _3036_/S _2943_/S1 vssd1 vssd1 vccd1 vccd1
+ _2918_/X sky130_fd_sc_hd__mux4_1
X_5706_ _5706_/CLK _5706_/D vssd1 vssd1 vccd1 vccd1 _5706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3898_ _3887_/X _3896_/X _3897_/X _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3898_/X sky130_fd_sc_hd__a22o_1
X_2849_ _5395_/Q _2849_/A1 _2851_/S vssd1 vssd1 vccd1 vccd1 _5395_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5637_ _5637_/CLK _5637_/D vssd1 vssd1 vccd1 vccd1 _5637_/Q sky130_fd_sc_hd__dfxtp_1
X_5568_ _5568_/CLK _5568_/D vssd1 vssd1 vccd1 vccd1 _5568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold141 hold76/X vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__buf_2
Xhold130 _3627_/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__buf_2
Xhold152 hold163/X vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__buf_2
XFILLER_144_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold163 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__buf_2
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 _4360_/A sky130_fd_sc_hd__buf_2
X_5499_ _5499_/CLK _5499_/D vssd1 vssd1 vccd1 vccd1 _5499_/Q sky130_fd_sc_hd__dfxtp_1
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__buf_2
XFILLER_144_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout621 _5319_/Q vssd1 vssd1 vccd1 vccd1 _2850_/A1 sky130_fd_sc_hd__buf_2
Xfanout610 _5321_/Q vssd1 vssd1 vccd1 vccd1 _3594_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout632 hold711/A vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__buf_4
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__buf_2
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout643 hold137/X vssd1 vssd1 vccd1 vccd1 hold1459/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4884__469 _5252_/CLK vssd1 vssd1 vccd1 vccd1 _5605_/CLK sky130_fd_sc_hd__inv_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4778__363 _5019_/CLK vssd1 vssd1 vccd1 vccd1 _5469_/CLK sky130_fd_sc_hd__inv_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3821_ _4355_/A _5020_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _5020_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3752_ _3752_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3752_/X sky130_fd_sc_hd__and2_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3683_ _5256_/Q _3688_/B vssd1 vssd1 vccd1 vccd1 _3683_/X sky130_fd_sc_hd__and2_1
XFILLER_118_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2703_ _3571_/A _3388_/B vssd1 vssd1 vccd1 vccd1 _2711_/S sky130_fd_sc_hd__or2_4
XFILLER_145_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2634_ _2778_/A _2634_/B vssd1 vssd1 vccd1 vccd1 _2673_/B sky130_fd_sc_hd__nand2_1
X_5422_ _5422_/CLK _5422_/D vssd1 vssd1 vccd1 vccd1 _5422_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput224 _3686_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__clkbuf_2
Xoutput213 _3676_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_145_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput235 _3663_/B vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__clkbuf_2
XFILLER_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5353_ _5353_/CLK _5353_/D vssd1 vssd1 vccd1 vccd1 _5353_/Q sky130_fd_sc_hd__dfxtp_1
X_2565_ _3579_/A0 _5647_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5647_/D sky130_fd_sc_hd__mux2_1
Xoutput257 _3658_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__clkbuf_2
Xoutput246 _3648_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput268 _3625_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4304_ _4264_/B _4308_/A2 _4308_/B1 _2446_/Y vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__o22a_1
XFILLER_141_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2496_ _2496_/A _2496_/B _2496_/C vssd1 vssd1 vccd1 vccd1 _2497_/D sky130_fd_sc_hd__or3_4
Xoutput279 _5851_/X vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_12
X_5284_ _5284_/CLK _5284_/D vssd1 vssd1 vccd1 vccd1 _5284_/Q sky130_fd_sc_hd__dfxtp_1
X_4571__156 _4432__17/A vssd1 vssd1 vccd1 vccd1 _5221_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4235_ _5340_/Q _4360_/B _4164_/B _4234_/X _4244_/S vssd1 vssd1 vccd1 vccd1 _5561_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4166_ _4167_/B _4167_/C _4253_/A vssd1 vssd1 vccd1 vccd1 _4169_/C sky130_fd_sc_hd__a21o_1
XFILLER_110_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3117_ _3593_/A1 _5351_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5351_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4097_ _5557_/Q _5530_/Q _4222_/B vssd1 vssd1 vccd1 vccd1 _4165_/B sky130_fd_sc_hd__and3_1
X_4612__197 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5286_/CLK sky130_fd_sc_hd__inv_2
XFILLER_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3048_ _3596_/A1 _2895_/Y _3047_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5376_/D sky130_fd_sc_hd__o211a_1
XFILLER_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4999_ _5739_/CLK _4999_/D vssd1 vssd1 vccd1 vccd1 _4999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout440 split3/A vssd1 vssd1 vccd1 vccd1 _4093_/B sky130_fd_sc_hd__buf_4
XFILLER_48_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout473 _3097_/B vssd1 vssd1 vccd1 vccd1 _2945_/A sky130_fd_sc_hd__buf_6
XFILLER_93_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout484 split1/A vssd1 vssd1 vccd1 vccd1 split5/A sky130_fd_sc_hd__buf_6
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout462 _3355_/B vssd1 vssd1 vccd1 vccd1 _3320_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout451 _3140_/X vssd1 vssd1 vccd1 vccd1 _3353_/B sky130_fd_sc_hd__buf_4
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout495 _3298_/B1 vssd1 vssd1 vccd1 vccd1 _3128_/B sky130_fd_sc_hd__buf_6
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_88_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4454__39/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5291_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4020_ _4021_/B _4065_/B _4029_/C vssd1 vssd1 vccd1 vccd1 _4020_/X sky130_fd_sc_hd__and3_1
X_4428__13 _4472__57/A vssd1 vssd1 vccd1 vccd1 _4979_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3804_ hold277/X _5255_/Q _3810_/A3 hold349/X _5004_/Q vssd1 vssd1 vccd1 vccd1 _5004_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3735_ _4998_/Q _3750_/B vssd1 vssd1 vccd1 vccd1 _3735_/X sky130_fd_sc_hd__or2_1
XFILLER_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3666_ _3666_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3666_/X sky130_fd_sc_hd__and2_1
X_5405_ _5405_/CLK _5405_/D vssd1 vssd1 vccd1 vccd1 _5405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3597_ _5026_/Q _3597_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5026_/D sky130_fd_sc_hd__mux2_1
X_2617_ _5370_/Q _2867_/B vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__xor2_2
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5336_ _5336_/CLK _5336_/D vssd1 vssd1 vccd1 vccd1 _5336_/Q sky130_fd_sc_hd__dfxtp_1
X_2548_ _5662_/Q _2853_/A1 _2555_/S vssd1 vssd1 vccd1 vccd1 _5662_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2812 _4090_/X vssd1 vssd1 vccd1 vccd1 hold2812/X sky130_fd_sc_hd__buf_2
Xhold2801 hold2801/A vssd1 vssd1 vccd1 vccd1 hold2801/X sky130_fd_sc_hd__buf_2
X_5267_ _5267_/CLK _5267_/D vssd1 vssd1 vccd1 vccd1 _5267_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2856 _4088_/X vssd1 vssd1 vccd1 vccd1 hold2856/X sky130_fd_sc_hd__buf_2
X_4218_ _5738_/Q _4181_/B _4186_/B _3836_/A _4165_/Y vssd1 vssd1 vccd1 vccd1 _4220_/B
+ sky130_fd_sc_hd__o221a_2
X_2479_ _5333_/Q _5332_/Q _5331_/Q vssd1 vssd1 vccd1 vccd1 _2486_/A sky130_fd_sc_hd__and3_1
X_5198_ _5198_/CLK _5198_/D vssd1 vssd1 vccd1 vccd1 _5198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2889 _2499_/X vssd1 vssd1 vccd1 vccd1 _4410_/A1 sky130_fd_sc_hd__buf_2
X_4149_ _4149_/A _4149_/B _4149_/C _4149_/D vssd1 vssd1 vccd1 vccd1 _4162_/C sky130_fd_sc_hd__and4_1
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4512__97 _5084_/CLK vssd1 vssd1 vccd1 vccd1 _5154_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940__525 _5244_/CLK vssd1 vssd1 vccd1 vccd1 _5661_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3520_ _5143_/Q _3610_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5143_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3451_ _3614_/A1 _5211_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5211_/D sky130_fd_sc_hd__mux2_1
Xmax_cap459 _2615_/Y vssd1 vssd1 vccd1 vccd1 _3832_/A3 sky130_fd_sc_hd__clkbuf_2
XFILLER_143_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3382_ _5298_/Q _3574_/A0 _3387_/S vssd1 vssd1 vccd1 vccd1 _5298_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5121_ _5121_/CLK _5121_/D vssd1 vssd1 vccd1 vccd1 _5121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2119 hold2119/A vssd1 vssd1 vccd1 vccd1 _3870_/B1 sky130_fd_sc_hd__buf_2
XFILLER_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _5052_/CLK _5052_/D vssd1 vssd1 vccd1 vccd1 _5052_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1418 hold2714/X vssd1 vssd1 vccd1 vccd1 hold2075/A sky130_fd_sc_hd__buf_2
Xhold1429 hold2090/X vssd1 vssd1 vccd1 vccd1 hold2091/A sky130_fd_sc_hd__buf_2
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4003_ _5676_/Q _5675_/Q _5674_/Q _5673_/Q vssd1 vssd1 vccd1 vccd1 _4011_/A sky130_fd_sc_hd__nand4_1
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4683__268 _4425__10/A vssd1 vssd1 vccd1 vccd1 _5372_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3718_ _3718_/A1 _3716_/X _3717_/X split2/X vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__o211a_1
X_3649_ _3649_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3649_/X sky130_fd_sc_hd__or2_1
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4577__162 _4433__18/A vssd1 vssd1 vccd1 vccd1 _5227_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5319_ _5684_/CLK _5319_/D vssd1 vssd1 vccd1 vccd1 _5319_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__buf_2
Xhold2620 hold2620/A vssd1 vssd1 vccd1 vccd1 hold774/A sky130_fd_sc_hd__buf_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__buf_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__buf_2
Xhold2664 hold2664/A vssd1 vssd1 vccd1 vccd1 hold2664/X sky130_fd_sc_hd__buf_2
Xhold2642 hold2642/A vssd1 vssd1 vccd1 vccd1 hold2642/X sky130_fd_sc_hd__buf_2
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__buf_2
Xhold56 hold91/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__buf_2
XFILLER_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1930 _4376_/X vssd1 vssd1 vccd1 vccd1 hold1930/X sky130_fd_sc_hd__buf_2
Xhold1952 _4374_/X vssd1 vssd1 vccd1 vccd1 hold1952/X sky130_fd_sc_hd__buf_2
Xhold1963 hold181/X vssd1 vssd1 vccd1 vccd1 _3960_/B sky130_fd_sc_hd__buf_2
Xhold1941 _4383_/X vssd1 vssd1 vccd1 vccd1 hold1941/X sky130_fd_sc_hd__buf_2
Xhold2697 hold2697/A vssd1 vssd1 vccd1 vccd1 hold377/A sky130_fd_sc_hd__buf_2
Xhold2675 hold2675/A vssd1 vssd1 vccd1 vccd1 hold2675/X sky130_fd_sc_hd__buf_2
Xhold2686 _3791_/X vssd1 vssd1 vccd1 vccd1 hold2686/X sky130_fd_sc_hd__buf_2
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__buf_2
Xhold67 hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__buf_2
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__buf_2
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924__509 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5645_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4818__403 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5509_/CLK sky130_fd_sc_hd__inv_2
XANTENNA_9 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _3004_/C1 _2941_/X _3075_/B1 vssd1 vssd1 vccd1 vccd1 _2951_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4506__91/A
+ sky130_fd_sc_hd__clkbuf_16
X_5670_ _5725_/CLK _5670_/D vssd1 vssd1 vccd1 vccd1 _5670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2882_ _5368_/Q _2883_/B vssd1 vssd1 vccd1 vccd1 _3094_/B sky130_fd_sc_hd__xnor2_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3503_ _5158_/Q _3584_/A0 _3507_/S vssd1 vssd1 vccd1 vccd1 _5158_/D sky130_fd_sc_hd__mux2_1
Xhold504 hold504/A vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__buf_2
Xhold526 _3879_/X vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__buf_2
XFILLER_116_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3434_ _3526_/A _3589_/B vssd1 vssd1 vccd1 vccd1 _3442_/S sky130_fd_sc_hd__nor2_8
XFILLER_89_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold537 _3891_/X vssd1 vssd1 vccd1 vccd1 _5072_/D sky130_fd_sc_hd__buf_2
Xhold548 hold548/A vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__buf_2
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3365_ _3584_/A0 _5314_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5314_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5252_/CLK _5104_/D vssd1 vssd1 vccd1 vccd1 _5104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1204 hold1893/X vssd1 vssd1 vccd1 vccd1 hold1894/A sky130_fd_sc_hd__buf_2
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3296_ _5656_/Q _5386_/Q _3327_/S vssd1 vssd1 vccd1 vccd1 _3297_/B sky130_fd_sc_hd__mux2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/CLK _5035_/D vssd1 vssd1 vccd1 vccd1 _5035_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1226 hold1928/X vssd1 vssd1 vccd1 vccd1 hold1929/A sky130_fd_sc_hd__buf_2
Xhold1248 hold2285/X vssd1 vssd1 vccd1 vccd1 hold2286/A sky130_fd_sc_hd__buf_2
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _5868_/A vssd1 vssd1 vccd1 vccd1 _5868_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput102 probe_out[6] vssd1 vssd1 vccd1 vccd1 _5843_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput124 probe_out[8] vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__clkbuf_2
Xinput113 probe_out[7] vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__clkbuf_2
Xinput135 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _3661_/A sky130_fd_sc_hd__buf_4
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2472 hold2472/A vssd1 vssd1 vccd1 vccd1 hold2472/X sky130_fd_sc_hd__buf_2
XFILLER_56_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput157 input157/A vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__buf_4
Xinput146 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _3662_/A sky130_fd_sc_hd__buf_4
Xinput168 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__buf_8
Xhold2461 hold42/X vssd1 vssd1 vccd1 vccd1 hold2461/X sky130_fd_sc_hd__buf_2
Xhold2450 hold2450/A vssd1 vssd1 vccd1 vccd1 hold2450/X sky130_fd_sc_hd__buf_2
Xhold1771 hold2484/X vssd1 vssd1 vccd1 vccd1 hold2485/A sky130_fd_sc_hd__buf_2
XFILLER_57_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput179 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _4351_/B sky130_fd_sc_hd__buf_8
Xhold1782 hold2501/X vssd1 vssd1 vccd1 vccd1 hold2502/A sky130_fd_sc_hd__buf_2
XFILLER_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _3145_/X _3148_/X _3149_/X _3334_/A1 _3169_/B vssd1 vssd1 vccd1 vccd1 _3150_/X
+ sky130_fd_sc_hd__o221a_2
X_3081_ _3081_/A _3081_/B vssd1 vssd1 vccd1 vccd1 _3089_/A sky130_fd_sc_hd__nor2_1
X_4946__531 _4965__550/A vssd1 vssd1 vccd1 vccd1 _5704_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3983_ _3647_/A _5252_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3983_/X sky130_fd_sc_hd__mux2_1
X_5722_ _5722_/CLK _5722_/D vssd1 vssd1 vccd1 vccd1 _5722_/Q sky130_fd_sc_hd__dfxtp_1
X_2934_ _2883_/X _2931_/X _2933_/X _2929_/X vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__a31o_2
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2865_ _2867_/B _3063_/S vssd1 vssd1 vccd1 vccd1 _2865_/X sky130_fd_sc_hd__or2_1
X_5653_ _5653_/CLK _5653_/D vssd1 vssd1 vccd1 vccd1 _5653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5584_ _5584_/CLK _5584_/D vssd1 vssd1 vccd1 vccd1 _5584_/Q sky130_fd_sc_hd__dfxtp_1
XCaravelHost_730 vssd1 vssd1 vccd1 vccd1 partID[14] CaravelHost_730/LO sky130_fd_sc_hd__conb_1
Xhold301 _3931_/X vssd1 vssd1 vccd1 vccd1 hold327/A sky130_fd_sc_hd__buf_2
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2796_ _3396_/A0 _5441_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5441_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold356 hold356/A vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__buf_2
Xhold367 hold367/A vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__buf_2
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3417_ _3590_/A1 _5241_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5241_/D sky130_fd_sc_hd__mux2_1
X_4397_ _3637_/A _4357_/B _4398_/A2 vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__a21bo_1
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3348_ _5332_/Q _2489_/Y split3/X vssd1 vssd1 vccd1 vccd1 _3349_/B sky130_fd_sc_hd__o21ai_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1001 hold1556/X vssd1 vssd1 vccd1 vccd1 hold1557/A sky130_fd_sc_hd__buf_2
Xhold1012 hold1578/X vssd1 vssd1 vccd1 vccd1 hold1579/A sky130_fd_sc_hd__buf_2
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 hold1588/X vssd1 vssd1 vccd1 vccd1 hold1589/A sky130_fd_sc_hd__buf_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4689__274 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5378_/CLK sky130_fd_sc_hd__inv_2
Xhold1045 _3624_/A vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__buf_2
X_3279_ _5466_/Q _3331_/A2 _3237_/B _5624_/Q _3171_/A vssd1 vssd1 vccd1 vccd1 _3279_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _5019_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 _5018_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1078 hold2806/X vssd1 vssd1 vccd1 vccd1 hold2807/A sky130_fd_sc_hd__buf_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2280 hold2831/X vssd1 vssd1 vccd1 vccd1 hold2832/A sky130_fd_sc_hd__buf_2
XFILLER_91_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2291 hold2291/A vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__buf_2
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1590 hold46/X vssd1 vssd1 vccd1 vccd1 hold1590/X sky130_fd_sc_hd__buf_2
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2650_ _5594_/Q _3576_/A0 _2653_/S vssd1 vssd1 vccd1 vccd1 _5594_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2581_ _3576_/A0 _5634_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5634_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4320_ _5680_/Q _5664_/Q _5663_/Q vssd1 vssd1 vccd1 vccd1 _4320_/X sky130_fd_sc_hd__and3_1
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4251_ _5743_/Q _4023_/B _4270_/B _5741_/Q vssd1 vssd1 vccd1 vccd1 _4251_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3202_ _3320_/C1 _3201_/X _3336_/A1 vssd1 vssd1 vccd1 vccd1 _3202_/X sky130_fd_sc_hd__a21o_1
X_4182_ _5530_/Q _4177_/X _4184_/B vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3133_ _5504_/Q _5496_/Q _5488_/Q _5512_/Q _3281_/S _3130_/B vssd1 vssd1 vccd1 vccd1
+ _3133_/X sky130_fd_sc_hd__mux4_1
X_3064_ _2460_/A _5186_/Q _2866_/B _5194_/Q _3064_/C1 vssd1 vssd1 vccd1 vccd1 _3064_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4473__58 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5115_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4723__308 _4731__316/A vssd1 vssd1 vccd1 vccd1 _5414_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3966_ _5378_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__and2_1
X_2917_ _5119_/Q _5167_/Q _5352_/Q _5231_/Q _2944_/S0 _3066_/S vssd1 vssd1 vccd1 vccd1
+ _2917_/X sky130_fd_sc_hd__mux4_2
X_5705_ _5705_/CLK _5705_/D vssd1 vssd1 vccd1 vccd1 _5705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3897_ _5747_/Q _3914_/C _3897_/C vssd1 vssd1 vccd1 vccd1 _3897_/X sky130_fd_sc_hd__and3_1
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5636_ _5636_/CLK _5636_/D vssd1 vssd1 vccd1 vccd1 _5636_/Q sky130_fd_sc_hd__dfxtp_1
X_2848_ _5396_/Q _2848_/A1 _2851_/S vssd1 vssd1 vccd1 vccd1 _5396_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5567_ _5567_/CLK _5567_/D vssd1 vssd1 vccd1 vccd1 _5567_/Q sky130_fd_sc_hd__dfxtp_1
X_2779_ _2779_/A _3607_/A vssd1 vssd1 vccd1 vccd1 _2787_/S sky130_fd_sc_hd__nor2_8
XFILLER_117_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 _3988_/S sky130_fd_sc_hd__buf_2
XFILLER_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold153 hold165/X vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__buf_2
X_5498_ _5498_/CLK _5498_/D vssd1 vssd1 vccd1 vccd1 _5498_/Q sky130_fd_sc_hd__dfxtp_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__buf_2
Xhold142 hold164/X vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__buf_2
X_4617__202 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5294_/CLK sky130_fd_sc_hd__inv_2
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__buf_2
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__buf_2
Xhold175 hold34/X vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__buf_2
XFILLER_132_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout611 _5321_/Q vssd1 vssd1 vccd1 vccd1 _3612_/A1 sky130_fd_sc_hd__buf_2
Xfanout600 _2916_/A1 vssd1 vssd1 vccd1 vccd1 _3501_/A1 sky130_fd_sc_hd__buf_2
Xfanout622 _3606_/A1 vssd1 vssd1 vccd1 vccd1 _3597_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout633 hold875/A vssd1 vssd1 vccd1 vccd1 hold710/A sky130_fd_sc_hd__buf_4
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__buf_2
Xfanout644 _4360_/A vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__buf_8
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3820_ _4354_/A _5019_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _5019_/D sky130_fd_sc_hd__mux2_1
X_3751_ _3824_/A1 _3749_/X _3750_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3751_/X sky130_fd_sc_hd__o211a_4
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2702_ _5521_/Q _3579_/A0 _2702_/S vssd1 vssd1 vccd1 vccd1 _5521_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3682_ _5255_/Q _3682_/B vssd1 vssd1 vccd1 vccd1 _3682_/X sky130_fd_sc_hd__and2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2633_ _5383_/Q _4358_/B vssd1 vssd1 vccd1 vccd1 _3081_/B sky130_fd_sc_hd__nand2_4
X_5421_ _5421_/CLK _5421_/D vssd1 vssd1 vccd1 vccd1 _5421_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput225 _3687_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__clkbuf_2
Xoutput214 _3677_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__clkbuf_2
X_4420__5 _4423__8/A vssd1 vssd1 vccd1 vccd1 _4971_/CLK sky130_fd_sc_hd__inv_2
X_5352_ _5352_/CLK _5352_/D vssd1 vssd1 vccd1 vccd1 _5352_/Q sky130_fd_sc_hd__dfxtp_1
X_2564_ _3578_/A0 _5648_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5648_/D sky130_fd_sc_hd__mux2_1
Xoutput258 _3631_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput247 _3630_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput236 _3629_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4303_ _4302_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5671_/D sky130_fd_sc_hd__and2b_1
Xoutput269 _3626_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2495_ _2495_/A _2495_/B _2495_/C _2495_/D vssd1 vssd1 vccd1 vccd1 _2496_/C sky130_fd_sc_hd__or4_1
X_5283_ _5283_/CLK _5283_/D vssd1 vssd1 vccd1 vccd1 _5283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4234_ _5561_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4234_/X sky130_fd_sc_hd__or2_1
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4165_ _5529_/Q _4165_/B vssd1 vssd1 vccd1 vccd1 _4165_/Y sky130_fd_sc_hd__nor2_1
X_3116_ _3592_/A1 _5352_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5352_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _5556_/Q _5555_/Q vssd1 vssd1 vccd1 vccd1 _4222_/B sky130_fd_sc_hd__and2_1
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3047_ _2863_/A _5376_/Q _3094_/A _3046_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _3047_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4998_ _5739_/CLK _4998_/D vssd1 vssd1 vccd1 vccd1 _4998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3949_ _5253_/Q _5106_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _5106_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5619_ _5619_/CLK _5619_/D vssd1 vssd1 vccd1 vccd1 _5619_/Q sky130_fd_sc_hd__dfxtp_1
X_4851__436 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5572_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout430 _3753_/X vssd1 vssd1 vccd1 vccd1 _3774_/B1 sky130_fd_sc_hd__buf_8
Xfanout441 split3/X vssd1 vssd1 vccd1 vccd1 _3277_/C1 sky130_fd_sc_hd__clkbuf_2
Xfanout474 _3097_/B vssd1 vssd1 vccd1 vccd1 _3029_/B1 sky130_fd_sc_hd__buf_6
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout452 _3139_/Y vssd1 vssd1 vccd1 vccd1 _3334_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout463 _3355_/B vssd1 vssd1 vccd1 vccd1 _3323_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout485 split1/X vssd1 vssd1 vccd1 vccd1 hold821/A sky130_fd_sc_hd__buf_4
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout496 _3127_/X vssd1 vssd1 vccd1 vccd1 _3298_/B1 sky130_fd_sc_hd__buf_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4745__330 _5005_/CLK vssd1 vssd1 vccd1 vccd1 _5436_/CLK sky130_fd_sc_hd__inv_2
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4594__179 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5268_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_57_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _5005_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4443__28 _5001_/CLK vssd1 vssd1 vccd1 vccd1 _5037_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3803_ hold277/X _5254_/Q _3810_/A3 hold349/X _5003_/Q vssd1 vssd1 vccd1 vccd1 _5003_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3734_ _5081_/Q input9/X _3763_/B vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3665_ _3665_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__and2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5404_ _5404_/CLK _5404_/D vssd1 vssd1 vccd1 vccd1 _5404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2616_ _4352_/A split1/A _2615_/Y _3931_/A vssd1 vssd1 vccd1 vccd1 _4094_/C sky130_fd_sc_hd__a31oi_4
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3596_ _5027_/Q _3596_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5027_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5335_ _5335_/CLK _5335_/D vssd1 vssd1 vccd1 vccd1 _5335_/Q sky130_fd_sc_hd__dfxtp_4
X_2547_ _2852_/A _3571_/A vssd1 vssd1 vccd1 vccd1 _2555_/S sky130_fd_sc_hd__nor2_8
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2813 hold2813/A vssd1 vssd1 vccd1 vccd1 hold2813/X sky130_fd_sc_hd__buf_2
X_5266_ _5266_/CLK _5266_/D vssd1 vssd1 vccd1 vccd1 _5266_/Q sky130_fd_sc_hd__dfxtp_1
X_2478_ _5332_/Q _5331_/Q vssd1 vssd1 vccd1 vccd1 _2545_/A sky130_fd_sc_hd__nand2_4
XFILLER_102_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4217_ _4217_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _5554_/D sky130_fd_sc_hd__nor2_1
X_5197_ _5197_/CLK _5197_/D vssd1 vssd1 vccd1 vccd1 _5197_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2868 _4087_/X vssd1 vssd1 vccd1 vccd1 hold2868/X sky130_fd_sc_hd__buf_2
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4148_ _4171_/C _4148_/B vssd1 vssd1 vccd1 vccd1 _4149_/D sky130_fd_sc_hd__and2_1
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4729__314 _4731__316/A vssd1 vssd1 vccd1 vccd1 _5420_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _5682_/Q _5681_/Q vssd1 vssd1 vccd1 vccd1 _4080_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_104_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5553_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4522__107 _4439__24/A vssd1 vssd1 vccd1 vccd1 _5164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap405 _3598_/A vssd1 vssd1 vccd1 vccd1 _3526_/A sky130_fd_sc_hd__buf_12
Xhold708 hold872/X vssd1 vssd1 vccd1 vccd1 hold873/A sky130_fd_sc_hd__buf_2
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3450_ _3613_/A1 _5212_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5212_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3381_ _5299_/Q _3564_/A1 _3387_/S vssd1 vssd1 vccd1 vccd1 _5299_/D sky130_fd_sc_hd__mux2_1
X_5120_ _5120_/CLK _5120_/D vssd1 vssd1 vccd1 vccd1 _5120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2109 _3784_/X vssd1 vssd1 vccd1 vccd1 hold2109/X sky130_fd_sc_hd__buf_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5051_ _5051_/CLK _5051_/D vssd1 vssd1 vccd1 vccd1 _5051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4002_ _5674_/Q _5673_/Q vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__and2_2
XFILLER_78_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1419 hold2076/X vssd1 vssd1 vccd1 vccd1 hold2077/A sky130_fd_sc_hd__buf_2
XFILLER_84_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _5884_/A vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3717_ _4992_/Q _3729_/B vssd1 vssd1 vccd1 vccd1 _3717_/X sky130_fd_sc_hd__or2_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3648_ _3648_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__or2_1
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3579_ _3579_/A0 _5042_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5042_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5318_ _5684_/CLK _5318_/D vssd1 vssd1 vccd1 vccd1 _5318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2621 hold774/X vssd1 vssd1 vccd1 vccd1 hold2621/X sky130_fd_sc_hd__buf_2
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__buf_2
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5249_ _5739_/CLK _5249_/D vssd1 vssd1 vccd1 vccd1 _5249_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__buf_2
Xhold1920 hold1920/A vssd1 vssd1 vccd1 vccd1 hold853/A sky130_fd_sc_hd__buf_2
Xhold2654 _4092_/X vssd1 vssd1 vccd1 vccd1 hold2654/X sky130_fd_sc_hd__buf_2
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__buf_2
Xhold2643 hold2643/A vssd1 vssd1 vccd1 vccd1 hold2643/X sky130_fd_sc_hd__buf_2
Xhold2665 hold2665/A vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__buf_2
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__buf_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5697_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1931 hold1931/A vssd1 vssd1 vccd1 vccd1 hold590/A sky130_fd_sc_hd__buf_2
Xhold1953 hold1953/A vssd1 vssd1 vccd1 vccd1 hold804/A sky130_fd_sc_hd__buf_2
X_4963__548 _4964__549/A vssd1 vssd1 vccd1 vccd1 _5721_/CLK sky130_fd_sc_hd__inv_2
Xhold1942 hold1942/A vssd1 vssd1 vccd1 vccd1 hold863/A sky130_fd_sc_hd__buf_2
Xhold2698 hold377/X vssd1 vssd1 vccd1 vccd1 hold2698/X sky130_fd_sc_hd__buf_2
Xhold2687 hold2687/A vssd1 vssd1 vccd1 vccd1 hold2687/X sky130_fd_sc_hd__buf_2
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__buf_2
Xhold68 hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__buf_2
Xhold57 hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__buf_2
XFILLER_84_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1964 _3958_/X vssd1 vssd1 vccd1 vccd1 hold1964/X sky130_fd_sc_hd__buf_2
Xhold1986 hold2617/X vssd1 vssd1 vccd1 vccd1 hold2618/A sky130_fd_sc_hd__buf_2
XFILLER_44_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1975 hold2604/X vssd1 vssd1 vccd1 vccd1 hold2605/A sky130_fd_sc_hd__buf_2
XFILLER_17_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4857__442 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5578_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2950_ _2945_/A _2940_/X _2949_/X vssd1 vssd1 vccd1 vccd1 _2950_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2881_ _2947_/S _2878_/X _2880_/X vssd1 vssd1 vccd1 vccd1 _2881_/X sky130_fd_sc_hd__a21o_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_wb_clk_i clkbuf_4_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5738_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3502_ _5159_/Q _3538_/A0 _3507_/S vssd1 vssd1 vccd1 vccd1 _5159_/D sky130_fd_sc_hd__mux2_1
Xhold505 hold505/A vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__buf_2
Xhold527 _3880_/X vssd1 vssd1 vccd1 vccd1 _5070_/D sky130_fd_sc_hd__buf_2
XFILLER_143_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3433_ _5226_/Q _3597_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5226_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5252_/CLK _5103_/D vssd1 vssd1 vccd1 vccd1 _5103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3364_ _3538_/A0 _5315_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5315_/D sky130_fd_sc_hd__mux2_1
X_4650__235 _5751_/CLK vssd1 vssd1 vccd1 vccd1 _5336_/CLK sky130_fd_sc_hd__inv_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1205 hold1895/X vssd1 vssd1 vccd1 vccd1 hold1896/A sky130_fd_sc_hd__buf_2
XFILLER_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _2482_/B _5302_/Q _5051_/Q _3326_/B2 _3326_/C1 vssd1 vssd1 vccd1 vccd1 _3295_/X
+ sky130_fd_sc_hd__o221a_1
X_5034_ _5034_/CLK _5034_/D vssd1 vssd1 vccd1 vccd1 _5034_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1227 hold1930/X vssd1 vssd1 vccd1 vccd1 hold1931/A sky130_fd_sc_hd__buf_2
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5867_ _5867_/A vssd1 vssd1 vccd1 vccd1 _5867_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput125 probe_out[90] vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__clkbuf_2
Xinput114 probe_out[80] vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__clkbuf_2
Xinput103 probe_out[70] vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__clkbuf_2
X_4479__64 _4509__94/A vssd1 vssd1 vccd1 vccd1 _5121_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput136 input136/A vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__buf_6
Xhold2440 hold2440/A vssd1 vssd1 vccd1 vccd1 hold2440/X sky130_fd_sc_hd__buf_2
XFILLER_102_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2473 hold2473/A vssd1 vssd1 vccd1 vccd1 hold2473/X sky130_fd_sc_hd__buf_2
Xhold2451 hold2451/A vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__buf_2
Xinput169 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _3639_/A sky130_fd_sc_hd__clkbuf_8
Xhold2462 hold2462/A vssd1 vssd1 vccd1 vccd1 hold2462/X sky130_fd_sc_hd__buf_2
Xinput147 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _2492_/D sky130_fd_sc_hd__clkbuf_2
Xinput158 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _2493_/B sky130_fd_sc_hd__clkbuf_2
Xhold2484 hold2838/X vssd1 vssd1 vccd1 vccd1 hold2484/X sky130_fd_sc_hd__buf_2
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1772 hold2486/X vssd1 vssd1 vccd1 vccd1 hold2487/A sky130_fd_sc_hd__buf_2
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1783 hold2503/X vssd1 vssd1 vccd1 vccd1 hold2504/A sky130_fd_sc_hd__buf_2
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4634__219 _4514__99/A vssd1 vssd1 vccd1 vccd1 _5312_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3080_ _5374_/Q _5383_/Q _3080_/B1 _3081_/B vssd1 vssd1 vccd1 vccd1 _5374_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3982_ _3646_/A _5251_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3982_/X sky130_fd_sc_hd__mux2_1
X_4528__113 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5170_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2933_ _3029_/B1 _2926_/X _2932_/X vssd1 vssd1 vccd1 vccd1 _2933_/X sky130_fd_sc_hd__a21o_2
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5721_ _5721_/CLK _5721_/D vssd1 vssd1 vccd1 vccd1 _5721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2864_ _2867_/B _3063_/S vssd1 vssd1 vccd1 vccd1 _2866_/A sky130_fd_sc_hd__nand2_2
X_5652_ _5652_/CLK _5652_/D vssd1 vssd1 vccd1 vccd1 _5652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5583_ _5583_/CLK _5583_/D vssd1 vssd1 vccd1 vccd1 _5583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2795_ _3395_/A0 _5442_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5442_/D sky130_fd_sc_hd__mux2_1
XCaravelHost_720 vssd1 vssd1 vccd1 vccd1 CaravelHost_720/HI versionID[2] sky130_fd_sc_hd__conb_1
XCaravelHost_731 vssd1 vssd1 vccd1 vccd1 partID[15] CaravelHost_731/LO sky130_fd_sc_hd__conb_1
Xhold302 hold319/X vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__buf_2
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold357 hold357/A vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__buf_2
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3416_ _3508_/A _3589_/B vssd1 vssd1 vccd1 vccd1 _3424_/S sky130_fd_sc_hd__or2_4
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold379 hold379/A vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__buf_2
X_4396_ _5746_/Q _4398_/A2 _4395_/X _3778_/A vssd1 vssd1 vccd1 vccd1 _4396_/X sky130_fd_sc_hd__o211a_1
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ split3/X _3347_/B _3347_/C vssd1 vssd1 vccd1 vccd1 _5333_/D sky130_fd_sc_hd__and3_1
XFILLER_140_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1002 hold1558/X vssd1 vssd1 vccd1 vccd1 hold1559/A sky130_fd_sc_hd__buf_2
Xhold1013 hold1580/X vssd1 vssd1 vccd1 vccd1 hold1581/A sky130_fd_sc_hd__buf_2
Xhold1024 hold1590/X vssd1 vssd1 vccd1 vccd1 hold1591/A sky130_fd_sc_hd__buf_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 hold1119/X vssd1 vssd1 vccd1 vccd1 hold1120/A sky130_fd_sc_hd__buf_2
X_5017_ _5734_/CLK hold59/X vssd1 vssd1 vccd1 vccd1 _5017_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1035 hold2790/X vssd1 vssd1 vccd1 vccd1 hold2791/A sky130_fd_sc_hd__buf_2
Xhold1046 hold196/X vssd1 vssd1 vccd1 vccd1 hold149/A sky130_fd_sc_hd__buf_2
X_3278_ _5514_/Q _5283_/Q _3330_/S vssd1 vssd1 vccd1 vccd1 _3278_/X sky130_fd_sc_hd__mux2_2
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1068 hold2799/X vssd1 vssd1 vccd1 vccd1 hold2800/A sky130_fd_sc_hd__buf_2
Xhold1079 hold2196/X vssd1 vssd1 vccd1 vccd1 hold2197/A sky130_fd_sc_hd__buf_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5919_ _5919_/A vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2281 hold2281/A vssd1 vssd1 vccd1 vccd1 hold2281/X sky130_fd_sc_hd__buf_2
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2270 hold30/X vssd1 vssd1 vccd1 vccd1 hold2270/X sky130_fd_sc_hd__buf_2
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1580 _3933_/X vssd1 vssd1 vccd1 vccd1 hold1580/X sky130_fd_sc_hd__buf_2
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2292 hold27/X vssd1 vssd1 vccd1 vccd1 hold2292/X sky130_fd_sc_hd__buf_2
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1591 hold1591/A vssd1 vssd1 vccd1 vccd1 _3942_/A0 sky130_fd_sc_hd__buf_2
XFILLER_57_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2580_ _3575_/A0 _5635_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5635_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4250_ _4246_/Y _4247_/X _4248_/X _4249_/X _4016_/B vssd1 vssd1 vccd1 vccd1 _4268_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_141_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4181_ _5738_/Q _4181_/B vssd1 vssd1 vccd1 vccd1 _4184_/B sky130_fd_sc_hd__nor2_1
X_3201_ _5643_/Q _5635_/Q _5046_/Q _5651_/Q _3284_/S _3201_/S1 vssd1 vssd1 vccd1 vccd1
+ _3201_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3132_ _3132_/A _3138_/B vssd1 vssd1 vccd1 vccd1 _3132_/X sky130_fd_sc_hd__or2_1
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3063_ _4967_/Q _5178_/Q _3063_/S vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4762__347 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5453_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _5377_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _3965_/X sky130_fd_sc_hd__and2_1
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2916_ _2916_/A1 _2895_/Y _2915_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5381_/D sky130_fd_sc_hd__o211a_1
X_3896_ _3914_/C _5363_/Q _3897_/C _3855_/X vssd1 vssd1 vccd1 vccd1 _3896_/X sky130_fd_sc_hd__a31o_1
X_5704_ _5704_/CLK _5704_/D vssd1 vssd1 vccd1 vccd1 _5704_/Q sky130_fd_sc_hd__dfxtp_1
X_4803__388 _4898__483/A vssd1 vssd1 vccd1 vccd1 _5494_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2847_ _5397_/Q _5322_/Q _2851_/S vssd1 vssd1 vccd1 vccd1 _5397_/D sky130_fd_sc_hd__mux2_1
X_5635_ _5635_/CLK _5635_/D vssd1 vssd1 vccd1 vccd1 _5635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold110 _3983_/X vssd1 vssd1 vccd1 vccd1 _5252_/D sky130_fd_sc_hd__buf_2
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2778_ _2778_/A _3091_/A vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__nand2_8
X_5566_ _5566_/CLK _5566_/D vssd1 vssd1 vccd1 vccd1 _5566_/Q sky130_fd_sc_hd__dfxtp_1
Xhold121 _3982_/X vssd1 vssd1 vccd1 vccd1 _5251_/D sky130_fd_sc_hd__buf_2
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4656__241 _4459__44/A vssd1 vssd1 vccd1 vccd1 _5342_/CLK sky130_fd_sc_hd__inv_2
Xhold143 hold168/X vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__buf_2
X_5497_ _5497_/CLK _5497_/D vssd1 vssd1 vccd1 vccd1 _5497_/Q sky130_fd_sc_hd__dfxtp_1
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__buf_2
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__buf_2
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__buf_2
Xhold154 hold167/X vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__buf_2
XFILLER_144_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout623 _3606_/A1 vssd1 vssd1 vccd1 vccd1 _3615_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout601 _5324_/Q vssd1 vssd1 vccd1 vccd1 _2916_/A1 sky130_fd_sc_hd__buf_6
Xfanout612 _5321_/Q vssd1 vssd1 vccd1 vccd1 _3603_/A1 sky130_fd_sc_hd__buf_4
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__buf_2
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__buf_2
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _3645_/A _3778_/B _4370_/X vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__a21bo_1
Xfanout645 _4390_/A vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__buf_6
Xfanout634 hold875/A vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4449__34 _4449__34/A vssd1 vssd1 vccd1 vccd1 _5043_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _5003_/Q _3750_/B vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__or2_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2701_ _5522_/Q _3569_/A1 _2702_/S vssd1 vssd1 vccd1 vccd1 _5522_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3681_ _5254_/Q _3682_/B vssd1 vssd1 vccd1 vccd1 _3681_/X sky130_fd_sc_hd__and2_1
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2632_ _5383_/Q _4358_/B vssd1 vssd1 vccd1 vccd1 _2634_/B sky130_fd_sc_hd__and2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5420_ _5420_/CLK _5420_/D vssd1 vssd1 vccd1 vccd1 _5420_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput226 _3688_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput215 _3678_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5351_ _5351_/CLK _5351_/D vssd1 vssd1 vccd1 vccd1 _5351_/Q sky130_fd_sc_hd__dfxtp_1
X_2563_ _3577_/A0 _5649_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5649_/D sky130_fd_sc_hd__mux2_1
Xoutput259 _3659_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__clkbuf_2
Xoutput248 _3649_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput237 _3639_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__clkbuf_2
X_4302_ _4253_/B _4308_/A2 _4308_/B1 _4034_/A vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__o22a_1
X_5282_ _5282_/CLK _5282_/D vssd1 vssd1 vccd1 vccd1 _5282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _5339_/Q _4360_/B _4164_/B _4232_/X _4244_/S vssd1 vssd1 vccd1 vccd1 _5560_/D
+ sky130_fd_sc_hd__o311a_1
X_2494_ _2494_/A _2494_/B input155/X input156/X vssd1 vssd1 vccd1 vccd1 _2496_/B sky130_fd_sc_hd__or4bb_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4164_ _4360_/B _4164_/B vssd1 vssd1 vccd1 vccd1 _4242_/B sky130_fd_sc_hd__nor2_4
X_3115_ _3591_/A1 _5353_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5353_/D sky130_fd_sc_hd__mux2_1
X_4095_ _4095_/A _4095_/B vssd1 vssd1 vccd1 vccd1 _4095_/X sky130_fd_sc_hd__and2_1
XFILLER_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046_ _3094_/B _3042_/X _3043_/X _3045_/X vssd1 vssd1 vccd1 vccd1 _3046_/X sky130_fd_sc_hd__a31o_1
XFILLER_82_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4997_ _5248_/CLK _4997_/D vssd1 vssd1 vccd1 vccd1 _4997_/Q sky130_fd_sc_hd__dfxtp_1
X_3948_ _5252_/Q _5105_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _3948_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3879_ _4399_/B _3876_/X _3878_/X hold554/X vssd1 vssd1 vccd1 vccd1 _3879_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5618_ _5618_/CLK _5618_/D vssd1 vssd1 vccd1 vccd1 _5618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5549_ _5551_/CLK _5549_/D vssd1 vssd1 vccd1 vccd1 _5549_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4890__475 _4898__483/A vssd1 vssd1 vccd1 vccd1 _5611_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout431 _3621_/X vssd1 vssd1 vccd1 vccd1 _3638_/B sky130_fd_sc_hd__buf_4
Xfanout420 _4319_/B vssd1 vssd1 vccd1 vccd1 _4082_/A sky130_fd_sc_hd__buf_4
XFILLER_59_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout475 _2870_/X vssd1 vssd1 vccd1 vccd1 _3097_/B sky130_fd_sc_hd__buf_6
XFILLER_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout442 _4091_/A vssd1 vssd1 vccd1 vccd1 split3/A sky130_fd_sc_hd__buf_6
Xfanout464 _3132_/X vssd1 vssd1 vccd1 vccd1 _3355_/B sky130_fd_sc_hd__buf_4
Xfanout453 _3139_/Y vssd1 vssd1 vccd1 vccd1 _3336_/A1 sky130_fd_sc_hd__buf_2
Xfanout497 _2868_/Y vssd1 vssd1 vccd1 vccd1 _2870_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout486 _2498_/X vssd1 vssd1 vccd1 vccd1 split1/A sky130_fd_sc_hd__buf_8
XFILLER_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_97_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4819__404/A
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_26_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4509__94/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3802_ hold277/X _5253_/Q _3810_/A3 hold349/X _5002_/Q vssd1 vssd1 vccd1 vccd1 _3802_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3733_ _3733_/A1 _3731_/X _3732_/X _3777_/A3 vssd1 vssd1 vccd1 vccd1 _3733_/X sky130_fd_sc_hd__o211a_1
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3664_ _3664_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3664_/X sky130_fd_sc_hd__and2_1
XFILLER_109_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4874__459 _4898__483/A vssd1 vssd1 vccd1 vccd1 _5595_/CLK sky130_fd_sc_hd__inv_2
XFILLER_146_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5403_ _5403_/CLK _5403_/D vssd1 vssd1 vccd1 vccd1 _5403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2615_ _4369_/A _3888_/A _4399_/C _3852_/A vssd1 vssd1 vccd1 vccd1 _2615_/Y sky130_fd_sc_hd__nor4_4
X_3595_ _5028_/Q _3595_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5028_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5334_ _5334_/CLK _5334_/D vssd1 vssd1 vccd1 vccd1 _5334_/Q sky130_fd_sc_hd__dfxtp_4
X_2546_ split3/A _3349_/A vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__nand2_8
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5265_ _5265_/CLK _5265_/D vssd1 vssd1 vccd1 vccd1 _5265_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2814 hold2814/A vssd1 vssd1 vccd1 vccd1 hold2814/X sky130_fd_sc_hd__buf_2
X_2477_ _5335_/Q _5330_/Q vssd1 vssd1 vccd1 vccd1 _3122_/C sky130_fd_sc_hd__xnor2_2
Xhold2803 _3797_/X vssd1 vssd1 vccd1 vccd1 hold2803/X sky130_fd_sc_hd__buf_2
XFILLER_141_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5196_ _5196_/CLK _5196_/D vssd1 vssd1 vccd1 vccd1 _5196_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2825 _3778_/X vssd1 vssd1 vccd1 vccd1 hold2825/X sky130_fd_sc_hd__buf_2
X_4216_ _5554_/Q _4209_/B _4186_/X _4107_/B vssd1 vssd1 vccd1 vccd1 _4217_/B sky130_fd_sc_hd__o2bb2a_1
Xhold2869 _4390_/A vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__buf_2
X_4147_ _4128_/B _4128_/C _5749_/Q vssd1 vssd1 vccd1 vccd1 _4148_/B sky130_fd_sc_hd__a21bo_1
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4768__353 _5734_/CLK vssd1 vssd1 vccd1 vccd1 _5459_/CLK sky130_fd_sc_hd__inv_2
X_4078_ _4078_/A _4324_/A vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__nor2_4
XFILLER_56_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3029_ _5059_/Q _3073_/B2 _3029_/B1 _3028_/X vssd1 vssd1 vccd1 vccd1 _3029_/X sky130_fd_sc_hd__o211a_1
XFILLER_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4809__394 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5500_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4561__146 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5211_/CLK sky130_fd_sc_hd__inv_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold709 hold874/X vssd1 vssd1 vccd1 vccd1 hold875/A sky130_fd_sc_hd__buf_2
X_4602__187 _4456__41/A vssd1 vssd1 vccd1 vccd1 _5276_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3380_ _5300_/Q _3572_/A0 _3387_/S vssd1 vssd1 vccd1 vccd1 _5300_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5050_ _5050_/CLK _5050_/D vssd1 vssd1 vccd1 vccd1 _5050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4503__88 _4422__7/A vssd1 vssd1 vccd1 vccd1 _5145_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4001_ _4350_/A split1/X _4001_/A3 _4390_/A vssd1 vssd1 vccd1 vccd1 _4001_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5883_ _5883_/A vssd1 vssd1 vccd1 vccd1 _5883_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3716_ _5075_/Q input34/X _3728_/S vssd1 vssd1 vccd1 vccd1 _3716_/X sky130_fd_sc_hd__mux2_4
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3647_ _3647_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3647_/X sky130_fd_sc_hd__or2_1
X_3578_ _3578_/A0 _5043_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5043_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5317_ _5317_/CLK _5317_/D vssd1 vssd1 vccd1 vccd1 _5317_/Q sky130_fd_sc_hd__dfxtp_1
X_2529_ _3392_/A0 _5712_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5712_/D sky130_fd_sc_hd__mux2_1
Xhold2622 hold2622/A vssd1 vssd1 vccd1 vccd1 hold2622/X sky130_fd_sc_hd__buf_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__buf_2
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__buf_2
XFILLER_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2655 hold2655/A vssd1 vssd1 vccd1 vccd1 hold2655/X sky130_fd_sc_hd__buf_2
Xhold1910 hold858/X vssd1 vssd1 vccd1 vccd1 hold1910/X sky130_fd_sc_hd__buf_2
Xhold2633 _3793_/X vssd1 vssd1 vccd1 vccd1 hold2633/X sky130_fd_sc_hd__buf_2
Xhold2644 hold2644/A vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__buf_2
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__buf_2
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__buf_2
X_5248_ _5248_/CLK _5248_/D vssd1 vssd1 vccd1 vccd1 _5248_/Q sky130_fd_sc_hd__dfxtp_1
X_5179_ _5179_/CLK _5179_/D vssd1 vssd1 vccd1 vccd1 _5179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1932 hold590/X vssd1 vssd1 vccd1 vccd1 hold1932/X sky130_fd_sc_hd__buf_2
Xhold1954 hold804/X vssd1 vssd1 vccd1 vccd1 hold1954/X sky130_fd_sc_hd__buf_2
XFILLER_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1943 hold863/X vssd1 vssd1 vccd1 vccd1 hold1943/X sky130_fd_sc_hd__buf_2
Xhold1921 hold853/X vssd1 vssd1 vccd1 vccd1 hold1921/X sky130_fd_sc_hd__buf_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2666 hold253/X vssd1 vssd1 vccd1 vccd1 hold2666/X sky130_fd_sc_hd__buf_2
Xhold2688 hold2688/A vssd1 vssd1 vccd1 vccd1 hold2688/X sky130_fd_sc_hd__buf_2
Xhold69 hold96/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__buf_2
Xhold58 hold78/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__buf_2
Xhold1965 hold1965/A vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__buf_2
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1987 hold2619/X vssd1 vssd1 vccd1 vccd1 hold2620/A sky130_fd_sc_hd__buf_2
Xhold1976 hold2606/X vssd1 vssd1 vccd1 vccd1 hold2607/A sky130_fd_sc_hd__buf_2
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1998 hold2633/X vssd1 vssd1 vccd1 vccd1 hold2634/A sky130_fd_sc_hd__buf_2
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4896__481 _4921__506/A vssd1 vssd1 vccd1 vccd1 _5617_/CLK sky130_fd_sc_hd__inv_2
XFILLER_125_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2880_ _2945_/A _2879_/X _2919_/B vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__a21o_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3501_ _5160_/Q _3501_/A1 _3507_/S vssd1 vssd1 vccd1 vccd1 _5160_/D sky130_fd_sc_hd__mux2_1
Xhold506 hold506/A vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__buf_2
Xhold517 _4001_/Y vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__buf_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3432_ _5227_/Q _3596_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5227_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4432__17/A
+ sky130_fd_sc_hd__clkbuf_16
X_3363_ _3501_/A1 _5316_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5316_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5102_ _5383_/CLK _5102_/D vssd1 vssd1 vccd1 vccd1 _5102_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1206 hold1897/X vssd1 vssd1 vccd1 vccd1 hold1898/A sky130_fd_sc_hd__buf_2
X_3294_ _3325_/A _3294_/B vssd1 vssd1 vccd1 vccd1 _3294_/X sky130_fd_sc_hd__or2_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/CLK _5033_/D vssd1 vssd1 vccd1 vccd1 _5033_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1228 hold1932/X vssd1 vssd1 vccd1 vccd1 hold1933/A sky130_fd_sc_hd__buf_2
Xhold1239 hold1948/X vssd1 vssd1 vccd1 vccd1 hold1949/A sky130_fd_sc_hd__buf_2
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5866_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930__515 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5651_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput126 probe_out[91] vssd1 vssd1 vccd1 vccd1 _5928_/A sky130_fd_sc_hd__clkbuf_2
Xinput115 probe_out[81] vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__clkbuf_2
Xinput104 probe_out[71] vssd1 vssd1 vccd1 vccd1 _5908_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2430 hold2430/A vssd1 vssd1 vccd1 vccd1 hold2430/X sky130_fd_sc_hd__buf_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2441 hold2441/A vssd1 vssd1 vccd1 vccd1 hold2441/X sky130_fd_sc_hd__buf_2
Xinput137 input137/A vssd1 vssd1 vccd1 vccd1 _3672_/A sky130_fd_sc_hd__buf_6
Xhold2463 hold2463/A vssd1 vssd1 vccd1 vccd1 hold2463/X sky130_fd_sc_hd__buf_2
Xinput148 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _2492_/C sky130_fd_sc_hd__clkbuf_2
Xinput159 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _2493_/A sky130_fd_sc_hd__clkbuf_2
Xhold2452 hold48/X vssd1 vssd1 vccd1 vccd1 hold2452/X sky130_fd_sc_hd__buf_2
Xhold2485 hold2485/A vssd1 vssd1 vccd1 vccd1 hold2485/X sky130_fd_sc_hd__buf_2
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2474 hold2474/A vssd1 vssd1 vccd1 vccd1 hold810/A sky130_fd_sc_hd__buf_2
Xhold1762 hold2471/X vssd1 vssd1 vccd1 vccd1 hold2472/A sky130_fd_sc_hd__buf_2
XFILLER_57_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4494__79 _4510__95/A vssd1 vssd1 vccd1 vccd1 _5136_/CLK sky130_fd_sc_hd__inv_2
Xhold1773 hold2488/X vssd1 vssd1 vccd1 vccd1 hold2489/A sky130_fd_sc_hd__buf_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4673__258 _5007_/CLK vssd1 vssd1 vccd1 vccd1 _5361_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4714__299 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5405_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4567__152 _4508__93/A vssd1 vssd1 vccd1 vccd1 _5217_/CLK sky130_fd_sc_hd__inv_2
X_3981_ _3645_/A _5250_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _5250_/D sky130_fd_sc_hd__mux2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2932_ _3004_/C1 _2925_/X _3075_/B1 vssd1 vssd1 vccd1 vccd1 _2932_/X sky130_fd_sc_hd__a21o_1
X_5720_ _5720_/CLK _5720_/D vssd1 vssd1 vccd1 vccd1 _5720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4608__193 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5282_/CLK sky130_fd_sc_hd__inv_2
X_2863_ _2863_/A _3962_/B vssd1 vssd1 vccd1 vccd1 _2863_/Y sky130_fd_sc_hd__nor2_1
X_5651_ _5651_/CLK _5651_/D vssd1 vssd1 vccd1 vccd1 _5651_/Q sky130_fd_sc_hd__dfxtp_1
X_5582_ _5582_/CLK _5582_/D vssd1 vssd1 vccd1 vccd1 _5582_/Q sky130_fd_sc_hd__dfxtp_1
X_2794_ _3394_/A0 _5443_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5443_/D sky130_fd_sc_hd__mux2_1
XCaravelHost_721 vssd1 vssd1 vccd1 vccd1 CaravelHost_721/HI versionID[3] sky130_fd_sc_hd__conb_1
XCaravelHost_710 vssd1 vssd1 vccd1 vccd1 CaravelHost_710/HI manufacturerID[10] sky130_fd_sc_hd__conb_1
Xhold303 _3946_/X vssd1 vssd1 vccd1 vccd1 _5103_/D sky130_fd_sc_hd__buf_2
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold358 hold358/A vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__buf_2
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3415_ _5373_/Q _3453_/C _3443_/B vssd1 vssd1 vccd1 vccd1 _3589_/B sky130_fd_sc_hd__or3b_4
X_4395_ _3638_/A _4357_/B _4398_/A2 vssd1 vssd1 vccd1 vccd1 _4395_/X sky130_fd_sc_hd__a21bo_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _3346_/A _3349_/A vssd1 vssd1 vccd1 vccd1 _3347_/C sky130_fd_sc_hd__or2_1
XFILLER_140_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1014 hold1582/X vssd1 vssd1 vccd1 vccd1 hold1583/A sky130_fd_sc_hd__buf_2
Xhold1003 hold2410/X vssd1 vssd1 vccd1 vccd1 hold2411/A sky130_fd_sc_hd__buf_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 hold1592/X vssd1 vssd1 vccd1 vccd1 hold1593/A sky130_fd_sc_hd__buf_2
Xhold1058 hold1121/X vssd1 vssd1 vccd1 vccd1 hold1122/A sky130_fd_sc_hd__buf_2
X_3277_ _3277_/A1 _3159_/B _3276_/X _3277_/C1 vssd1 vssd1 vccd1 vccd1 _5339_/D sky130_fd_sc_hd__o211a_1
Xhold1047 hold149/X vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__buf_2
XFILLER_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5016_ _5016_/CLK _5016_/D vssd1 vssd1 vccd1 vccd1 _5016_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1036 hold675/X vssd1 vssd1 vccd1 vccd1 hold1643/A sky130_fd_sc_hd__buf_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1069 hold2187/X vssd1 vssd1 vccd1 vccd1 hold2188/A sky130_fd_sc_hd__buf_2
XFILLER_39_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5918_ _5918_/A vssd1 vssd1 vccd1 vccd1 _5918_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _5849_/A vssd1 vssd1 vccd1 vccd1 _5849_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2282 hold2282/A vssd1 vssd1 vccd1 vccd1 hold2282/X sky130_fd_sc_hd__buf_2
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2271 hold2271/A vssd1 vssd1 vccd1 vccd1 hold974/A sky130_fd_sc_hd__buf_2
Xhold2260 hold24/X vssd1 vssd1 vccd1 vccd1 hold2260/X sky130_fd_sc_hd__buf_2
XFILLER_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1570 hold23/X vssd1 vssd1 vccd1 vccd1 hold1570/X sky130_fd_sc_hd__buf_2
Xhold2293 hold2293/A vssd1 vssd1 vccd1 vccd1 hold980/A sky130_fd_sc_hd__buf_2
Xhold1592 _3942_/X vssd1 vssd1 vccd1 vccd1 hold1592/X sky130_fd_sc_hd__buf_2
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1581 hold1581/A vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__buf_2
XFILLER_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4180_ _3836_/A _4178_/C _4179_/X vssd1 vssd1 vccd1 vccd1 _5530_/D sky130_fd_sc_hd__a21oi_1
X_3200_ _5611_/Q _5595_/Q _5579_/Q _5619_/Q _3281_/S _3130_/B vssd1 vssd1 vccd1 vccd1
+ _3200_/X sky130_fd_sc_hd__mux4_2
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3131_ _3132_/A _3138_/B vssd1 vssd1 vccd1 vccd1 _3131_/Y sky130_fd_sc_hd__nor2_4
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3062_ _3094_/B _3051_/Y _3054_/Y _3061_/X vssd1 vssd1 vccd1 vccd1 _3077_/A sky130_fd_sc_hd__a31o_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _5376_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _5203_/D sky130_fd_sc_hd__and2_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2915_ _2863_/A _5381_/Q _3094_/A _2914_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _2915_/X
+ sky130_fd_sc_hd__a221o_1
X_3895_ _4399_/B _3893_/X hold555/X vssd1 vssd1 vccd1 vccd1 _3895_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5703_ _5703_/CLK _5703_/D vssd1 vssd1 vccd1 vccd1 _5703_/Q sky130_fd_sc_hd__dfxtp_1
X_2846_ _5398_/Q _3538_/A0 _2851_/S vssd1 vssd1 vccd1 vccd1 _5398_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5634_ _5634_/CLK _5634_/D vssd1 vssd1 vccd1 vccd1 _5634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2777_ _2777_/A _3081_/B vssd1 vssd1 vccd1 vccd1 _3091_/A sky130_fd_sc_hd__nor2_4
X_5565_ _5565_/CLK _5565_/D vssd1 vssd1 vccd1 vccd1 _5565_/Q sky130_fd_sc_hd__dfxtp_1
Xhold100 hold73/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__buf_2
XFILLER_144_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold111 hold122/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__buf_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__buf_2
X_5496_ _5496_/CLK _5496_/D vssd1 vssd1 vccd1 vccd1 _5496_/Q sky130_fd_sc_hd__dfxtp_1
Xhold144 hold172/X vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__buf_2
X_4695__280 _4941__526/A vssd1 vssd1 vccd1 vccd1 _5386_/CLK sky130_fd_sc_hd__inv_2
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__buf_2
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__buf_2
Xhold155 hold169/X vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__buf_2
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__buf_2
XFILLER_144_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout613 _5321_/Q vssd1 vssd1 vccd1 vccd1 _2848_/A1 sky130_fd_sc_hd__buf_2
XFILLER_113_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout624 _3543_/A0 vssd1 vssd1 vccd1 vccd1 _3606_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout602 _5323_/Q vssd1 vssd1 vccd1 vccd1 _3592_/A1 sky130_fd_sc_hd__buf_4
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__buf_2
Xhold188 hold294/X vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__buf_2
XFILLER_144_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4378_ _5738_/Q _4370_/X _4378_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4378_/X sky130_fd_sc_hd__o211a_1
Xfanout646 _4390_/A vssd1 vssd1 vccd1 vccd1 hold599/A sky130_fd_sc_hd__buf_2
Xfanout635 _3824_/A1 vssd1 vssd1 vccd1 vccd1 _3718_/A1 sky130_fd_sc_hd__buf_6
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _5417_/Q _2482_/B _3237_/B _5409_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _3329_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4464__49 _4424__9/A vssd1 vssd1 vccd1 vccd1 _5058_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4936__521 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5657_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2090 hold441/X vssd1 vssd1 vccd1 vccd1 hold2090/X sky130_fd_sc_hd__buf_2
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2700_ _5523_/Q _3568_/A1 _2702_/S vssd1 vssd1 vccd1 vccd1 _5523_/D sky130_fd_sc_hd__mux2_1
X_3680_ _5253_/Q _3682_/B vssd1 vssd1 vccd1 vccd1 _3680_/X sky130_fd_sc_hd__and2_1
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4679__264 _4432__17/A vssd1 vssd1 vccd1 vccd1 _5368_/CLK sky130_fd_sc_hd__inv_2
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2631_ _2617_/X _2621_/X _2627_/X _2630_/X vssd1 vssd1 vccd1 vccd1 _4358_/B sky130_fd_sc_hd__a211o_4
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput216 _3679_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5350_ _5350_/CLK _5350_/D vssd1 vssd1 vccd1 vccd1 _5350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2562_ _3576_/A0 _5650_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5650_/D sky130_fd_sc_hd__mux2_1
Xoutput249 _3650_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__clkbuf_2
Xoutput238 _3640_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput227 _3663_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4301_ _4300_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5670_/D sky130_fd_sc_hd__and2b_1
X_5281_ _5281_/CLK _5281_/D vssd1 vssd1 vccd1 vccd1 _5281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4232_ _5560_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__or2_1
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2493_ _2493_/A _2493_/B input167/X vssd1 vssd1 vccd1 vccd1 _2496_/A sky130_fd_sc_hd__or3b_4
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4163_ _5738_/Q _4186_/A vssd1 vssd1 vccd1 vccd1 _4164_/B sky130_fd_sc_hd__nand2_8
X_3114_ _3590_/A1 _5354_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5354_/D sky130_fd_sc_hd__mux2_1
X_4094_ _5738_/Q _5309_/Q _4094_/C vssd1 vssd1 vccd1 vccd1 _4094_/X sky130_fd_sc_hd__and3_1
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3045_ _3045_/A1 _3026_/X _3029_/X _3044_/X _2883_/X vssd1 vssd1 vccd1 vccd1 _3045_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _5551_/CLK _4996_/D vssd1 vssd1 vccd1 vccd1 _4996_/Q sky130_fd_sc_hd__dfxtp_1
X_3947_ _5251_/Q _5104_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _5104_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3878_ _5733_/Q _3857_/Y _3877_/X _3887_/B _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3878_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2829_ _3392_/A0 _5413_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5413_/D sky130_fd_sc_hd__mux2_1
X_5617_ _5617_/CLK _5617_/D vssd1 vssd1 vccd1 vccd1 _5617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5548_ _5551_/CLK _5548_/D vssd1 vssd1 vccd1 vccd1 _5548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4509__94 _4509__94/A vssd1 vssd1 vccd1 vccd1 _5151_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5479_ _5479_/CLK _5479_/D vssd1 vssd1 vccd1 vccd1 _5479_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout432 _3621_/X vssd1 vssd1 vccd1 vccd1 _3642_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout421 hold506/A vssd1 vssd1 vccd1 vccd1 hold483/A sky130_fd_sc_hd__buf_4
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout410 _4182_/X vssd1 vssd1 vccd1 vccd1 _4209_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout454 _2875_/X vssd1 vssd1 vccd1 vccd1 _2919_/B sky130_fd_sc_hd__buf_8
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout443 _4409_/B vssd1 vssd1 vccd1 vccd1 _4415_/A3 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout465 _3282_/C1 vssd1 vssd1 vccd1 vccd1 _3240_/S sky130_fd_sc_hd__clkbuf_8
Xfanout498 _2866_/B vssd1 vssd1 vccd1 vccd1 _3041_/A2 sky130_fd_sc_hd__buf_6
Xfanout476 _3064_/C1 vssd1 vssd1 vccd1 vccd1 _2947_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout487 _2498_/X vssd1 vssd1 vccd1 vccd1 _4389_/B sky130_fd_sc_hd__buf_6
XFILLER_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_66_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3801_ hold277/X _5252_/Q _3810_/A3 hold349/X _5001_/Q vssd1 vssd1 vccd1 vccd1 _5001_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3732_ _4997_/Q _3732_/B vssd1 vssd1 vccd1 vccd1 _3732_/X sky130_fd_sc_hd__or2_1
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3663_ _3663_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3663_/X sky130_fd_sc_hd__and2_1
X_5402_ _5402_/CLK _5402_/D vssd1 vssd1 vccd1 vccd1 _5402_/Q sky130_fd_sc_hd__dfxtp_1
X_2614_ _5373_/Q _2625_/A _3453_/C vssd1 vssd1 vccd1 vccd1 _2779_/A sky130_fd_sc_hd__nand3_4
XFILLER_133_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3594_ _5029_/Q _3594_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5029_/D sky130_fd_sc_hd__mux2_1
X_5333_ _5333_/CLK _5333_/D vssd1 vssd1 vccd1 vccd1 _5333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2545_ _2545_/A _3350_/B vssd1 vssd1 vccd1 vccd1 _3349_/A sky130_fd_sc_hd__nor2_8
XFILLER_130_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5264_ _5265_/CLK _5264_/D vssd1 vssd1 vccd1 vccd1 _5264_/Q sky130_fd_sc_hd__dfxtp_1
X_2476_ _3122_/B _3122_/A _3123_/A vssd1 vssd1 vccd1 vccd1 _2487_/A sky130_fd_sc_hd__mux2_1
Xhold2804 hold2804/A vssd1 vssd1 vccd1 vccd1 hold2804/X sky130_fd_sc_hd__buf_2
X_5195_ _5195_/CLK _5195_/D vssd1 vssd1 vccd1 vccd1 _5195_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2826 hold2826/A vssd1 vssd1 vccd1 vccd1 hold2826/X sky130_fd_sc_hd__buf_2
X_4215_ _4217_/A _4215_/B vssd1 vssd1 vccd1 vccd1 _5553_/D sky130_fd_sc_hd__nor2_1
X_4146_ _4130_/A _4130_/B _5750_/Q vssd1 vssd1 vccd1 vccd1 _4171_/C sky130_fd_sc_hd__a21bo_1
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4077_ _5663_/Q _5664_/Q vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__nand2b_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _4976_/Q _2868_/Y _3027_/X _3034_/A vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__o22a_1
X_4434__19 _4439__24/A vssd1 vssd1 vccd1 vccd1 _5028_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4979_ _4979_/CLK _4979_/D vssd1 vssd1 vccd1 vccd1 _4979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4731__316/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4000_ _3980_/A _5292_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__mux2_1
XFILLER_84_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4841__426 _5001_/CLK vssd1 vssd1 vccd1 vccd1 _5534_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5882_ _5882_/A vssd1 vssd1 vccd1 vccd1 _5882_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3715_ _3718_/A1 _3713_/X _3714_/X split2/X vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__o211a_1
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3646_ _3646_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__or2_1
X_4735__320 _4744__329/A vssd1 vssd1 vccd1 vccd1 _5426_/CLK sky130_fd_sc_hd__inv_2
X_3577_ _3577_/A0 _5044_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5044_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5316_ _5316_/CLK _5316_/D vssd1 vssd1 vccd1 vccd1 _5316_/Q sky130_fd_sc_hd__dfxtp_1
X_2528_ _3391_/A0 _5713_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5713_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5247_ _5247_/CLK _5247_/D vssd1 vssd1 vccd1 vccd1 _5247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2459_ _5369_/Q vssd1 vssd1 vccd1 vccd1 _2776_/A sky130_fd_sc_hd__inv_2
Xhold1900 hold1900/A vssd1 vssd1 vccd1 vccd1 _5742_/D sky130_fd_sc_hd__buf_2
Xhold2656 hold2656/A vssd1 vssd1 vccd1 vccd1 hold2656/X sky130_fd_sc_hd__buf_2
Xhold1911 hold1911/A vssd1 vssd1 vccd1 vccd1 _5744_/D sky130_fd_sc_hd__buf_2
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__buf_2
Xhold2645 hold243/X vssd1 vssd1 vccd1 vccd1 hold2645/X sky130_fd_sc_hd__buf_2
Xhold2634 hold2634/A vssd1 vssd1 vccd1 vccd1 hold2634/X sky130_fd_sc_hd__buf_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__buf_2
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__buf_2
X_5178_ _5178_/CLK _5178_/D vssd1 vssd1 vccd1 vccd1 _5178_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1933 hold1933/A vssd1 vssd1 vccd1 vccd1 _5737_/D sky130_fd_sc_hd__buf_2
XFILLER_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1922 hold1922/A vssd1 vssd1 vccd1 vccd1 _5741_/D sky130_fd_sc_hd__buf_2
Xhold1944 hold1944/A vssd1 vssd1 vccd1 vccd1 _5740_/D sky130_fd_sc_hd__buf_2
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__buf_2
Xhold2689 hold2689/A vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__buf_2
Xhold2678 _3792_/X vssd1 vssd1 vccd1 vccd1 hold2678/X sky130_fd_sc_hd__buf_2
Xhold2667 hold2667/A vssd1 vssd1 vccd1 vccd1 hold2667/X sky130_fd_sc_hd__buf_2
XFILLER_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__buf_2
Xhold1955 hold1955/A vssd1 vssd1 vccd1 vccd1 _5736_/D sky130_fd_sc_hd__buf_2
Xhold1966 hold182/X vssd1 vssd1 vccd1 vccd1 hold1966/X sky130_fd_sc_hd__buf_2
X_4129_ _5543_/Q _4132_/B _5544_/Q vssd1 vssd1 vccd1 vccd1 _4130_/B sky130_fd_sc_hd__a21o_1
Xhold1988 hold2621/X vssd1 vssd1 vccd1 vccd1 hold2622/A sky130_fd_sc_hd__buf_2
Xhold1977 hold2608/X vssd1 vssd1 vccd1 vccd1 hold2609/A sky130_fd_sc_hd__buf_2
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1999 hold2635/X vssd1 vssd1 vccd1 vccd1 hold2636/A sky130_fd_sc_hd__buf_2
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4584__169 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5234_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3500_ _5161_/Q _3599_/A1 _3507_/S vssd1 vssd1 vccd1 vccd1 _5161_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4719__304 _4941__526/A vssd1 vssd1 vccd1 vccd1 _5410_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3431_ _5228_/Q _3595_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5228_/D sky130_fd_sc_hd__mux2_1
X_3362_ _3536_/A0 _5317_/Q _3369_/S vssd1 vssd1 vccd1 vccd1 _5317_/D sky130_fd_sc_hd__mux2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5101_ _5383_/CLK _5101_/D vssd1 vssd1 vccd1 vccd1 _5101_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1207 hold1899/X vssd1 vssd1 vccd1 vccd1 hold1900/A sky130_fd_sc_hd__buf_2
X_3293_ _5522_/Q _5275_/Q _3324_/S vssd1 vssd1 vccd1 vccd1 _3294_/B sky130_fd_sc_hd__mux2_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5032_ _5032_/CLK _5032_/D vssd1 vssd1 vccd1 vccd1 _5032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1218 hold1882/X vssd1 vssd1 vccd1 vccd1 hold1883/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_81_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4964__549/A sky130_fd_sc_hd__clkbuf_16
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5542_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5934_ _5934_/A vssd1 vssd1 vccd1 vccd1 _5934_/X sky130_fd_sc_hd__clkbuf_4
X_5865_ _5865_/A vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3629_ _4350_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3629_/X sky130_fd_sc_hd__or2_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput127 probe_out[92] vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__clkbuf_2
Xinput116 probe_out[82] vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__clkbuf_2
Xinput105 probe_out[72] vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__clkbuf_2
Xhold2431 hold2431/A vssd1 vssd1 vccd1 vccd1 hold2431/X sky130_fd_sc_hd__buf_2
Xhold2420 hold2420/A vssd1 vssd1 vccd1 vccd1 hold997/A sky130_fd_sc_hd__buf_2
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2464 hold2464/A vssd1 vssd1 vccd1 vccd1 input140/A sky130_fd_sc_hd__buf_2
Xhold2442 hold2442/A vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__buf_2
Xhold2453 hold2453/A vssd1 vssd1 vccd1 vccd1 hold2453/X sky130_fd_sc_hd__buf_2
Xinput138 input138/A vssd1 vssd1 vccd1 vccd1 _3673_/A sky130_fd_sc_hd__buf_4
Xinput149 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _2495_/B sky130_fd_sc_hd__clkbuf_2
Xhold2486 hold2486/A vssd1 vssd1 vccd1 vccd1 hold2486/X sky130_fd_sc_hd__buf_2
Xhold2497 hold2850/X vssd1 vssd1 vccd1 vccd1 hold2497/X sky130_fd_sc_hd__buf_2
Xhold2475 hold810/X vssd1 vssd1 vccd1 vccd1 hold2475/X sky130_fd_sc_hd__buf_2
XFILLER_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1730 hold2407/X vssd1 vssd1 vccd1 vccd1 hold2408/A sky130_fd_sc_hd__buf_2
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1763 hold2473/X vssd1 vssd1 vccd1 vccd1 hold2474/A sky130_fd_sc_hd__buf_2
Xhold1774 hold2490/X vssd1 vssd1 vccd1 vccd1 hold2491/A sky130_fd_sc_hd__buf_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3980_ _3980_/A _3989_/B vssd1 vssd1 vccd1 vccd1 _3980_/Y sky130_fd_sc_hd__nand2_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _3029_/B1 _2921_/X _2930_/X vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5650_ _5650_/CLK _5650_/D vssd1 vssd1 vccd1 vccd1 _5650_/Q sky130_fd_sc_hd__dfxtp_1
X_2862_ _2862_/A _2862_/B _2862_/C _2862_/D vssd1 vssd1 vccd1 vccd1 _3962_/B sky130_fd_sc_hd__and4_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5581_ _5581_/CLK _5581_/D vssd1 vssd1 vccd1 vccd1 _5581_/Q sky130_fd_sc_hd__dfxtp_1
X_2793_ _3393_/A0 _5444_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5444_/D sky130_fd_sc_hd__mux2_1
XCaravelHost_711 vssd1 vssd1 vccd1 vccd1 CaravelHost_711/HI partID[1] sky130_fd_sc_hd__conb_1
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_722 vssd1 vssd1 vccd1 vccd1 core1Index[0] CaravelHost_722/LO sky130_fd_sc_hd__conb_1
X_4953__538 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5711_/CLK sky130_fd_sc_hd__inv_2
XCaravelHost_700 vssd1 vssd1 vccd1 vccd1 CaravelHost_700/HI manufacturerID[0] sky130_fd_sc_hd__conb_1
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold359 _3813_/X vssd1 vssd1 vccd1 vccd1 _5013_/D sky130_fd_sc_hd__buf_2
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold348 hold372/X vssd1 vssd1 vccd1 vccd1 hold364/A sky130_fd_sc_hd__buf_2
X_3414_ _5266_/Q _3579_/A0 _3414_/S vssd1 vssd1 vccd1 vccd1 _5266_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4394_ _5745_/Q _4398_/A2 _4394_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4394_/X sky130_fd_sc_hd__o211a_1
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3344_/A _3347_/B _3344_/Y split3/X vssd1 vssd1 vccd1 vccd1 _5334_/D sky130_fd_sc_hd__o211a_1
X_3276_ _5339_/Q _3125_/A _3156_/X _3275_/X vssd1 vssd1 vccd1 vccd1 _3276_/X sky130_fd_sc_hd__a211o_1
Xhold1004 hold2414/X vssd1 vssd1 vccd1 vccd1 hold2415/A sky130_fd_sc_hd__buf_2
Xhold1015 hold2458/X vssd1 vssd1 vccd1 vccd1 hold2459/A sky130_fd_sc_hd__buf_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4847__432 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5568_/CLK sky130_fd_sc_hd__inv_2
Xhold1026 hold1594/X vssd1 vssd1 vccd1 vccd1 hold1595/A sky130_fd_sc_hd__buf_2
Xhold1037 hold2591/X vssd1 vssd1 vccd1 vccd1 hold2592/A sky130_fd_sc_hd__buf_2
Xhold1048 hold197/X vssd1 vssd1 vccd1 vccd1 _3827_/C sky130_fd_sc_hd__buf_2
X_5015_ _5016_/CLK _5015_/D vssd1 vssd1 vccd1 vccd1 _5015_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1059 _3955_/Y vssd1 vssd1 vccd1 vccd1 _3958_/A2 sky130_fd_sc_hd__buf_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5917_ _5917_/A vssd1 vssd1 vccd1 vccd1 _5917_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5848_ _5848_/A vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2261 hold2261/A vssd1 vssd1 vccd1 vccd1 hold968/A sky130_fd_sc_hd__buf_2
Xhold2250 hold2250/A vssd1 vssd1 vccd1 vccd1 hold962/A sky130_fd_sc_hd__buf_2
Xhold2272 hold974/X vssd1 vssd1 vccd1 vccd1 hold2272/X sky130_fd_sc_hd__buf_2
Xhold2283 hold2283/A vssd1 vssd1 vccd1 vccd1 hold662/A sky130_fd_sc_hd__buf_2
Xhold1571 hold1571/A vssd1 vssd1 vccd1 vccd1 _5089_/D sky130_fd_sc_hd__buf_2
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1560 hold2409/X vssd1 vssd1 vccd1 vccd1 hold2410/A sky130_fd_sc_hd__buf_2
Xhold2294 hold980/X vssd1 vssd1 vccd1 vccd1 hold2294/X sky130_fd_sc_hd__buf_2
Xhold1593 hold1593/A vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__buf_2
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1582 hold41/X vssd1 vssd1 vccd1 vccd1 hold1582/X sky130_fd_sc_hd__buf_2
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4640__225 _4921__506/A vssd1 vssd1 vccd1 vccd1 _5326_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3130_ _5328_/Q _3130_/B _3281_/S vssd1 vssd1 vccd1 vccd1 _3138_/B sky130_fd_sc_hd__and3_2
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3061_ _2883_/X _3057_/Y _3060_/Y _3043_/A vssd1 vssd1 vccd1 vccd1 _3061_/X sky130_fd_sc_hd__a31o_1
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ _5375_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _5202_/D sky130_fd_sc_hd__and2_1
X_2914_ _2883_/X _2909_/X _2913_/X _2905_/X vssd1 vssd1 vccd1 vccd1 _2914_/X sky130_fd_sc_hd__a31o_2
X_3894_ _3844_/A _3955_/A _5073_/Q hold554/X vssd1 vssd1 vccd1 vccd1 _3894_/X sky130_fd_sc_hd__a31o_1
X_5702_ _5702_/CLK _5702_/D vssd1 vssd1 vccd1 vccd1 _5702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2845_ _5399_/Q _3501_/A1 _2851_/S vssd1 vssd1 vccd1 vccd1 _5399_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5633_ _5633_/CLK _5633_/D vssd1 vssd1 vccd1 vccd1 _5633_/Q sky130_fd_sc_hd__dfxtp_1
X_5564_ _5564_/CLK _5564_/D vssd1 vssd1 vccd1 vccd1 _5564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2776_ _2776_/A _3081_/B vssd1 vssd1 vccd1 vccd1 _3093_/A sky130_fd_sc_hd__nor2_1
Xhold101 hold74/X vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__buf_2
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold134 _3980_/Y vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__buf_2
XFILLER_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__buf_2
X_5495_ _5495_/CLK _5495_/D vssd1 vssd1 vccd1 vccd1 _5495_/Q sky130_fd_sc_hd__dfxtp_1
Xhold112 hold124/X vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__buf_2
XFILLER_144_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold145 hold176/X vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__buf_2
Xhold167 hold33/X vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__buf_2
Xhold156 hold171/X vssd1 vssd1 vccd1 vccd1 hold172/A sky130_fd_sc_hd__buf_2
Xfanout603 _5323_/Q vssd1 vssd1 vccd1 vccd1 _3610_/A1 sky130_fd_sc_hd__buf_2
Xfanout614 _5320_/Q vssd1 vssd1 vccd1 vccd1 _3595_/A1 sky130_fd_sc_hd__buf_4
X_4377_ _3646_/A _4389_/B _4370_/X vssd1 vssd1 vccd1 vccd1 _4377_/X sky130_fd_sc_hd__a21bo_1
XFILLER_59_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__buf_2
Xhold189 hold296/X vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__buf_2
XFILLER_113_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout625 _5318_/Q vssd1 vssd1 vccd1 vccd1 _3543_/A0 sky130_fd_sc_hd__buf_4
XFILLER_98_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout647 _4360_/A vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__buf_6
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3328_/A _3328_/B vssd1 vssd1 vccd1 vccd1 _3328_/X sky130_fd_sc_hd__or2_1
Xfanout636 _3824_/A1 vssd1 vssd1 vccd1 vccd1 _3733_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3259_ _5268_/Q _5295_/Q _3290_/S vssd1 vssd1 vccd1 vccd1 _3259_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4624__209 _4456__41/A vssd1 vssd1 vccd1 vccd1 _5301_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4518__103 _5007_/CLK vssd1 vssd1 vccd1 vccd1 _5160_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold690 hold690/A vssd1 vssd1 vccd1 vccd1 _4357_/B sky130_fd_sc_hd__buf_2
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2091 hold2091/A vssd1 vssd1 vccd1 vccd1 _4989_/D sky130_fd_sc_hd__buf_2
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _2861_/A _2777_/A _3081_/A _2861_/B _2862_/C vssd1 vssd1 vccd1 vccd1 _2630_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput206 _5025_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__clkbuf_2
Xoutput217 _3680_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2561_ _3575_/A0 _5651_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5651_/D sky130_fd_sc_hd__mux2_1
Xoutput239 _3641_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput228 _3664_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4300_ _4048_/Y _4308_/A2 _4308_/B1 _2448_/Y vssd1 vssd1 vccd1 vccd1 _4300_/X sky130_fd_sc_hd__o22a_1
X_5280_ _5280_/CLK _5280_/D vssd1 vssd1 vccd1 vccd1 _5280_/Q sky130_fd_sc_hd__dfxtp_1
X_2492_ _2492_/A _2492_/B _2492_/C _2492_/D vssd1 vssd1 vccd1 vccd1 _2497_/C sky130_fd_sc_hd__or4_2
XFILLER_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _5338_/Q _4360_/B _4164_/B _4230_/X _4244_/S vssd1 vssd1 vccd1 vccd1 _5559_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _4177_/B _4170_/A _4162_/C _4162_/D vssd1 vssd1 vccd1 vccd1 _4186_/B sky130_fd_sc_hd__and4_4
X_3113_ _3508_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3121_/S sky130_fd_sc_hd__or2_4
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4093_ _5566_/Q _4093_/B _4093_/C _5738_/Q vssd1 vssd1 vccd1 vccd1 _4093_/X sky130_fd_sc_hd__and4b_1
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3044_ _3034_/X _3035_/X _3075_/B1 _3032_/X vssd1 vssd1 vccd1 vccd1 _3044_/X sky130_fd_sc_hd__a211o_1
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4995_ _5246_/CLK _4995_/D vssd1 vssd1 vccd1 vccd1 _4995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3946_ _5250_/Q _5103_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _3946_/X sky130_fd_sc_hd__mux2_1
X_4959__544 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5717_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3877_ _3998_/A1 _5206_/Q _3882_/A3 _3855_/X vssd1 vssd1 vccd1 vccd1 _3877_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5616_ _5616_/CLK _5616_/D vssd1 vssd1 vccd1 vccd1 _5616_/Q sky130_fd_sc_hd__dfxtp_1
X_2828_ _3391_/A0 _5414_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5414_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5547_ _5551_/CLK _5547_/D vssd1 vssd1 vccd1 vccd1 _5547_/Q sky130_fd_sc_hd__dfxtp_1
X_2759_ _3389_/A0 _5472_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5472_/D sky130_fd_sc_hd__mux2_1
X_5478_ _5478_/CLK _5478_/D vssd1 vssd1 vccd1 vccd1 _5478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout422 _4000_/S vssd1 vssd1 vccd1 vccd1 _3999_/S sky130_fd_sc_hd__buf_8
Xfanout411 _3901_/X vssd1 vssd1 vccd1 vccd1 _3921_/C1 sky130_fd_sc_hd__buf_6
Xfanout433 _3660_/B vssd1 vssd1 vccd1 vccd1 _3659_/B sky130_fd_sc_hd__clkbuf_4
Xfanout455 _2875_/X vssd1 vssd1 vccd1 vccd1 _3075_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout444 _4381_/X vssd1 vssd1 vccd1 vccd1 _4398_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout466 _3131_/Y vssd1 vssd1 vccd1 vccd1 _3282_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout499 _3031_/B1 vssd1 vssd1 vccd1 vccd1 _2866_/B sky130_fd_sc_hd__buf_6
Xfanout477 _3004_/C1 vssd1 vssd1 vccd1 vccd1 _3064_/C1 sky130_fd_sc_hd__buf_4
Xfanout488 _2498_/X vssd1 vssd1 vccd1 vccd1 _3778_/B sky130_fd_sc_hd__buf_2
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4752__337 _5734_/CLK vssd1 vssd1 vccd1 vccd1 _5443_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4646__231 _5553_/CLK vssd1 vssd1 vccd1 vccd1 _5332_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3800_ hold277/X _5251_/Q _3810_/A3 hold349/X _5000_/Q vssd1 vssd1 vccd1 vccd1 _5000_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _5080_/Q input8/X _3763_/B vssd1 vssd1 vccd1 vccd1 _3731_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4419__4/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _3662_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3662_/X sky130_fd_sc_hd__and2_1
XFILLER_119_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5401_ _5401_/CLK _5401_/D vssd1 vssd1 vccd1 vccd1 _5401_/Q sky130_fd_sc_hd__dfxtp_1
X_3593_ _5030_/Q _3593_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5030_/D sky130_fd_sc_hd__mux2_1
X_2613_ _3339_/A1 _5607_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5607_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5332_ _5332_/CLK _5332_/D vssd1 vssd1 vccd1 vccd1 _5332_/Q sky130_fd_sc_hd__dfxtp_4
X_2544_ _5335_/Q _3344_/A _5333_/Q vssd1 vssd1 vccd1 vccd1 _2852_/A sky130_fd_sc_hd__or3b_4
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5263_ _5265_/CLK _5263_/D vssd1 vssd1 vccd1 vccd1 _5263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2475_ _3350_/A _3312_/S vssd1 vssd1 vccd1 vccd1 _3122_/B sky130_fd_sc_hd__nand2_1
Xhold2805 hold2805/A vssd1 vssd1 vccd1 vccd1 hold2805/X sky130_fd_sc_hd__buf_2
X_5194_ _5194_/CLK _5194_/D vssd1 vssd1 vccd1 vccd1 _5194_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2838 _4084_/X vssd1 vssd1 vccd1 vccd1 hold2838/X sky130_fd_sc_hd__buf_2
X_4214_ _5553_/Q _4209_/B _4210_/C _4151_/Y vssd1 vssd1 vccd1 vccd1 _4215_/B sky130_fd_sc_hd__o2bb2a_1
X_4145_ _4145_/A _4171_/B _4145_/C vssd1 vssd1 vccd1 vccd1 _4149_/C sky130_fd_sc_hd__and3_1
XFILLER_29_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4076_ _5663_/Q _5664_/Q vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__and2b_1
X_3027_ _5035_/Q _5532_/Q _3072_/S vssd1 vssd1 vccd1 vccd1 _3027_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _4978_/CLK _4978_/D vssd1 vssd1 vccd1 vccd1 _4978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3929_ _3959_/A _3959_/B _3960_/A _5088_/Q hold711/A vssd1 vssd1 vccd1 vccd1 _3929_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4880__465 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5881_ _5881_/A vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3714_ _4991_/Q _3729_/B vssd1 vssd1 vccd1 vccd1 _3714_/X sky130_fd_sc_hd__or2_1
XFILLER_146_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3645_ _3645_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3645_/X sky130_fd_sc_hd__or2_1
XFILLER_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3576_ _3576_/A0 _5045_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5045_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5315_ _5315_/CLK _5315_/D vssd1 vssd1 vccd1 vccd1 _5315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2527_ _3390_/A0 _5714_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5714_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2458_ _3443_/B vssd1 vssd1 vccd1 vccd1 _2625_/A sky130_fd_sc_hd__clkinv_2
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5246_ _5246_/CLK _5246_/D vssd1 vssd1 vccd1 vccd1 _5246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__buf_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__buf_2
Xhold2646 hold2646/A vssd1 vssd1 vccd1 vccd1 hold2646/X sky130_fd_sc_hd__buf_2
Xhold2635 hold2635/A vssd1 vssd1 vccd1 vccd1 hold2635/X sky130_fd_sc_hd__buf_2
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__buf_2
XFILLER_96_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5177_ _5177_/CLK _5177_/D vssd1 vssd1 vccd1 vccd1 _5177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2657 hold2657/A vssd1 vssd1 vccd1 vccd1 hold682/A sky130_fd_sc_hd__buf_2
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__buf_2
Xhold2679 hold2679/A vssd1 vssd1 vccd1 vccd1 hold2679/X sky130_fd_sc_hd__buf_2
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1967 hold1967/A vssd1 vssd1 vccd1 vccd1 _5111_/D sky130_fd_sc_hd__buf_2
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _5749_/Q _4128_/B _4128_/C vssd1 vssd1 vccd1 vccd1 _4171_/A sky130_fd_sc_hd__nand3b_1
Xhold1978 hold1978/A vssd1 vssd1 vccd1 vccd1 _5699_/D sky130_fd_sc_hd__buf_2
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4059_ _5753_/Q _4259_/B _4259_/C vssd1 vssd1 vccd1 vccd1 _4059_/X sky130_fd_sc_hd__and3_1
Xhold1989 hold1989/A vssd1 vssd1 vccd1 vccd1 _5698_/D sky130_fd_sc_hd__buf_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4864__449 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5585_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758__343 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5449_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3430_ _5229_/Q _3594_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5229_/D sky130_fd_sc_hd__mux2_1
X_3361_ _3508_/A _3535_/B vssd1 vssd1 vccd1 vccd1 _3369_/S sky130_fd_sc_hd__or2_4
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5100_ _5383_/CLK _5100_/D vssd1 vssd1 vccd1 vccd1 _5100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5031_ _5031_/CLK _5031_/D vssd1 vssd1 vccd1 vccd1 _5031_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3357_/B _3290_/X _3291_/X _3323_/C1 vssd1 vssd1 vccd1 vccd1 _3292_/X sky130_fd_sc_hd__o211a_1
Xhold1219 hold1884/X vssd1 vssd1 vccd1 vccd1 hold1885/A sky130_fd_sc_hd__buf_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5933_ _5933_/A vssd1 vssd1 vccd1 vccd1 _5933_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_50_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5002_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5864_ _5864_/A vssd1 vssd1 vccd1 vccd1 _5864_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3628_ _3628_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3628_/X sky130_fd_sc_hd__and2_1
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3559_ _5060_/Q _3604_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5060_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4551__136 _4423__8/A vssd1 vssd1 vccd1 vccd1 _5193_/CLK sky130_fd_sc_hd__inv_2
Xinput117 probe_out[83] vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__clkbuf_2
Xinput106 probe_out[73] vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__clkbuf_2
Xhold2410 hold2410/A vssd1 vssd1 vccd1 vccd1 hold2410/X sky130_fd_sc_hd__buf_2
Xhold2421 hold997/X vssd1 vssd1 vccd1 vccd1 hold2421/X sky130_fd_sc_hd__buf_2
Xinput128 probe_out[93] vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__clkbuf_2
X_5229_ _5229_/CLK _5229_/D vssd1 vssd1 vccd1 vccd1 _5229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1720 hold2382/X vssd1 vssd1 vccd1 vccd1 hold2383/A sky130_fd_sc_hd__buf_2
Xhold2443 hold45/X vssd1 vssd1 vccd1 vccd1 hold2443/X sky130_fd_sc_hd__buf_2
Xhold2454 hold2454/A vssd1 vssd1 vccd1 vccd1 hold2454/X sky130_fd_sc_hd__buf_2
Xinput139 input139/A vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__buf_4
Xhold2432 hold2432/A vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__buf_2
Xhold2476 hold2476/A vssd1 vssd1 vccd1 vccd1 hold2476/X sky130_fd_sc_hd__buf_2
Xhold2498 hold2498/A vssd1 vssd1 vccd1 vccd1 hold2498/X sky130_fd_sc_hd__buf_2
Xhold2487 hold2487/A vssd1 vssd1 vccd1 vccd1 hold793/A sky130_fd_sc_hd__buf_2
Xhold1753 hold2562/X vssd1 vssd1 vccd1 vccd1 hold2563/A sky130_fd_sc_hd__buf_2
Xhold2465 _3675_/A vssd1 vssd1 vccd1 vccd1 hold2465/X sky130_fd_sc_hd__buf_2
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1764 hold2475/X vssd1 vssd1 vccd1 vccd1 hold2476/A sky130_fd_sc_hd__buf_2
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2930_ _3073_/C1 _2920_/X _3045_/A1 vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4423__8 _4423__8/A vssd1 vssd1 vccd1 vccd1 _4974_/CLK sky130_fd_sc_hd__inv_2
X_2861_ _2861_/A _2861_/B vssd1 vssd1 vccd1 vccd1 _2862_/D sky130_fd_sc_hd__nor2_1
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5580_ _5580_/CLK _5580_/D vssd1 vssd1 vccd1 vccd1 _5580_/Q sky130_fd_sc_hd__dfxtp_1
X_2792_ _3392_/A0 _5445_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5445_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XCaravelHost_712 vssd1 vssd1 vccd1 vccd1 CaravelHost_712/HI partID[3] sky130_fd_sc_hd__conb_1
XCaravelHost_701 vssd1 vssd1 vccd1 vccd1 CaravelHost_701/HI manufacturerID[1] sky130_fd_sc_hd__conb_1
XCaravelHost_723 vssd1 vssd1 vccd1 vccd1 partID[0] CaravelHost_723/LO sky130_fd_sc_hd__conb_1
Xhold316 hold327/X vssd1 vssd1 vccd1 vccd1 hold328/A sky130_fd_sc_hd__buf_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold349 hold349/A vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__buf_2
Xhold327 hold327/A vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__buf_2
X_3413_ _5267_/Q _3578_/A0 _3414_/S vssd1 vssd1 vccd1 vccd1 _5267_/D sky130_fd_sc_hd__mux2_1
X_4393_ _3639_/A _4389_/B _4398_/A2 vssd1 vssd1 vccd1 vccd1 _4393_/X sky130_fd_sc_hd__a21bo_1
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3344_/A _3347_/B vssd1 vssd1 vccd1 vccd1 _3344_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1005 hold2418/X vssd1 vssd1 vccd1 vccd1 hold1565/A sky130_fd_sc_hd__buf_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3272_/X _3274_/X _3357_/A vssd1 vssd1 vccd1 vccd1 _3275_/X sky130_fd_sc_hd__o21a_1
X_5014_ _5265_/CLK _5014_/D vssd1 vssd1 vccd1 vccd1 _5014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1038 hold2595/X vssd1 vssd1 vccd1 vccd1 hold2596/A sky130_fd_sc_hd__buf_2
Xhold1049 _3827_/X vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__buf_2
Xhold1027 hold2449/X vssd1 vssd1 vccd1 vccd1 hold2450/A sky130_fd_sc_hd__buf_2
Xhold1016 hold2462/X vssd1 vssd1 vccd1 vccd1 hold2463/A sky130_fd_sc_hd__buf_2
X_4886__471 _4897__482/A vssd1 vssd1 vccd1 vccd1 _5607_/CLK sky130_fd_sc_hd__inv_2
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5916_ _5916_/A vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5847_ _5847_/A vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold872 hold879/X vssd1 vssd1 vccd1 vccd1 hold872/X sky130_fd_sc_hd__buf_2
XFILLER_89_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2240 hold956/X vssd1 vssd1 vccd1 vccd1 hold2240/X sky130_fd_sc_hd__buf_2
Xhold2251 hold962/X vssd1 vssd1 vccd1 vccd1 hold2251/X sky130_fd_sc_hd__buf_2
Xhold2262 hold968/X vssd1 vssd1 vccd1 vccd1 hold2262/X sky130_fd_sc_hd__buf_2
Xhold2273 hold2273/A vssd1 vssd1 vccd1 vccd1 input164/A sky130_fd_sc_hd__buf_2
Xhold2284 hold662/X vssd1 vssd1 vccd1 vccd1 hold2284/X sky130_fd_sc_hd__buf_2
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1550 hold2423/X vssd1 vssd1 vccd1 vccd1 hold2424/A sky130_fd_sc_hd__buf_2
Xhold1561 hold2411/X vssd1 vssd1 vccd1 vccd1 hold2412/A sky130_fd_sc_hd__buf_2
Xhold2295 hold2295/A vssd1 vssd1 vccd1 vccd1 input165/A sky130_fd_sc_hd__buf_2
Xhold1594 hold47/X vssd1 vssd1 vccd1 vccd1 hold1594/X sky130_fd_sc_hd__buf_2
Xhold1583 hold1583/A vssd1 vssd1 vccd1 vccd1 _5090_/D sky130_fd_sc_hd__buf_2
XFILLER_45_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1572 hold2429/X vssd1 vssd1 vccd1 vccd1 hold2430/A sky130_fd_sc_hd__buf_2
XFILLER_45_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3060_ _3099_/B _3058_/X _3059_/X vssd1 vssd1 vccd1 vccd1 _3060_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4920__505 _4921__506/A vssd1 vssd1 vccd1 vccd1 _5641_/CLK sky130_fd_sc_hd__inv_2
X_3962_ _4390_/A _3962_/B vssd1 vssd1 vccd1 vccd1 _3962_/Y sky130_fd_sc_hd__nor2_4
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701_ _5701_/CLK _5701_/D vssd1 vssd1 vccd1 vccd1 _5701_/Q sky130_fd_sc_hd__dfxtp_1
X_2913_ _3004_/C1 _2910_/X _2912_/X vssd1 vssd1 vccd1 vccd1 _2913_/X sky130_fd_sc_hd__a21o_2
X_3893_ _5748_/Q _3888_/Y _3892_/X _3887_/X vssd1 vssd1 vccd1 vccd1 _3893_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2844_ _5400_/Q _3536_/A0 _2851_/S vssd1 vssd1 vccd1 vccd1 _5400_/D sky130_fd_sc_hd__mux2_1
X_5632_ _5632_/CLK _5632_/D vssd1 vssd1 vccd1 vccd1 _5632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5563_ _5564_/CLK _5563_/D vssd1 vssd1 vccd1 vccd1 _5563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2775_ _3396_/A0 _5457_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5457_/D sky130_fd_sc_hd__mux2_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__buf_2
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold113 hold126/X vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__buf_2
X_5494_ _5494_/CLK _5494_/D vssd1 vssd1 vccd1 vccd1 _5494_/Q sky130_fd_sc_hd__dfxtp_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__buf_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold146 hold160/X vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__buf_2
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__buf_2
Xhold157 hold173/X vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__buf_2
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout604 _3538_/A0 vssd1 vssd1 vccd1 vccd1 _3601_/A1 sky130_fd_sc_hd__buf_4
Xfanout615 _5320_/Q vssd1 vssd1 vccd1 vccd1 _3613_/A1 sky130_fd_sc_hd__buf_2
XFILLER_113_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4376_ _5737_/Q _4370_/X _4376_/B1 hold875/X vssd1 vssd1 vccd1 vccd1 _4376_/X sky130_fd_sc_hd__o211a_1
Xhold179 hold297/X vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__buf_2
Xfanout648 _4360_/A vssd1 vssd1 vccd1 vccd1 hold367/A sky130_fd_sc_hd__clkbuf_8
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout626 _5291_/Q vssd1 vssd1 vccd1 vccd1 _3914_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout637 _2466_/Y vssd1 vssd1 vccd1 vccd1 _3824_/A1 sky130_fd_sc_hd__buf_12
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _5655_/Q _5385_/Q _3327_/S vssd1 vssd1 vccd1 vccd1 _3328_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3325_/A _3256_/X _3257_/X vssd1 vssd1 vccd1 vccd1 _3258_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3189_ _5644_/Q _5636_/Q _5047_/Q _5652_/Q _3284_/S _3201_/S1 vssd1 vssd1 vccd1 vccd1
+ _3189_/X sky130_fd_sc_hd__mux4_2
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663__248 _4478__63/A vssd1 vssd1 vccd1 vccd1 _5351_/CLK sky130_fd_sc_hd__inv_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4704__289 _4744__329/A vssd1 vssd1 vccd1 vccd1 _5395_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4557__142 _4421__6/A vssd1 vssd1 vccd1 vccd1 _5199_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold691 _4400_/X vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__buf_2
XFILLER_134_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2070 hold2070/A vssd1 vssd1 vccd1 vccd1 _5346_/D sky130_fd_sc_hd__buf_2
Xhold2081 _3786_/X vssd1 vssd1 vccd1 vccd1 hold2081/X sky130_fd_sc_hd__buf_2
XFILLER_94_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1380 hold2136/X vssd1 vssd1 vccd1 vccd1 hold2137/A sky130_fd_sc_hd__buf_2
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput207 _3661_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2560_ _2743_/A0 _5652_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5652_/D sky130_fd_sc_hd__mux2_1
Xoutput229 _3665_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput218 _3662_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2491_ _3844_/A _5111_/Q vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__nand2_4
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4230_ _5559_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__or2_1
X_4161_ _4152_/Y _4153_/X _4170_/B _4157_/X _4160_/Y vssd1 vssd1 vccd1 vccd1 _4162_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3112_ _5373_/Q _3443_/B _3453_/C vssd1 vssd1 vccd1 vccd1 _3544_/B sky130_fd_sc_hd__or3_4
X_4092_ _3928_/A _4361_/B _3897_/C _4357_/C _4401_/A vssd1 vssd1 vccd1 vccd1 _4092_/X
+ sky130_fd_sc_hd__o2111a_1
X_3043_ _3043_/A _3043_/B _3043_/C vssd1 vssd1 vccd1 vccd1 _3043_/X sky130_fd_sc_hd__or3_1
XFILLER_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _5246_/CLK _4994_/D vssd1 vssd1 vccd1 vccd1 _4994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3945_ _5249_/Q _5102_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _5102_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ _5751_/Q _3998_/A1 _3882_/A3 _3887_/A vssd1 vssd1 vccd1 vccd1 _3876_/X sky130_fd_sc_hd__a31o_1
X_5615_ _5615_/CLK _5615_/D vssd1 vssd1 vccd1 vccd1 _5615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2827_ _3390_/A0 _5415_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5415_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5546_ _5546_/CLK _5546_/D vssd1 vssd1 vccd1 vccd1 _5546_/Q sky130_fd_sc_hd__dfxtp_1
X_2758_ _3370_/A _3388_/B vssd1 vssd1 vccd1 vccd1 _2766_/S sky130_fd_sc_hd__or2_4
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5477_ _5477_/CLK _5477_/D vssd1 vssd1 vccd1 vccd1 _5477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2689_ _3603_/A1 _5534_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5534_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout423 _3953_/S vssd1 vssd1 vccd1 vccd1 _4000_/S sky130_fd_sc_hd__buf_6
Xfanout412 _3353_/A vssd1 vssd1 vccd1 vccd1 _3357_/A sky130_fd_sc_hd__clkbuf_4
Xfanout434 _3621_/X vssd1 vssd1 vccd1 vccd1 _3660_/B sky130_fd_sc_hd__buf_4
Xfanout456 _2874_/Y vssd1 vssd1 vccd1 vccd1 _3043_/A sky130_fd_sc_hd__buf_6
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4359_ _5374_/Q _4365_/A vssd1 vssd1 vccd1 vccd1 _5725_/D sky130_fd_sc_hd__and2_1
Xfanout445 _4381_/X vssd1 vssd1 vccd1 vccd1 _4389_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout478 _3004_/C1 vssd1 vssd1 vccd1 vccd1 _3073_/C1 sky130_fd_sc_hd__buf_6
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout489 _3795_/B1 vssd1 vssd1 vccd1 vccd1 _3796_/B1 sky130_fd_sc_hd__buf_8
Xfanout467 _3131_/Y vssd1 vssd1 vccd1 vccd1 _3316_/C1 sky130_fd_sc_hd__buf_6
XFILLER_86_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5754_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4791__376 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5482_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4685__270 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _3733_/A1 _3728_/X _3729_/X split2/A vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__o211a_1
XFILLER_146_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _3661_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3661_/X sky130_fd_sc_hd__and2_1
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5400_ _5400_/CLK _5400_/D vssd1 vssd1 vccd1 vccd1 _5400_/Q sky130_fd_sc_hd__dfxtp_1
X_3592_ _5031_/Q _3592_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5031_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_75_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5565_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2612_ _3569_/A1 _5608_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5608_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2543_ _3579_/A0 _5700_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5700_/D sky130_fd_sc_hd__mux2_1
X_5331_ _5331_/CLK _5331_/D vssd1 vssd1 vccd1 vccd1 _5331_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5262_ _5262_/CLK _5262_/D vssd1 vssd1 vccd1 vccd1 _5262_/Q sky130_fd_sc_hd__dfxtp_1
X_2474_ _3350_/A _3312_/S vssd1 vssd1 vccd1 vccd1 _3122_/A sky130_fd_sc_hd__or2_1
X_5193_ _5193_/CLK _5193_/D vssd1 vssd1 vccd1 vccd1 _5193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4213_ _4217_/A _4213_/B vssd1 vssd1 vccd1 vccd1 _5552_/D sky130_fd_sc_hd__nor2_1
Xhold2806 hold2806/A vssd1 vssd1 vccd1 vccd1 hold2806/X sky130_fd_sc_hd__buf_2
X_4144_ _4142_/X _4143_/Y _4137_/Y _4138_/Y _4139_/X vssd1 vssd1 vccd1 vccd1 _4145_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4926__511 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5647_/CLK sky130_fd_sc_hd__inv_2
X_4075_ _4075_/A _4075_/B _4074_/C _4074_/D vssd1 vssd1 vccd1 vccd1 _4078_/A sky130_fd_sc_hd__or4bb_4
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3026_ _3034_/A _3024_/X _3025_/X vssd1 vssd1 vccd1 vccd1 _3026_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4977_ _4977_/CLK _4977_/D vssd1 vssd1 vccd1 vccd1 _4977_/Q sky130_fd_sc_hd__dfxtp_1
X_3928_ _3928_/A _4281_/A _4361_/B _4091_/B vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__or4b_2
XFILLER_126_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3859_ _4399_/B _3847_/X _3858_/X _4361_/A vssd1 vssd1 vccd1 vccd1 _3859_/X sky130_fd_sc_hd__a31o_1
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5529_ _5557_/CLK _5529_/D vssd1 vssd1 vccd1 vccd1 _5529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4669__254 _5004_/CLK vssd1 vssd1 vccd1 vccd1 _5357_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_122_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5016_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5880_ _5880_/A vssd1 vssd1 vccd1 vccd1 _5880_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3713_ _5074_/Q input33/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3713_/X sky130_fd_sc_hd__mux2_4
XFILLER_147_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3644_ _3644_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__or2_1
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3575_ _3575_/A0 _5046_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5046_/D sky130_fd_sc_hd__mux2_1
X_5314_ _5314_/CLK _5314_/D vssd1 vssd1 vccd1 vccd1 _5314_/Q sky130_fd_sc_hd__dfxtp_1
X_2526_ _3389_/A0 _5715_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5715_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2457_ _5530_/Q vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__inv_2
X_5245_ _5246_/CLK _5245_/D vssd1 vssd1 vccd1 vccd1 _5245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__buf_2
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2625 _4390_/X vssd1 vssd1 vccd1 vccd1 hold2625/X sky130_fd_sc_hd__buf_2
Xhold2636 hold2636/A vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__buf_2
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__buf_2
XFILLER_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5176_ _5176_/CLK _5176_/D vssd1 vssd1 vccd1 vccd1 _5176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2658 hold682/X vssd1 vssd1 vccd1 vccd1 hold2658/X sky130_fd_sc_hd__buf_2
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__buf_2
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4127_ _4128_/B _4128_/C vssd1 vssd1 vccd1 vccd1 _4127_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4058_ _4259_/B _4259_/C vssd1 vssd1 vccd1 vccd1 _4058_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3009_ _5172_/Q _5236_/Q _3040_/S vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput390 _3762_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4797__382 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5488_/CLK sky130_fd_sc_hd__inv_2
XFILLER_143_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3360_ _3281_/S _3353_/A _3359_/Y vssd1 vssd1 vccd1 vccd1 _5326_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/CLK _5030_/D vssd1 vssd1 vccd1 vccd1 _5030_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _5701_/Q _3331_/A2 _3326_/B2 _5717_/Q vssd1 vssd1 vccd1 vccd1 _3291_/X sky130_fd_sc_hd__o22a_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5932_ _5932_/A vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5863_ _5863_/A vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_90_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4875__460/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3627_ _3627_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3627_/X sky130_fd_sc_hd__and2_1
XFILLER_119_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3558_ _5061_/Q _3603_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5061_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2509_ _5097_/Q _5098_/Q _3930_/C _5089_/Q vssd1 vssd1 vccd1 vccd1 _2510_/C sky130_fd_sc_hd__or4b_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput118 probe_out[84] vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__clkbuf_2
Xinput107 probe_out[74] vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4590__175 _4438__23/A vssd1 vssd1 vccd1 vccd1 _5240_/CLK sky130_fd_sc_hd__inv_2
X_3489_ _3597_/A1 _5170_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5170_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2422 hold2422/A vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__buf_2
Xhold2411 hold2411/A vssd1 vssd1 vccd1 vccd1 hold2411/X sky130_fd_sc_hd__buf_2
Xinput129 probe_out[94] vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__clkbuf_2
X_5228_ _5228_/CLK _5228_/D vssd1 vssd1 vccd1 vccd1 _5228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1710 hold2228/X vssd1 vssd1 vccd1 vccd1 hold2229/A sky130_fd_sc_hd__buf_2
Xhold2455 hold2455/A vssd1 vssd1 vccd1 vccd1 input139/A sky130_fd_sc_hd__buf_2
Xhold2433 hold39/X vssd1 vssd1 vccd1 vccd1 hold2433/X sky130_fd_sc_hd__buf_2
Xhold2444 hold2444/A vssd1 vssd1 vccd1 vccd1 hold2444/X sky130_fd_sc_hd__buf_2
X_5159_ _5159_/CLK _5159_/D vssd1 vssd1 vccd1 vccd1 _5159_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2488 hold793/X vssd1 vssd1 vccd1 vccd1 hold2488/X sky130_fd_sc_hd__buf_2
Xhold2477 hold2477/A vssd1 vssd1 vccd1 vccd1 hold2477/X sky130_fd_sc_hd__buf_2
XFILLER_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1721 hold2384/X vssd1 vssd1 vccd1 vccd1 hold2385/A sky130_fd_sc_hd__buf_2
Xhold2499 hold2499/A vssd1 vssd1 vccd1 vccd1 hold2499/X sky130_fd_sc_hd__buf_2
Xhold1765 hold2477/X vssd1 vssd1 vccd1 vccd1 hold2478/A sky130_fd_sc_hd__buf_2
XFILLER_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1754 hold2564/X vssd1 vssd1 vccd1 vccd1 hold2565/A sky130_fd_sc_hd__buf_2
Xhold1798 hold2510/X vssd1 vssd1 vccd1 vccd1 hold2511/A sky130_fd_sc_hd__buf_2
XFILLER_72_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_80 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4831__416 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4725__310 _5247_/CLK vssd1 vssd1 vccd1 vccd1 _5416_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2860_ _5385_/Q _3396_/A0 _2860_/S vssd1 vssd1 vccd1 vccd1 _5385_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2791_ _3409_/A1 _5446_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5446_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XCaravelHost_713 vssd1 vssd1 vccd1 vccd1 CaravelHost_713/HI partID[5] sky130_fd_sc_hd__conb_1
XCaravelHost_702 vssd1 vssd1 vccd1 vccd1 CaravelHost_702/HI manufacturerID[2] sky130_fd_sc_hd__conb_1
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XCaravelHost_724 vssd1 vssd1 vccd1 vccd1 partID[2] CaravelHost_724/LO sky130_fd_sc_hd__conb_1
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__buf_2
XFILLER_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold328 hold328/A vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__buf_2
X_3412_ _5268_/Q _3568_/A1 _3414_/S vssd1 vssd1 vccd1 vccd1 _5268_/D sky130_fd_sc_hd__mux2_1
X_4574__159 _4438__23/A vssd1 vssd1 vccd1 vccd1 _5224_/CLK sky130_fd_sc_hd__inv_2
X_4392_ _5744_/Q _4398_/A2 _4392_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4392_/X sky130_fd_sc_hd__o211a_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _2545_/A _3350_/B _3562_/B _3342_/X _4093_/B vssd1 vssd1 vccd1 vccd1 _5335_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1006 hold1566/X vssd1 vssd1 vccd1 vccd1 hold1567/A sky130_fd_sc_hd__buf_2
XFILLER_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3336_/A1 _3255_/X _3258_/X _3273_/X _3136_/X vssd1 vssd1 vccd1 vccd1 _3274_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_112_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5013_ _5262_/CLK _5013_/D vssd1 vssd1 vccd1 vccd1 _5013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1039 hold1648/X vssd1 vssd1 vccd1 vccd1 hold1649/A sky130_fd_sc_hd__buf_2
Xhold1028 hold2453/X vssd1 vssd1 vccd1 vccd1 hold2454/A sky130_fd_sc_hd__buf_2
Xhold1017 hold1600/X vssd1 vssd1 vccd1 vccd1 hold1601/A sky130_fd_sc_hd__buf_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5915_ _5915_/A vssd1 vssd1 vccd1 vccd1 _5915_/X sky130_fd_sc_hd__clkbuf_4
X_5846_ _5846_/A vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ _3041_/B1 _2987_/X _2988_/X vssd1 vssd1 vccd1 vccd1 _3012_/B sky130_fd_sc_hd__o21a_1
XFILLER_10_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold862 hold862/A vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__buf_2
Xhold873 hold873/A vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__buf_2
XFILLER_143_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2230 hold641/X vssd1 vssd1 vccd1 vccd1 hold2230/X sky130_fd_sc_hd__buf_2
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2263 hold2263/A vssd1 vssd1 vccd1 vccd1 input163/A sky130_fd_sc_hd__buf_2
Xhold2252 hold2252/A vssd1 vssd1 vccd1 vccd1 input162/A sky130_fd_sc_hd__buf_2
Xhold2241 hold2241/A vssd1 vssd1 vccd1 vccd1 input161/A sky130_fd_sc_hd__buf_2
Xhold2285 hold2285/A vssd1 vssd1 vccd1 vccd1 hold2285/X sky130_fd_sc_hd__buf_2
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2274 _3668_/A vssd1 vssd1 vccd1 vccd1 hold2274/X sky130_fd_sc_hd__buf_2
Xhold1551 hold2425/X vssd1 vssd1 vccd1 vccd1 hold2426/A sky130_fd_sc_hd__buf_2
Xhold1562 hold2413/X vssd1 vssd1 vccd1 vccd1 hold2414/A sky130_fd_sc_hd__buf_2
Xhold1540 hold2394/X vssd1 vssd1 vccd1 vccd1 hold2395/A sky130_fd_sc_hd__buf_2
Xhold2296 _3669_/A vssd1 vssd1 vccd1 vccd1 hold2296/X sky130_fd_sc_hd__buf_2
X_4475__60 _4507__92/A vssd1 vssd1 vccd1 vccd1 _5117_/CLK sky130_fd_sc_hd__inv_2
Xhold1595 hold1595/A vssd1 vssd1 vccd1 vccd1 _5099_/D sky130_fd_sc_hd__buf_2
XFILLER_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1584 hold2439/X vssd1 vssd1 vccd1 vccd1 hold2440/A sky130_fd_sc_hd__buf_2
Xhold1573 hold2431/X vssd1 vssd1 vccd1 vccd1 hold2432/A sky130_fd_sc_hd__buf_2
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4421__6/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _3829_/A _3829_/B _4403_/B1 vssd1 vssd1 vccd1 vccd1 _3961_/Y sky130_fd_sc_hd__a21oi_1
X_2912_ _3029_/B1 _2911_/X _2919_/B vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5700_ _5700_/CLK _5700_/D vssd1 vssd1 vccd1 vccd1 _5700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3892_ _4401_/A _5209_/Q _3897_/C _3855_/X vssd1 vssd1 vccd1 vccd1 _3892_/X sky130_fd_sc_hd__a31o_1
X_2843_ _3607_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2851_/S sky130_fd_sc_hd__nor2_8
X_5631_ _5631_/CLK _5631_/D vssd1 vssd1 vccd1 vccd1 _5631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5562_ _5564_/CLK _5562_/D vssd1 vssd1 vccd1 vccd1 _5562_/Q sky130_fd_sc_hd__dfxtp_1
X_2774_ _3395_/A0 _5458_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5458_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold103 hold139/X vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__buf_2
X_5493_ _5493_/CLK _5493_/D vssd1 vssd1 vccd1 vccd1 _5493_/Q sky130_fd_sc_hd__dfxtp_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__buf_2
Xhold114 hold128/X vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__buf_2
Xhold158 hold175/X vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__buf_2
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__buf_2
Xhold147 _3978_/X vssd1 vssd1 vccd1 vccd1 _5248_/D sky130_fd_sc_hd__buf_2
Xfanout605 _5323_/Q vssd1 vssd1 vccd1 vccd1 _3538_/A0 sky130_fd_sc_hd__buf_2
X_4375_ _3647_/A _3778_/B _4370_/X vssd1 vssd1 vccd1 vccd1 _4375_/X sky130_fd_sc_hd__a21bo_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__buf_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout616 _5320_/Q vssd1 vssd1 vccd1 vccd1 _3604_/A1 sky130_fd_sc_hd__buf_4
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout649 _4360_/A vssd1 vssd1 vccd1 vccd1 hold379/A sky130_fd_sc_hd__clkbuf_4
Xfanout627 _4401_/A vssd1 vssd1 vccd1 vccd1 _3998_/A1 sky130_fd_sc_hd__buf_4
XFILLER_59_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3326_ _2482_/B _5301_/Q _5050_/Q _3326_/B2 _3326_/C1 vssd1 vssd1 vccd1 vccd1 _3326_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout638 _4351_/A vssd1 vssd1 vccd1 vccd1 _3711_/B sky130_fd_sc_hd__buf_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _5617_/Q _2464_/A _3128_/B _5609_/Q _3316_/C1 vssd1 vssd1 vccd1 vccd1 _3257_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3188_ _5612_/Q _5596_/Q _5580_/Q _5620_/Q _3318_/S _3130_/B vssd1 vssd1 vccd1 vccd1
+ _3188_/X sky130_fd_sc_hd__mux4_2
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4596__181 _4460__45/A vssd1 vssd1 vccd1 vccd1 _5270_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold692 _4402_/X vssd1 vssd1 vccd1 vccd1 _5748_/D sky130_fd_sc_hd__buf_2
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2082 hold2082/A vssd1 vssd1 vccd1 vccd1 hold445/A sky130_fd_sc_hd__buf_2
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4943__528 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5701_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1381 hold2138/X vssd1 vssd1 vccd1 vccd1 hold2139/A sky130_fd_sc_hd__buf_2
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4837__422 _4463__48/A vssd1 vssd1 vccd1 vccd1 _5528_/CLK sky130_fd_sc_hd__inv_2
Xoutput208 _3671_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__clkbuf_2
Xoutput219 _3681_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2490_ _3844_/A _3955_/A vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__and2_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4253_/A _4160_/B vssd1 vssd1 vccd1 vccd1 _4160_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3111_ _5355_/Q _3543_/A0 _3111_/S vssd1 vssd1 vccd1 vccd1 _5355_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ _4091_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4357_/C sky130_fd_sc_hd__and2_4
X_3042_ _3039_/X _3041_/X _2919_/B _3038_/X vssd1 vssd1 vccd1 vccd1 _3042_/X sky130_fd_sc_hd__a211o_1
XFILLER_95_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _5244_/CLK _4993_/D vssd1 vssd1 vccd1 vccd1 _4993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3944_ _3944_/A0 _5101_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3944_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3875_ _5069_/Q _3959_/A _3875_/B1 vssd1 vssd1 vccd1 vccd1 _3875_/X sky130_fd_sc_hd__a21o_1
X_5614_ _5614_/CLK _5614_/D vssd1 vssd1 vccd1 vccd1 _5614_/Q sky130_fd_sc_hd__dfxtp_1
X_2826_ _3389_/A0 _5416_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5416_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5545_ _5546_/CLK _5545_/D vssd1 vssd1 vccd1 vccd1 _5545_/Q sky130_fd_sc_hd__dfxtp_2
X_2757_ _3396_/A0 _5473_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5473_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2688_ _3602_/A1 _5535_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5535_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ _5476_/CLK _5476_/D vssd1 vssd1 vccd1 vccd1 _5476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout413 _3125_/Y vssd1 vssd1 vccd1 vccd1 _3353_/A sky130_fd_sc_hd__buf_4
Xfanout457 _2874_/Y vssd1 vssd1 vccd1 vccd1 _3045_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout435 _2863_/Y vssd1 vssd1 vccd1 vccd1 _3094_/A sky130_fd_sc_hd__buf_4
X_4358_ _4358_/A _4358_/B vssd1 vssd1 vccd1 vccd1 _4358_/Y sky130_fd_sc_hd__nor2_2
Xfanout424 hold317/X vssd1 vssd1 vccd1 vccd1 hold318/A sky130_fd_sc_hd__clkbuf_16
Xfanout446 _3619_/Y vssd1 vssd1 vccd1 vccd1 _3931_/B sky130_fd_sc_hd__buf_8
X_4630__215 _4463__48/A vssd1 vssd1 vccd1 vccd1 _5307_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout479 _2869_/Y vssd1 vssd1 vccd1 vccd1 _3004_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4289_ _4283_/C _4322_/B _4288_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5664_/D sky130_fd_sc_hd__o211a_1
X_3309_ _5513_/Q _5282_/Q _3330_/S vssd1 vssd1 vccd1 vccd1 _3309_/X sky130_fd_sc_hd__mux2_2
Xfanout468 _3131_/Y vssd1 vssd1 vccd1 vccd1 _3326_/C1 sky130_fd_sc_hd__buf_4
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4445__30 _4468__53/A vssd1 vssd1 vccd1 vccd1 _5039_/CLK sky130_fd_sc_hd__inv_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3660_ _3660_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3660_/X sky130_fd_sc_hd__or2_1
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3591_ _5032_/Q _3591_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5032_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2611_ _3577_/A0 _5609_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5609_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2542_ _3569_/A1 _5701_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5701_/D sky130_fd_sc_hd__mux2_1
X_5330_ _5330_/CLK _5330_/D vssd1 vssd1 vccd1 vccd1 _5330_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5261_ _5261_/CLK _5261_/D vssd1 vssd1 vccd1 vccd1 _5261_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4962__547/A sky130_fd_sc_hd__clkbuf_8
XFILLER_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4212_ _5552_/Q _4209_/B _4210_/C _4155_/B vssd1 vssd1 vccd1 vccd1 _4213_/B sky130_fd_sc_hd__o2bb2a_1
X_2473_ _5332_/Q _3127_/A vssd1 vssd1 vccd1 vccd1 _3123_/A sky130_fd_sc_hd__xor2_1
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5192_ _5192_/CLK _5192_/D vssd1 vssd1 vccd1 vccd1 _5192_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_44_wb_clk_i _4676__261/A vssd1 vssd1 vccd1 vccd1 _5383_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2807 hold2807/A vssd1 vssd1 vccd1 vccd1 hold2807/X sky130_fd_sc_hd__buf_2
XFILLER_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4143_ _4142_/B _4142_/C _5753_/Q vssd1 vssd1 vccd1 vccd1 _4143_/Y sky130_fd_sc_hd__a21oi_1
X_4074_ _4075_/A _4075_/B _4074_/C _4074_/D vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__and4bb_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4965__550 _4965__550/A vssd1 vssd1 vccd1 vccd1 _5723_/CLK sky130_fd_sc_hd__inv_2
X_3025_ _5600_/Q _5366_/Q _3073_/B2 _5584_/Q _3073_/C1 vssd1 vssd1 vccd1 vccd1 _3025_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4976_ _4976_/CLK _4976_/D vssd1 vssd1 vccd1 vccd1 _4976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3927_ _4399_/B _3927_/B vssd1 vssd1 vccd1 vccd1 _4091_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3858_ _3887_/B _3856_/X _3857_/Y _5729_/Q _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3858_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2809_ _3501_/A1 _5431_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5431_/D sky130_fd_sc_hd__mux2_1
X_3789_ _3789_/A1 _5021_/Q _3829_/A _3796_/B1 _4989_/Q vssd1 vssd1 vccd1 vccd1 _3789_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_119_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5528_ _5528_/CLK _5528_/D vssd1 vssd1 vccd1 vccd1 _5528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5459_ _5459_/CLK _5459_/D vssd1 vssd1 vccd1 vccd1 _5459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4949__534 _4965__550/A vssd1 vssd1 vccd1 vccd1 _5707_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3712_ _3718_/A1 _3710_/X _3711_/X split2/X vssd1 vssd1 vccd1 vccd1 _3712_/X sky130_fd_sc_hd__o211a_1
X_3643_ _3643_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3643_/X sky130_fd_sc_hd__or2_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5313_ _5313_/CLK _5313_/D vssd1 vssd1 vccd1 vccd1 _5313_/Q sky130_fd_sc_hd__dfxtp_1
X_3574_ _3574_/A0 _5047_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5047_/D sky130_fd_sc_hd__mux2_1
X_2525_ _3562_/A _2788_/A vssd1 vssd1 vccd1 vccd1 _2533_/S sky130_fd_sc_hd__or2_4
XFILLER_142_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2456_ _5548_/Q vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__inv_2
Xhold2604 _4357_/X vssd1 vssd1 vccd1 vccd1 hold2604/X sky130_fd_sc_hd__buf_2
X_5244_ _5244_/CLK _5244_/D vssd1 vssd1 vccd1 vccd1 _5244_/Q sky130_fd_sc_hd__dfxtp_1
X_5175_ _5175_/CLK _5175_/D vssd1 vssd1 vccd1 vccd1 _5175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2626 hold2626/A vssd1 vssd1 vccd1 vccd1 hold2626/X sky130_fd_sc_hd__buf_2
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__buf_2
Xhold2637 hold240/X vssd1 vssd1 vccd1 vccd1 hold2637/X sky130_fd_sc_hd__buf_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__buf_2
XFILLER_84_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2659 hold2659/A vssd1 vssd1 vccd1 vccd1 hold2659/X sky130_fd_sc_hd__buf_2
X_4126_ _5544_/Q _5543_/Q _4132_/B _5545_/Q vssd1 vssd1 vccd1 vccd1 _4128_/C sky130_fd_sc_hd__a31o_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _5666_/Q _5665_/Q _5667_/Q vssd1 vssd1 vccd1 vccd1 _4259_/C sky130_fd_sc_hd__a21o_1
X_3008_ _5220_/Q _2873_/B _2870_/B vssd1 vssd1 vccd1 vccd1 _3008_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4742__327 _5005_/CLK vssd1 vssd1 vccd1 vccd1 _5433_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4636__221 _4514__99/A vssd1 vssd1 vccd1 vccd1 _5314_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput380 _3739_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput391 _3764_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _5267_/Q _5294_/Q _3290_/S vssd1 vssd1 vccd1 vccd1 _3290_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _5931_/A vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5862_ _5862_/A vssd1 vssd1 vccd1 vccd1 _5862_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3626_ _3626_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3626_/X sky130_fd_sc_hd__and2_1
XFILLER_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3557_ _5062_/Q _3611_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5062_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2508_ _3930_/C _2512_/B _2512_/C _2512_/D vssd1 vssd1 vccd1 vccd1 _3850_/B sky130_fd_sc_hd__or4_2
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput108 probe_out[75] vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__clkbuf_2
X_5227_ _5227_/CLK _5227_/D vssd1 vssd1 vccd1 vccd1 _5227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3488_ _3596_/A1 _5171_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5171_/D sky130_fd_sc_hd__mux2_1
Xhold2401 _4408_/X vssd1 vssd1 vccd1 vccd1 hold2401/X sky130_fd_sc_hd__buf_2
Xhold2412 hold2412/A vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__buf_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput119 probe_out[85] vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__clkbuf_2
Xhold1711 hold2230/X vssd1 vssd1 vccd1 vccd1 hold2231/A sky130_fd_sc_hd__buf_2
X_2439_ _5679_/Q vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__inv_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2423 hold15/X vssd1 vssd1 vccd1 vccd1 hold2423/X sky130_fd_sc_hd__buf_2
Xhold2445 hold2445/A vssd1 vssd1 vccd1 vccd1 hold2445/X sky130_fd_sc_hd__buf_2
Xhold2434 hold2434/A vssd1 vssd1 vccd1 vccd1 hold2434/X sky130_fd_sc_hd__buf_2
XFILLER_130_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _5158_/CLK _5158_/D vssd1 vssd1 vccd1 vccd1 _5158_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2489 hold2489/A vssd1 vssd1 vccd1 vccd1 hold2489/X sky130_fd_sc_hd__buf_2
Xhold2478 hold2478/A vssd1 vssd1 vccd1 vccd1 _5318_/D sky130_fd_sc_hd__buf_2
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1744 hold2549/X vssd1 vssd1 vccd1 vccd1 hold2550/A sky130_fd_sc_hd__buf_2
Xhold2456 _3674_/A vssd1 vssd1 vccd1 vccd1 hold2456/X sky130_fd_sc_hd__buf_2
XFILLER_29_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5089_ _5730_/CLK _5089_/D vssd1 vssd1 vccd1 vccd1 _5089_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1755 hold2566/X vssd1 vssd1 vccd1 vccd1 hold2567/A sky130_fd_sc_hd__buf_2
X_4109_ _4132_/B _4119_/C _4104_/D _4114_/B _2455_/Y vssd1 vssd1 vccd1 vccd1 _4110_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1799 hold2512/X vssd1 vssd1 vccd1 vccd1 hold2513/A sky130_fd_sc_hd__buf_2
XFILLER_72_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_81 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_70 hold90/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4870__455 _4875__460/A vssd1 vssd1 vccd1 vccd1 _5591_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4911__496 _4449__34/A vssd1 vssd1 vccd1 vccd1 _5632_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4805__390 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5496_/CLK sky130_fd_sc_hd__inv_2
X_2790_ _2790_/A0 _5447_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5447_/D sky130_fd_sc_hd__mux2_1
XCaravelHost_703 vssd1 vssd1 vccd1 vccd1 CaravelHost_703/HI manufacturerID[3] sky130_fd_sc_hd__conb_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_714 vssd1 vssd1 vccd1 vccd1 CaravelHost_714/HI partID[7] sky130_fd_sc_hd__conb_1
XCaravelHost_725 vssd1 vssd1 vccd1 vccd1 partID[4] CaravelHost_725/LO sky130_fd_sc_hd__conb_1
XFILLER_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold318 hold318/A vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__buf_2
X_4391_ _3640_/A _4389_/B _4398_/A2 vssd1 vssd1 vccd1 vccd1 _4391_/X sky130_fd_sc_hd__a21bo_1
X_3411_ _5269_/Q _3576_/A0 _3414_/S vssd1 vssd1 vccd1 vccd1 _5269_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3342_ _5334_/Q _5333_/Q _3349_/A _5335_/Q vssd1 vssd1 vccd1 vccd1 _3342_/X sky130_fd_sc_hd__a31o_1
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3273_ _3263_/X _3264_/X _3353_/B _3261_/X vssd1 vssd1 vccd1 vccd1 _3273_/X sky130_fd_sc_hd__a211o_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5012_ _5265_/CLK _5012_/D vssd1 vssd1 vccd1 vccd1 _5012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1007 hold1568/X vssd1 vssd1 vccd1 vccd1 hold1569/A sky130_fd_sc_hd__buf_2
Xhold1018 hold1602/X vssd1 vssd1 vccd1 vccd1 hold1603/A sky130_fd_sc_hd__buf_2
Xhold1029 hold1612/X vssd1 vssd1 vccd1 vccd1 hold1613/A sky130_fd_sc_hd__buf_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5914_ _5914_/A vssd1 vssd1 vccd1 vccd1 _5914_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5845_ _5845_/A vssd1 vssd1 vccd1 vccd1 _5845_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2988_ _2867_/A _5132_/Q _3041_/A2 _5140_/Q _3064_/C1 vssd1 vssd1 vccd1 vccd1 _2988_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4854__439 _4875__460/A vssd1 vssd1 vccd1 vccd1 _5575_/CLK sky130_fd_sc_hd__inv_2
X_3609_ _4973_/Q _3609_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4973_/D sky130_fd_sc_hd__mux2_1
Xinput90 probe_out[59] vssd1 vssd1 vccd1 vccd1 _5896_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold863 hold863/A vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__buf_2
Xhold852 hold852/A vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__buf_2
Xhold841 hold841/A vssd1 vssd1 vccd1 vccd1 hold841/X sky130_fd_sc_hd__buf_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold874 hold874/A vssd1 vssd1 vccd1 vccd1 hold874/X sky130_fd_sc_hd__buf_2
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2220 hold2220/A vssd1 vssd1 vccd1 vccd1 hold2220/X sky130_fd_sc_hd__buf_2
XFILLER_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2231 hold2231/A vssd1 vssd1 vccd1 vccd1 hold2231/X sky130_fd_sc_hd__buf_2
XFILLER_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2242 _3665_/A vssd1 vssd1 vccd1 vccd1 hold2242/X sky130_fd_sc_hd__buf_2
Xhold2264 _3667_/A vssd1 vssd1 vccd1 vccd1 hold2264/X sky130_fd_sc_hd__buf_2
Xhold2253 _3666_/A vssd1 vssd1 vccd1 vccd1 hold2253/X sky130_fd_sc_hd__buf_2
X_4748__333 _5261_/CLK vssd1 vssd1 vccd1 vccd1 _5439_/CLK sky130_fd_sc_hd__inv_2
Xhold2286 hold2286/A vssd1 vssd1 vccd1 vccd1 hold2286/X sky130_fd_sc_hd__buf_2
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2297 hold2297/A vssd1 vssd1 vccd1 vccd1 hold981/A sky130_fd_sc_hd__buf_2
Xhold2275 hold2275/A vssd1 vssd1 vccd1 vccd1 hold975/A sky130_fd_sc_hd__buf_2
Xhold1552 hold2427/X vssd1 vssd1 vccd1 vccd1 hold2428/A sky130_fd_sc_hd__buf_2
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1530 hold37/X vssd1 vssd1 vccd1 vccd1 hold994/A sky130_fd_sc_hd__buf_2
Xhold1541 hold987/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__buf_2
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1574 hold2433/X vssd1 vssd1 vccd1 vccd1 hold2434/A sky130_fd_sc_hd__buf_2
Xhold1585 hold2441/X vssd1 vssd1 vccd1 vccd1 hold2442/A sky130_fd_sc_hd__buf_2
Xhold1563 hold2415/X vssd1 vssd1 vccd1 vccd1 hold2416/A sky130_fd_sc_hd__buf_2
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1596 hold2457/X vssd1 vssd1 vccd1 vccd1 hold2458/A sky130_fd_sc_hd__buf_2
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4490__75 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5132_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3960_ _3960_/A _3960_/B _3960_/C vssd1 vssd1 vccd1 vccd1 _3960_/X sky130_fd_sc_hd__and3_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2911_ _5431_/Q _5407_/Q _5399_/Q _5439_/Q _3069_/S _2942_/S1 vssd1 vssd1 vccd1 vccd1
+ _2911_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_69_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4514__99/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _4399_/B _3889_/X hold536/X vssd1 vssd1 vccd1 vccd1 _3891_/X sky130_fd_sc_hd__a21o_1
X_4541__126 _4421__6/A vssd1 vssd1 vccd1 vccd1 _5183_/CLK sky130_fd_sc_hd__inv_2
X_2842_ _3543_/A0 _5401_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5401_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5630_ _5630_/CLK _5630_/D vssd1 vssd1 vccd1 vccd1 _5630_/Q sky130_fd_sc_hd__dfxtp_1
X_5561_ _5564_/CLK _5561_/D vssd1 vssd1 vccd1 vccd1 _5561_/Q sky130_fd_sc_hd__dfxtp_1
X_2773_ _3394_/A0 _5459_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5459_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5492_ _5492_/CLK _5492_/D vssd1 vssd1 vccd1 vccd1 _5492_/Q sky130_fd_sc_hd__dfxtp_1
Xhold104 hold141/X vssd1 vssd1 vccd1 vccd1 _3989_/B sky130_fd_sc_hd__buf_2
Xhold126 hold51/X vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__buf_2
Xhold115 hold130/X vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__buf_2
Xhold159 hold177/X vssd1 vssd1 vccd1 vccd1 _3971_/A sky130_fd_sc_hd__buf_2
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__buf_2
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__buf_2
Xfanout606 _3584_/A0 vssd1 vssd1 vccd1 vccd1 _3611_/A1 sky130_fd_sc_hd__buf_4
X_4374_ _5736_/Q _4370_/X _4374_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4374_/X sky130_fd_sc_hd__o211a_1
Xfanout617 _5320_/Q vssd1 vssd1 vccd1 vccd1 _2849_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout628 _5290_/Q vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__buf_6
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3325_ _3325_/A _3325_/B vssd1 vssd1 vccd1 vccd1 _3325_/X sky130_fd_sc_hd__or2_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 _3732_/B vssd1 vssd1 vccd1 vccd1 _3729_/B sky130_fd_sc_hd__buf_6
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _5577_/Q _5593_/Q _3284_/S vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3187_ _3240_/S _3186_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3187_/X sky130_fd_sc_hd__a21o_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold682 hold682/A vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__buf_2
XFILLER_104_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2050 _3960_/X vssd1 vssd1 vccd1 vccd1 hold2050/X sky130_fd_sc_hd__buf_2
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1360 hold2695/X vssd1 vssd1 vccd1 vccd1 hold2696/A sky130_fd_sc_hd__buf_2
Xhold2083 hold445/X vssd1 vssd1 vccd1 vccd1 hold2083/X sky130_fd_sc_hd__buf_2
Xhold1393 hold2152/X vssd1 vssd1 vccd1 vccd1 hold2153/A sky130_fd_sc_hd__buf_2
Xhold1382 hold522/X vssd1 vssd1 vccd1 vccd1 _5069_/D sky130_fd_sc_hd__buf_2
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876__461 _4892__477/A vssd1 vssd1 vccd1 vccd1 _5597_/CLK sky130_fd_sc_hd__inv_2
Xoutput209 _3672_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5243_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3110_ _5356_/Q _3605_/A1 _3111_/S vssd1 vssd1 vccd1 vccd1 _5356_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4090_ _5691_/Q _4094_/C vssd1 vssd1 vccd1 vccd1 _4090_/X sky130_fd_sc_hd__and2_1
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3041_ _5027_/Q _3041_/A2 _3041_/B1 _3040_/X vssd1 vssd1 vccd1 vccd1 _3041_/X sky130_fd_sc_hd__o22a_1
XFILLER_95_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4992_ _5243_/CLK _4992_/D vssd1 vssd1 vccd1 vccd1 _4992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _3943_/A0 _5100_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3874_ _4369_/A _3871_/X _3873_/X _4361_/A vssd1 vssd1 vccd1 vccd1 _3874_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5613_ _5613_/CLK _5613_/D vssd1 vssd1 vccd1 vccd1 _5613_/Q sky130_fd_sc_hd__dfxtp_1
X_2825_ _3562_/A _2852_/A vssd1 vssd1 vccd1 vccd1 _2833_/S sky130_fd_sc_hd__or2_4
XFILLER_136_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5544_ _5546_/CLK _5544_/D vssd1 vssd1 vccd1 vccd1 _5544_/Q sky130_fd_sc_hd__dfxtp_2
X_2756_ _3395_/A0 _5474_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5474_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2687_ _3601_/A1 _5536_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5536_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5475_ _5475_/CLK _5475_/D vssd1 vssd1 vccd1 vccd1 _5475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout414 _3672_/B vssd1 vssd1 vccd1 vccd1 _3663_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout436 _2863_/Y vssd1 vssd1 vccd1 vccd1 _3099_/A sky130_fd_sc_hd__clkbuf_4
Xfanout447 _3619_/Y vssd1 vssd1 vccd1 vccd1 _3728_/S sky130_fd_sc_hd__buf_6
Xfanout425 _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3923_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4357_ _4357_/A _4357_/B _4357_/C vssd1 vssd1 vccd1 vccd1 _4357_/X sky130_fd_sc_hd__and3_1
XFILLER_140_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4288_ _5663_/Q _4269_/B _5664_/Q vssd1 vssd1 vccd1 vccd1 _4288_/X sky130_fd_sc_hd__a21o_1
X_3308_ _3308_/A1 _3159_/B _3307_/X _4093_/B vssd1 vssd1 vccd1 vccd1 _5338_/D sky130_fd_sc_hd__o211a_1
Xfanout469 _3301_/A1 vssd1 vssd1 vccd1 vccd1 _3328_/A sky130_fd_sc_hd__buf_4
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3239_ _3171_/A _3238_/X _3235_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3239_/X sky130_fd_sc_hd__a211o_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4710__295 _5002_/CLK vssd1 vssd1 vccd1 vccd1 _5401_/CLK sky130_fd_sc_hd__inv_2
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4460__45 _4460__45/A vssd1 vssd1 vccd1 vccd1 _5054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3590_ _5033_/Q _3590_/A1 _3597_/S vssd1 vssd1 vccd1 vccd1 _5033_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2610_ _3567_/A1 _5610_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5610_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2541_ _3568_/A1 _5702_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5702_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _5261_/CLK _5260_/D vssd1 vssd1 vccd1 vccd1 _5260_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2472_ _3346_/A _3344_/A _5335_/Q vssd1 vssd1 vccd1 vccd1 _3406_/A sky130_fd_sc_hd__or3b_4
XFILLER_114_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4653__238 _5726_/CLK vssd1 vssd1 vccd1 vccd1 _5339_/CLK sky130_fd_sc_hd__inv_2
X_4211_ _4209_/Y _4210_/X _4217_/A vssd1 vssd1 vccd1 vccd1 _5551_/D sky130_fd_sc_hd__a21oi_1
XFILLER_141_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5191_ _5191_/CLK _5191_/D vssd1 vssd1 vccd1 vccd1 _5191_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2819 _4089_/X vssd1 vssd1 vccd1 vccd1 hold2819/X sky130_fd_sc_hd__buf_2
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4142_ _5753_/Q _4142_/B _4142_/C vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__and3_1
XFILLER_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4073_ _4042_/X _4073_/B _4073_/C _4073_/D vssd1 vssd1 vccd1 vccd1 _4074_/C sky130_fd_sc_hd__and4b_1
XFILLER_56_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3024_ _5450_/Q _5568_/Q _3024_/S vssd1 vssd1 vccd1 vccd1 _3024_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_84_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4960__545/A sky130_fd_sc_hd__clkbuf_16
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i _4676__261/A vssd1 vssd1 vccd1 vccd1 _5731_/CLK sky130_fd_sc_hd__clkbuf_16
X_4547__132 _4419__4/A vssd1 vssd1 vccd1 vccd1 _5189_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4975_ _4975_/CLK _4975_/D vssd1 vssd1 vccd1 vccd1 _4975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3926_ _5087_/Q _3926_/A2 _3901_/X vssd1 vssd1 vccd1 vccd1 _5087_/D sky130_fd_sc_hd__a21o_1
XFILLER_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3857_ _3888_/A _3857_/B vssd1 vssd1 vccd1 vccd1 _3857_/Y sky130_fd_sc_hd__nor2_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2808_ _3536_/A0 _5432_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5432_/D sky130_fd_sc_hd__mux2_1
X_3788_ _3789_/A1 _5020_/Q _3829_/A _3796_/B1 _4988_/Q vssd1 vssd1 vccd1 vccd1 _3788_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_117_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5527_ _5527_/CLK _5527_/D vssd1 vssd1 vccd1 vccd1 _5527_/Q sky130_fd_sc_hd__dfxtp_1
X_2739_ _3339_/A1 _5489_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5489_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _5458_/CLK _5458_/D vssd1 vssd1 vccd1 vccd1 _5458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4409_ _5752_/Q _4409_/B vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__or2_1
X_5389_ _5389_/CLK _5389_/D vssd1 vssd1 vccd1 vccd1 _5389_/Q sky130_fd_sc_hd__dfxtp_1
X_4505__90 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5147_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3711_ _4990_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__or2_1
X_3642_ _3642_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3642_/X sky130_fd_sc_hd__or2_1
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5312_ _5312_/CLK _5312_/D vssd1 vssd1 vccd1 vccd1 _5312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3573_ _3573_/A0 _5048_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5048_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2524_ _5335_/Q _3344_/A _3346_/A vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__or3_4
X_2455_ _5550_/Q vssd1 vssd1 vccd1 vccd1 _2455_/Y sky130_fd_sc_hd__inv_2
X_5243_ _5243_/CLK _5243_/D vssd1 vssd1 vccd1 vccd1 _5243_/Q sky130_fd_sc_hd__dfxtp_1
X_5174_ _5174_/CLK _5174_/D vssd1 vssd1 vccd1 vccd1 _5174_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2627 hold2627/A vssd1 vssd1 vccd1 vccd1 hold2627/X sky130_fd_sc_hd__buf_2
Xhold2605 hold2605/A vssd1 vssd1 vccd1 vccd1 hold2605/X sky130_fd_sc_hd__buf_2
Xhold2638 hold2638/A vssd1 vssd1 vccd1 vccd1 hold2638/X sky130_fd_sc_hd__buf_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__buf_2
Xhold1926 hold2768/X vssd1 vssd1 vccd1 vccd1 hold1926/X sky130_fd_sc_hd__buf_2
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1904 hold2756/X vssd1 vssd1 vccd1 vccd1 hold1904/X sky130_fd_sc_hd__buf_2
Xhold1915 hold2760/X vssd1 vssd1 vccd1 vccd1 hold1915/X sky130_fd_sc_hd__buf_2
X_4125_ _5545_/Q _5544_/Q _5543_/Q _4132_/B vssd1 vssd1 vccd1 vccd1 _4128_/B sky130_fd_sc_hd__nand4_2
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1948 hold2764/X vssd1 vssd1 vccd1 vccd1 hold1948/X sky130_fd_sc_hd__buf_2
Xhold1937 hold2772/X vssd1 vssd1 vccd1 vccd1 hold1937/X sky130_fd_sc_hd__buf_2
X_4056_ _5755_/Q _5665_/Q vssd1 vssd1 vccd1 vccd1 _4056_/X sky130_fd_sc_hd__xor2_1
X_3007_ _3099_/B _3005_/X _3006_/X vssd1 vssd1 vccd1 vccd1 _3007_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4781__366 _4909__494/A vssd1 vssd1 vccd1 vccd1 _5472_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4430__15 _4470__55/A vssd1 vssd1 vccd1 vccd1 _4981_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3909_ _5078_/Q _3926_/A2 _3923_/B1 _3908_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5078_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4675__260 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5364_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput370 _5934_/X vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_12
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput381 _3742_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__clkbuf_2
Xoutput392 _3766_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4916__501 _4453__38/A vssd1 vssd1 vccd1 vccd1 _5637_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4496__81 _4504__89/A vssd1 vssd1 vccd1 vccd1 _5138_/CLK sky130_fd_sc_hd__inv_2
XFILLER_120_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5930_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5930_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5861_ _5861_/A vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4659__244 _4432__17/A vssd1 vssd1 vccd1 vccd1 _5347_/CLK sky130_fd_sc_hd__inv_2
XFILLER_147_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3625_ hold90/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3625_/X sky130_fd_sc_hd__and2_1
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3556_ _5063_/Q _3601_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5063_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2507_ _5100_/Q _5101_/Q _5102_/Q _5099_/Q vssd1 vssd1 vccd1 vccd1 _2512_/D sky130_fd_sc_hd__or4b_4
XFILLER_130_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput109 probe_out[76] vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__clkbuf_2
X_5226_ _5226_/CLK _5226_/D vssd1 vssd1 vccd1 vccd1 _5226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3487_ _3595_/A1 _5172_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5172_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2402 hold2402/A vssd1 vssd1 vccd1 vccd1 hold2402/X sky130_fd_sc_hd__buf_2
Xhold2413 hold21/X vssd1 vssd1 vccd1 vccd1 hold2413/X sky130_fd_sc_hd__buf_2
X_2438_ _5681_/Q vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__inv_2
Xhold2446 hold2446/A vssd1 vssd1 vccd1 vccd1 input138/A sky130_fd_sc_hd__buf_2
Xhold2424 hold2424/A vssd1 vssd1 vccd1 vccd1 hold998/A sky130_fd_sc_hd__buf_2
Xhold2435 hold2435/A vssd1 vssd1 vccd1 vccd1 hold2435/X sky130_fd_sc_hd__buf_2
Xhold1701 hold2365/X vssd1 vssd1 vccd1 vccd1 hold2366/A sky130_fd_sc_hd__buf_2
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5157_ _5157_/CLK _5157_/D vssd1 vssd1 vccd1 vccd1 _5157_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1712 hold2232/X vssd1 vssd1 vccd1 vccd1 hold2233/A sky130_fd_sc_hd__buf_2
Xhold2457 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 hold2457/X sky130_fd_sc_hd__buf_2
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5088_ _5111_/CLK _5088_/D vssd1 vssd1 vccd1 vccd1 _5088_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1745 hold2551/X vssd1 vssd1 vccd1 vccd1 hold2552/A sky130_fd_sc_hd__buf_2
Xhold1756 hold2568/X vssd1 vssd1 vccd1 vccd1 hold2569/A sky130_fd_sc_hd__buf_2
X_4108_ _5549_/Q _4108_/B _4119_/C _4108_/D vssd1 vssd1 vccd1 vccd1 _4114_/B sky130_fd_sc_hd__nand4_4
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1789 hold2523/X vssd1 vssd1 vccd1 vccd1 hold2524/A sky130_fd_sc_hd__buf_2
X_4039_ _4052_/B _4052_/C vssd1 vssd1 vccd1 vccd1 _4039_/X sky130_fd_sc_hd__or2_2
XFILLER_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_60 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 hold90/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XCaravelHost_704 vssd1 vssd1 vccd1 vccd1 CaravelHost_704/HI manufacturerID[4] sky130_fd_sc_hd__conb_1
XFILLER_7_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_715 vssd1 vssd1 vccd1 vccd1 CaravelHost_715/HI partID[9] sky130_fd_sc_hd__conb_1
XCaravelHost_726 vssd1 vssd1 vccd1 vccd1 partID[6] CaravelHost_726/LO sky130_fd_sc_hd__conb_1
Xhold308 hold328/X vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__buf_2
Xhold319 hold319/A vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__buf_2
X_4390_ _4390_/A _4390_/B _4390_/C vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__or3_1
X_3410_ _5270_/Q _3566_/A1 _3414_/S vssd1 vssd1 vccd1 vccd1 _5270_/D sky130_fd_sc_hd__mux2_1
X_3341_ _3346_/A _3349_/A vssd1 vssd1 vccd1 vccd1 _3347_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3334_/A1 _3249_/X _3252_/X _3271_/X _3169_/B vssd1 vssd1 vccd1 vccd1 _3272_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5011_ _5262_/CLK _5011_/D vssd1 vssd1 vccd1 vccd1 _5011_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1019 hold1604/X vssd1 vssd1 vccd1 vccd1 hold1605/A sky130_fd_sc_hd__buf_2
XFILLER_94_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1008 hold1570/X vssd1 vssd1 vccd1 vccd1 hold1571/A sky130_fd_sc_hd__buf_2
XFILLER_39_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _5913_/A vssd1 vssd1 vccd1 vccd1 _5913_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5844_ _5844_/A vssd1 vssd1 vccd1 vccd1 _5844_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2987_ _5212_/Q _5148_/Q _3036_/S vssd1 vssd1 vccd1 vccd1 _2987_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4893__478 _4901__486/A vssd1 vssd1 vccd1 vccd1 _5614_/CLK sky130_fd_sc_hd__inv_2
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3608_ _4974_/Q _3608_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4974_/D sky130_fd_sc_hd__mux2_1
Xinput91 probe_out[5] vssd1 vssd1 vccd1 vccd1 _5842_/A sky130_fd_sc_hd__clkbuf_2
Xinput80 probe_out[4] vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__clkbuf_2
Xhold853 hold853/A vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__buf_2
Xhold842 hold842/A vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__buf_2
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3539_ _3584_/A0 _5126_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5126_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold875 hold875/A vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__buf_2
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2221 hold2221/A vssd1 vssd1 vccd1 vccd1 _5324_/D sky130_fd_sc_hd__buf_2
XFILLER_130_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2232 hold2232/A vssd1 vssd1 vccd1 vccd1 hold2232/X sky130_fd_sc_hd__buf_2
XFILLER_85_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5209_ _5731_/CLK _5209_/D vssd1 vssd1 vccd1 vccd1 _5209_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2254 hold2254/A vssd1 vssd1 vccd1 vccd1 hold963/A sky130_fd_sc_hd__buf_2
Xhold2243 hold2243/A vssd1 vssd1 vccd1 vccd1 hold957/A sky130_fd_sc_hd__buf_2
XFILLER_123_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2287 hold2287/A vssd1 vssd1 vccd1 vccd1 _5383_/D sky130_fd_sc_hd__buf_2
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1542 hold7/X vssd1 vssd1 vccd1 vccd1 hold988/A sky130_fd_sc_hd__buf_2
Xhold1520 _3938_/X vssd1 vssd1 vccd1 vccd1 hold983/A sky130_fd_sc_hd__buf_2
Xhold1531 hold994/X vssd1 vssd1 vccd1 vccd1 _3939_/A0 sky130_fd_sc_hd__buf_2
Xhold2265 hold2265/A vssd1 vssd1 vccd1 vccd1 hold969/A sky130_fd_sc_hd__buf_2
Xhold1553 hold999/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__buf_2
X_4787__372 _5697_/CLK vssd1 vssd1 vccd1 vccd1 _5478_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1575 hold2435/X vssd1 vssd1 vccd1 vccd1 hold2436/A sky130_fd_sc_hd__buf_2
Xhold1586 hold2443/X vssd1 vssd1 vccd1 vccd1 hold2444/A sky130_fd_sc_hd__buf_2
Xhold1564 hold2417/X vssd1 vssd1 vccd1 vccd1 hold2418/A sky130_fd_sc_hd__buf_2
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1597 hold2459/X vssd1 vssd1 vccd1 vccd1 hold2460/A sky130_fd_sc_hd__buf_2
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4466__51 _4469__54/A vssd1 vssd1 vccd1 vccd1 _5060_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2910_ _5128_/Q _5160_/Q _5316_/Q _5361_/Q _2941_/S0 _3072_/S vssd1 vssd1 vccd1 vccd1
+ _2910_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3890_ _3844_/A _3955_/A _5072_/Q hold554/X vssd1 vssd1 vccd1 vccd1 _3890_/X sky130_fd_sc_hd__a31o_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2841_ _2850_/A1 _5402_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5402_/D sky130_fd_sc_hd__mux2_1
X_4580__165 _4477__62/A vssd1 vssd1 vccd1 vccd1 _5230_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5560_ _5726_/CLK _5560_/D vssd1 vssd1 vccd1 vccd1 _5560_/Q sky130_fd_sc_hd__dfxtp_1
X_2772_ _3393_/A0 _5460_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5460_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4468__53/A
+ sky130_fd_sc_hd__clkbuf_16
X_5491_ _5491_/CLK _5491_/D vssd1 vssd1 vccd1 vccd1 _5491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold105 hold123/X vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__buf_2
Xhold116 hold132/X vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__buf_2
XFILLER_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__buf_2
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__buf_2
XFILLER_125_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4373_ _3648_/A _3778_/B _4370_/X vssd1 vssd1 vccd1 vccd1 _4373_/X sky130_fd_sc_hd__a21bo_1
Xfanout607 _3593_/A1 vssd1 vssd1 vccd1 vccd1 _3602_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout618 _5319_/Q vssd1 vssd1 vccd1 vccd1 _3596_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout629 _3920_/B vssd1 vssd1 vccd1 vccd1 _3924_/B sky130_fd_sc_hd__buf_4
X_3324_ _5521_/Q _5274_/Q _3324_/S vssd1 vssd1 vccd1 vccd1 _3325_/B sky130_fd_sc_hd__mux2_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3325_/A _3253_/X _3254_/X _3320_/C1 vssd1 vssd1 vccd1 vccd1 _3255_/X sky130_fd_sc_hd__o211a_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3186_ _5414_/Q _5390_/Q _5660_/Q _5422_/Q _3327_/S _3219_/S0 vssd1 vssd1 vccd1 vccd1
+ _3186_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4821__406 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5512_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5689_ _5691_/CLK _5689_/D vssd1 vssd1 vccd1 vccd1 _5689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4715__300 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5406_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold672 hold873/X vssd1 vssd1 vccd1 vccd1 hold874/A sky130_fd_sc_hd__buf_2
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2051 hold2051/A vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__buf_2
Xhold2040 hold2688/X vssd1 vssd1 vccd1 vccd1 hold2689/A sky130_fd_sc_hd__buf_2
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1361 hold2058/X vssd1 vssd1 vccd1 vccd1 hold2059/A sky130_fd_sc_hd__buf_2
Xhold2095 _3788_/X vssd1 vssd1 vccd1 vccd1 hold2095/X sky130_fd_sc_hd__buf_2
Xhold2084 hold2084/A vssd1 vssd1 vccd1 vccd1 _4986_/D sky130_fd_sc_hd__buf_2
XFILLER_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1394 hold2154/X vssd1 vssd1 vccd1 vccd1 hold2155/A sky130_fd_sc_hd__buf_2
Xhold1372 hold2125/X vssd1 vssd1 vccd1 vccd1 hold2126/A sky130_fd_sc_hd__buf_2
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4564__149 _4508__93/A vssd1 vssd1 vccd1 vccd1 _5214_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3040_ _5171_/Q _5235_/Q _3040_/S vssd1 vssd1 vccd1 vccd1 _3040_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _5243_/CLK _4991_/D vssd1 vssd1 vccd1 vccd1 _4991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3942_ _3942_/A0 _5099_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3942_/X sky130_fd_sc_hd__mux2_1
X_3873_ _5732_/Q _3857_/Y _3872_/X _3887_/B _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3873_/X
+ sky130_fd_sc_hd__a221o_1
X_5612_ _5612_/CLK _5612_/D vssd1 vssd1 vccd1 vccd1 _5612_/Q sky130_fd_sc_hd__dfxtp_1
X_2824_ _5692_/Q _5417_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5417_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5543_ _5543_/CLK _5543_/D vssd1 vssd1 vccd1 vccd1 _5543_/Q sky130_fd_sc_hd__dfxtp_4
X_2755_ _3394_/A0 _5475_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5475_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2686_ _3600_/A1 _5537_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5537_/D sky130_fd_sc_hd__mux2_1
X_5474_ _5474_/CLK _5474_/D vssd1 vssd1 vccd1 vccd1 _5474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4356_ _4356_/A _4357_/B _4357_/C vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__and3_1
Xfanout415 _3622_/Y vssd1 vssd1 vccd1 vccd1 _3672_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout448 _3619_/Y vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__buf_6
Xfanout437 _2778_/A vssd1 vssd1 vccd1 vccd1 _3080_/B1 sky130_fd_sc_hd__buf_4
Xfanout426 _3845_/Y vssd1 vssd1 vccd1 vccd1 _3925_/B1 sky130_fd_sc_hd__buf_6
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3307_ _5338_/Q _3125_/A _3156_/X _3306_/X vssd1 vssd1 vccd1 vccd1 _3307_/X sky130_fd_sc_hd__a211o_1
XFILLER_140_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4287_ _4269_/Y _4286_/Y _4285_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5663_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3238_ _5476_/Q _3331_/A2 _3328_/A _3236_/X _3237_/X vssd1 vssd1 vccd1 vccd1 _3238_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3169_ _3357_/A _3169_/B vssd1 vssd1 vccd1 vccd1 _3169_/Y sky130_fd_sc_hd__nand2_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4899__484 _4901__486/A vssd1 vssd1 vccd1 vccd1 _5620_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold480 hold501/X vssd1 vssd1 vccd1 vccd1 hold502/A sky130_fd_sc_hd__buf_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4436__21 _5730_/CLK vssd1 vssd1 vccd1 vccd1 _5030_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2540_ _3576_/A0 _5703_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5703_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4692__277 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5381_/CLK sky130_fd_sc_hd__inv_2
X_4210_ _4210_/A _4210_/B _4210_/C vssd1 vssd1 vccd1 vccd1 _4210_/X sky130_fd_sc_hd__or3_1
X_5190_ _5190_/CLK _5190_/D vssd1 vssd1 vccd1 vccd1 _5190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4141_ _4142_/B _4142_/C vssd1 vssd1 vccd1 vccd1 _4141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4072_ _5742_/Q _4270_/B _4070_/Y _4071_/X vssd1 vssd1 vccd1 vccd1 _4073_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3023_ _5115_/Q _3041_/A2 _2945_/A _3022_/X vssd1 vssd1 vccd1 vccd1 _3043_/C sky130_fd_sc_hd__o211a_1
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4586__171 _4439__24/A vssd1 vssd1 vccd1 vccd1 _5236_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4974_ _4974_/CLK _4974_/D vssd1 vssd1 vccd1 vccd1 _4974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5252_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3925_ _5086_/Q _2490_/X _3925_/B1 _3924_/X _3901_/X vssd1 vssd1 vccd1 vccd1 _5086_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3856_ _3998_/A1 _5202_/Q _3882_/A3 _3855_/X vssd1 vssd1 vccd1 vccd1 _3856_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2807_ _3589_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2815_/S sky130_fd_sc_hd__or2_4
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3787_ _3789_/A1 _5019_/Q _3829_/A _3796_/B1 _4987_/Q vssd1 vssd1 vccd1 vccd1 _3787_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_133_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5526_ _5526_/CLK _5526_/D vssd1 vssd1 vccd1 vccd1 _5526_/Q sky130_fd_sc_hd__dfxtp_1
X_2738_ _3308_/A1 _5490_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5490_/D sky130_fd_sc_hd__mux2_1
X_4933__518 _4455__40/A vssd1 vssd1 vccd1 vccd1 _5654_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5457_ _5457_/CLK _5457_/D vssd1 vssd1 vccd1 vccd1 _5457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4408_ _5751_/Q _4415_/A3 _4407_/X _4368_/A vssd1 vssd1 vccd1 vccd1 _4408_/X sky130_fd_sc_hd__o211a_1
X_2669_ _5578_/Q _3576_/A0 _2672_/S vssd1 vssd1 vccd1 vccd1 _5578_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5388_ _5388_/CLK _5388_/D vssd1 vssd1 vccd1 vccd1 _5388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4339_ _5687_/Q _4324_/X _4338_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5686_/D sky130_fd_sc_hd__o211a_1
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827__412 _5019_/CLK vssd1 vssd1 vccd1 vccd1 _5518_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3710_ _5073_/Q input32/X _3728_/S vssd1 vssd1 vccd1 vccd1 _3710_/X sky130_fd_sc_hd__mux2_4
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4620__205 _4965__550/A vssd1 vssd1 vccd1 vccd1 _5297_/CLK sky130_fd_sc_hd__inv_2
XFILLER_146_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3641_ _4389_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__or2_1
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3572_ _3572_/A0 _5049_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _5049_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5311_ _5311_/CLK _5311_/D vssd1 vssd1 vccd1 vccd1 _5311_/Q sky130_fd_sc_hd__dfxtp_1
X_2523_ _3579_/A0 _5716_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5716_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2454_ _5556_/Q vssd1 vssd1 vccd1 vccd1 _2454_/Y sky130_fd_sc_hd__inv_2
X_5242_ _5243_/CLK _5242_/D vssd1 vssd1 vccd1 vccd1 _5242_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_100_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5248_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5173_ _5173_/CLK _5173_/D vssd1 vssd1 vccd1 vccd1 _5173_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2628 hold2628/A vssd1 vssd1 vccd1 vccd1 hold459/A sky130_fd_sc_hd__buf_2
Xhold2617 _4356_/X vssd1 vssd1 vccd1 vccd1 hold2617/X sky130_fd_sc_hd__buf_2
Xhold2606 hold2606/A vssd1 vssd1 vccd1 vccd1 hold2606/X sky130_fd_sc_hd__buf_2
Xhold1927 hold1927/A vssd1 vssd1 vccd1 vccd1 hold589/A sky130_fd_sc_hd__buf_2
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1905 hold1905/A vssd1 vssd1 vccd1 vccd1 hold857/A sky130_fd_sc_hd__buf_2
Xhold1916 hold1916/A vssd1 vssd1 vccd1 vccd1 hold852/A sky130_fd_sc_hd__buf_2
X_4124_ _5544_/Q _5543_/Q _4132_/B vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__nand3_1
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1949 hold1949/A vssd1 vssd1 vccd1 vccd1 hold803/A sky130_fd_sc_hd__buf_2
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1938 hold1938/A vssd1 vssd1 vccd1 vccd1 hold862/A sky130_fd_sc_hd__buf_2
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4055_ _5754_/Q _4258_/B vssd1 vssd1 vccd1 vccd1 _4055_/X sky130_fd_sc_hd__xor2_1
X_3006_ _2867_/A _5188_/Q _2866_/B _5196_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3006_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3908_ _5743_/Q _3924_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3908_/X sky130_fd_sc_hd__and3_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3839_ _5557_/Q _3835_/X _3834_/X _5529_/Q vssd1 vssd1 vccd1 vccd1 _3839_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5509_ _5509_/CLK _5509_/D vssd1 vssd1 vccd1 vccd1 _5509_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput360 _5925_/X vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_12
XFILLER_10_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput371 _5846_/X vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_12
XFILLER_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput382 _3745_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput393 _3768_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4955__540 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5713_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5860_ _5860_/A vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3624_ _3624_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3624_/X sky130_fd_sc_hd__and2_1
X_4698__283 _5246_/CLK vssd1 vssd1 vccd1 vccd1 _5389_/CLK sky130_fd_sc_hd__inv_2
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3555_ _5064_/Q _3600_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5064_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2506_ _5107_/Q _5108_/Q _5109_/Q _5110_/Q vssd1 vssd1 vccd1 vccd1 _2512_/C sky130_fd_sc_hd__or4_4
XFILLER_130_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3486_ _3594_/A1 _5173_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5173_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5225_ _5225_/CLK _5225_/D vssd1 vssd1 vccd1 vccd1 _5225_/Q sky130_fd_sc_hd__dfxtp_1
X_2437_ _5683_/Q vssd1 vssd1 vccd1 vccd1 _4080_/A sky130_fd_sc_hd__inv_2
Xhold2403 hold2403/A vssd1 vssd1 vccd1 vccd1 hold2403/X sky130_fd_sc_hd__buf_2
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2436 hold2436/A vssd1 vssd1 vccd1 vccd1 input160/A sky130_fd_sc_hd__buf_2
Xhold2425 hold998/X vssd1 vssd1 vccd1 vccd1 hold2425/X sky130_fd_sc_hd__buf_2
Xhold2414 hold2414/A vssd1 vssd1 vccd1 vccd1 hold2414/X sky130_fd_sc_hd__buf_2
Xhold1702 hold2367/X vssd1 vssd1 vccd1 vccd1 hold2368/A sky130_fd_sc_hd__buf_2
XFILLER_111_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _5156_/CLK _5156_/D vssd1 vssd1 vccd1 vccd1 _5156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1735 hold2832/X vssd1 vssd1 vccd1 vccd1 hold2281/A sky130_fd_sc_hd__buf_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2447 _3673_/A vssd1 vssd1 vccd1 vccd1 hold2447/X sky130_fd_sc_hd__buf_2
Xhold2458 hold2458/A vssd1 vssd1 vccd1 vccd1 hold2458/X sky130_fd_sc_hd__buf_2
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5087_ _5684_/CLK _5087_/D vssd1 vssd1 vccd1 vccd1 _5087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1746 hold2553/X vssd1 vssd1 vccd1 vccd1 hold2554/A sky130_fd_sc_hd__buf_2
X_4107_ _5740_/Q _4107_/B vssd1 vssd1 vccd1 vccd1 _4177_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4038_ _4065_/B _4029_/C _5673_/Q vssd1 vssd1 vccd1 vccd1 _4052_/C sky130_fd_sc_hd__a21oi_1
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4939__524 _5246_/CLK vssd1 vssd1 vccd1 vccd1 _5660_/CLK sky130_fd_sc_hd__inv_2
XANTENNA_50 _3628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_61 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_83 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_716 vssd1 vssd1 vccd1 vccd1 CaravelHost_716/HI partID[12] sky130_fd_sc_hd__conb_1
XCaravelHost_727 vssd1 vssd1 vccd1 vccd1 partID[8] CaravelHost_727/LO sky130_fd_sc_hd__conb_1
XCaravelHost_705 vssd1 vssd1 vccd1 vccd1 CaravelHost_705/HI manufacturerID[5] sky130_fd_sc_hd__conb_1
XFILLER_144_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold309 hold318/X vssd1 vssd1 vccd1 vccd1 hold319/A sky130_fd_sc_hd__buf_2
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3340_ _5336_/Q _5345_/Q _3350_/B _4091_/A vssd1 vssd1 vccd1 vccd1 _5336_/D sky130_fd_sc_hd__o211a_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4732__317 _5246_/CLK vssd1 vssd1 vccd1 vccd1 _5423_/CLK sky130_fd_sc_hd__inv_2
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5010_ _5010_/CLK _5010_/D vssd1 vssd1 vccd1 vccd1 _5010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3266_/X _3267_/X _3270_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3271_/X sky130_fd_sc_hd__a211o_1
XFILLER_94_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1009 hold2430/X vssd1 vssd1 vccd1 vccd1 hold2431/A sky130_fd_sc_hd__buf_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5912_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5912_/X sky130_fd_sc_hd__clkbuf_4
X_4626__211 _5564_/CLK vssd1 vssd1 vccd1 vccd1 _5303_/CLK sky130_fd_sc_hd__inv_2
X_5843_ _5843_/A vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2986_ _3594_/A1 _2895_/Y _2985_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5378_/D sky130_fd_sc_hd__o211a_1
XFILLER_147_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3607_ _3607_/A _3607_/B vssd1 vssd1 vccd1 vccd1 _3615_/S sky130_fd_sc_hd__nor2_8
Xinput81 probe_out[50] vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__clkbuf_2
Xinput70 probe_out[40] vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__clkbuf_2
Xhold810 hold810/A vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__buf_2
Xhold821 hold821/A vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__buf_2
Xinput92 probe_out[60] vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__clkbuf_2
X_3538_ _3538_/A0 _5127_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5127_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3469_ _5188_/Q _3613_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5188_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2233 hold2233/A vssd1 vssd1 vccd1 vccd1 _5325_/D sky130_fd_sc_hd__buf_2
XFILLER_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _5731_/CLK _5208_/D vssd1 vssd1 vccd1 vccd1 _5208_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1510 hold32/X vssd1 vssd1 vccd1 vccd1 hold978/A sky130_fd_sc_hd__buf_2
Xhold2244 hold957/X vssd1 vssd1 vccd1 vccd1 hold2244/X sky130_fd_sc_hd__buf_2
Xhold2255 hold963/X vssd1 vssd1 vccd1 vccd1 hold2255/X sky130_fd_sc_hd__buf_2
X_5139_ _5139_/CLK _5139_/D vssd1 vssd1 vccd1 vccd1 _5139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1543 hold988/X vssd1 vssd1 vccd1 vccd1 _3940_/A0 sky130_fd_sc_hd__buf_2
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1532 _3939_/X vssd1 vssd1 vccd1 vccd1 hold995/A sky130_fd_sc_hd__buf_2
Xhold1521 hold983/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__buf_2
Xhold2266 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 hold2266/X sky130_fd_sc_hd__buf_2
Xhold2288 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 hold2288/X sky130_fd_sc_hd__buf_2
Xhold1554 hold16/X vssd1 vssd1 vccd1 vccd1 hold1554/X sky130_fd_sc_hd__buf_2
Xhold1576 hold2437/X vssd1 vssd1 vccd1 vccd1 hold2438/A sky130_fd_sc_hd__buf_2
Xhold1565 hold1565/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__buf_2
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5752_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1598 hold2461/X vssd1 vssd1 vccd1 vccd1 hold2462/A sky130_fd_sc_hd__buf_2
Xhold1587 hold2445/X vssd1 vssd1 vccd1 vccd1 hold2446/A sky130_fd_sc_hd__buf_2
XFILLER_16_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4481__66 _5004_/CLK vssd1 vssd1 vccd1 vccd1 _5123_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _2849_/A1 _5403_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5403_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2771_ _3392_/A0 _5461_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5461_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5490_ _5490_/CLK _5490_/D vssd1 vssd1 vccd1 vccd1 _5490_/Q sky130_fd_sc_hd__dfxtp_1
Xhold117 hold52/X vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__buf_2
Xhold106 hold127/X vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__buf_2
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold139 _3781_/Y vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_78_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4460__45/A sky130_fd_sc_hd__clkbuf_16
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__buf_2
XFILLER_125_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4372_ _5735_/Q _4370_/X _4372_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4372_/X sky130_fd_sc_hd__o211a_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _5319_/Q vssd1 vssd1 vccd1 vccd1 _3614_/A1 sky130_fd_sc_hd__buf_2
XFILLER_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout608 _3584_/A0 vssd1 vssd1 vccd1 vccd1 _3593_/A1 sky130_fd_sc_hd__buf_6
X_3323_ _3357_/B _3321_/X _3322_/X _3323_/C1 vssd1 vssd1 vccd1 vccd1 _3323_/X sky130_fd_sc_hd__o211a_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _5649_/Q _3331_/A2 _3128_/B _5641_/Q vssd1 vssd1 vccd1 vccd1 _3254_/X sky130_fd_sc_hd__o22a_1
XFILLER_67_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3185_ _3355_/B _3185_/B vssd1 vssd1 vccd1 vccd1 _3185_/X sky130_fd_sc_hd__and2_1
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4860__445 _4892__477/A vssd1 vssd1 vccd1 vccd1 _5581_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2969_ _2867_/A _5189_/Q _3041_/A2 _5197_/Q _3064_/C1 vssd1 vssd1 vccd1 vccd1 _2969_/X
+ sky130_fd_sc_hd__o221a_1
X_4901__486 _4901__486/A vssd1 vssd1 vccd1 vccd1 _5622_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5688_ _5691_/CLK _5688_/D vssd1 vssd1 vccd1 vccd1 _5688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold662 hold662/A vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__buf_2
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold673 hold710/X vssd1 vssd1 vccd1 vccd1 hold711/A sky130_fd_sc_hd__buf_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2030 hold2030/A vssd1 vssd1 vccd1 vccd1 _4990_/D sky130_fd_sc_hd__buf_2
XFILLER_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2052 hold200/X vssd1 vssd1 vccd1 vccd1 hold2052/X sky130_fd_sc_hd__buf_2
Xhold2041 hold2690/X vssd1 vssd1 vccd1 vccd1 hold2691/A sky130_fd_sc_hd__buf_2
XFILLER_94_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2096 hold2096/A vssd1 vssd1 vccd1 vccd1 hold449/A sky130_fd_sc_hd__buf_2
Xhold2074 hold2713/X vssd1 vssd1 vccd1 vccd1 hold2714/A sky130_fd_sc_hd__buf_2
Xhold1340 hold2675/X vssd1 vssd1 vccd1 vccd1 hold2030/A sky130_fd_sc_hd__buf_2
Xhold1395 hold2156/X vssd1 vssd1 vccd1 vccd1 hold2157/A sky130_fd_sc_hd__buf_2
Xhold1373 hold2127/X vssd1 vssd1 vccd1 vccd1 hold2128/A sky130_fd_sc_hd__buf_2
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4844__429 _4468__53/A vssd1 vssd1 vccd1 vccd1 _5537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4990_ _5243_/CLK _4990_/D vssd1 vssd1 vccd1 vccd1 _4990_/Q sky130_fd_sc_hd__dfxtp_1
X_3941_ _3941_/A0 _5098_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3941_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3872_ _4401_/A _5205_/Q _3897_/C _3855_/X vssd1 vssd1 vccd1 vccd1 _3872_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5611_ _5611_/CLK _5611_/D vssd1 vssd1 vccd1 vccd1 _5611_/Q sky130_fd_sc_hd__dfxtp_1
X_2823_ _3395_/A0 _5418_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5418_/D sky130_fd_sc_hd__mux2_1
X_5542_ _5542_/CLK _5542_/D vssd1 vssd1 vccd1 vccd1 _5542_/Q sky130_fd_sc_hd__dfxtp_1
X_2754_ _3402_/A1 _5476_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5476_/D sky130_fd_sc_hd__mux2_1
X_4738__323 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5429_/CLK sky130_fd_sc_hd__inv_2
X_2685_ _3599_/A1 _5538_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5538_/D sky130_fd_sc_hd__mux2_1
X_5473_ _5473_/CLK _5473_/D vssd1 vssd1 vccd1 vccd1 _5473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4355_ _4355_/A split5/X _4357_/C vssd1 vssd1 vccd1 vccd1 _4355_/X sky130_fd_sc_hd__and3_1
Xfanout416 _3622_/Y vssd1 vssd1 vccd1 vccd1 _3682_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout438 _4088_/B vssd1 vssd1 vccd1 vccd1 _2778_/A sky130_fd_sc_hd__buf_6
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout427 _4204_/A vssd1 vssd1 vccd1 vccd1 _4217_/A sky130_fd_sc_hd__buf_4
X_3306_ _3303_/X _3305_/X _3357_/A vssd1 vssd1 vccd1 vccd1 _3306_/X sky130_fd_sc_hd__o21a_1
Xfanout449 _3619_/Y vssd1 vssd1 vccd1 vccd1 _3773_/B sky130_fd_sc_hd__clkbuf_4
X_4286_ _5663_/Q _4286_/B vssd1 vssd1 vccd1 vccd1 _4286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _5711_/Q _3237_/B vssd1 vssd1 vccd1 vccd1 _3237_/X sky130_fd_sc_hd__or2_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3168_ _3316_/C1 _3165_/X _3167_/X vssd1 vssd1 vccd1 vccd1 _3168_/X sky130_fd_sc_hd__a21o_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3099_ _3099_/A _3099_/B vssd1 vssd1 vccd1 vccd1 _3099_/Y sky130_fd_sc_hd__nand2_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold481 hold503/X vssd1 vssd1 vccd1 vccd1 hold504/A sky130_fd_sc_hd__buf_2
Xhold470 _4404_/X vssd1 vssd1 vccd1 vccd1 _5749_/D sky130_fd_sc_hd__buf_2
XFILLER_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531__116 _4435__20/A vssd1 vssd1 vccd1 vccd1 _5173_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1170 hold1845/X vssd1 vssd1 vccd1 vccd1 hold1846/A sky130_fd_sc_hd__buf_2
XFILLER_58_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1192 hold2563/X vssd1 vssd1 vccd1 vccd1 hold2564/A sky130_fd_sc_hd__buf_2
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451__36 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5045_/CLK sky130_fd_sc_hd__inv_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2470_ _5384_/Q vssd1 vssd1 vccd1 vccd1 _2863_/A sky130_fd_sc_hd__inv_2
XFILLER_142_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4140_ _5540_/Q _5539_/Q _5541_/Q vssd1 vssd1 vccd1 vccd1 _4142_/C sky130_fd_sc_hd__a21o_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4071_ _5745_/Q _4071_/B _4071_/C vssd1 vssd1 vccd1 vccd1 _4071_/X sky130_fd_sc_hd__and3_1
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3022_ _5227_/Q _2870_/B _3021_/X _3041_/B1 vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__o22a_1
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4973_ _4973_/CLK _4973_/D vssd1 vssd1 vccd1 vccd1 _4973_/Q sky130_fd_sc_hd__dfxtp_1
X_3924_ _5735_/Q _3924_/B _5292_/Q vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__and3_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3855_ _3888_/C _3855_/B vssd1 vssd1 vccd1 vccd1 _3855_/X sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_93_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4455__40/A
+ sky130_fd_sc_hd__clkbuf_16
X_2806_ _5433_/Q _3543_/A0 _2806_/S vssd1 vssd1 vccd1 vccd1 _5433_/D sky130_fd_sc_hd__mux2_1
X_3786_ _3789_/A1 _5018_/Q _3829_/A _3796_/B1 _4986_/Q vssd1 vssd1 vccd1 vccd1 _3786_/X
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4478__63/A
+ sky130_fd_sc_hd__clkbuf_16
X_5525_ _5525_/CLK _5525_/D vssd1 vssd1 vccd1 vccd1 _5525_/Q sky130_fd_sc_hd__dfxtp_1
X_2737_ _3277_/A1 _5491_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5491_/D sky130_fd_sc_hd__mux2_1
X_5456_ _5456_/CLK _5456_/D vssd1 vssd1 vccd1 vccd1 _5456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2668_ _5579_/Q _3575_/A0 _2672_/S vssd1 vssd1 vccd1 vccd1 _5579_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4407_ _4354_/A split5/A _4415_/A3 vssd1 vssd1 vccd1 vccd1 _4407_/X sky130_fd_sc_hd__a21bo_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2599_ _2743_/A0 _5620_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5620_/D sky130_fd_sc_hd__mux2_1
X_5387_ _5387_/CLK _5387_/D vssd1 vssd1 vccd1 vccd1 _5387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4338_ _5686_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4338_/X sky130_fd_sc_hd__or2_1
XFILLER_115_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4269_ _4269_/A _4269_/B vssd1 vssd1 vccd1 vccd1 _4269_/Y sky130_fd_sc_hd__nor2_1
X_4866__451 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5587_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4907__492 _5022_/CLK vssd1 vssd1 vccd1 vccd1 _5628_/CLK sky130_fd_sc_hd__inv_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3640_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3640_/X sky130_fd_sc_hd__or2_1
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4700__285 _5246_/CLK vssd1 vssd1 vccd1 vccd1 _5391_/CLK sky130_fd_sc_hd__inv_2
X_3571_ _3571_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _3579_/S sky130_fd_sc_hd__or2_4
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5310_ _5310_/CLK _5310_/D vssd1 vssd1 vccd1 vccd1 _5310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2522_ _3569_/A1 _5717_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5717_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5241_ _5241_/CLK _5241_/D vssd1 vssd1 vccd1 vccd1 _5241_/Q sky130_fd_sc_hd__dfxtp_1
X_2453_ _5665_/Q vssd1 vssd1 vccd1 vccd1 _2453_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5172_ _5172_/CLK _5172_/D vssd1 vssd1 vccd1 vccd1 _5172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2629 hold459/X vssd1 vssd1 vccd1 vccd1 hold2629/X sky130_fd_sc_hd__buf_2
Xhold2618 hold2618/A vssd1 vssd1 vccd1 vccd1 hold2618/X sky130_fd_sc_hd__buf_2
Xhold2607 hold2607/A vssd1 vssd1 vccd1 vccd1 hold782/A sky130_fd_sc_hd__buf_2
Xhold1906 hold857/X vssd1 vssd1 vccd1 vccd1 hold1906/X sky130_fd_sc_hd__buf_2
Xhold1917 hold852/X vssd1 vssd1 vccd1 vccd1 hold1917/X sky130_fd_sc_hd__buf_2
X_4123_ _4122_/B _4122_/C _5747_/Q vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__a21oi_2
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
Xhold1928 hold589/X vssd1 vssd1 vccd1 vccd1 hold1928/X sky130_fd_sc_hd__buf_2
XFILLER_84_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4054_ _5666_/Q _5665_/Q vssd1 vssd1 vccd1 vccd1 _4258_/B sky130_fd_sc_hd__xnor2_4
XFILLER_69_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1939 hold862/X vssd1 vssd1 vccd1 vccd1 hold1939/X sky130_fd_sc_hd__buf_2
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3005_ _4969_/Q _5180_/Q _3005_/S vssd1 vssd1 vccd1 vccd1 _3005_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3907_ _5077_/Q _3926_/A2 _3923_/B1 _3906_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5077_/D
+ sky130_fd_sc_hd__a221o_1
X_3838_ _5530_/Q _5529_/Q vssd1 vssd1 vccd1 vccd1 _4181_/B sky130_fd_sc_hd__or2_4
XFILLER_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3769_ _3769_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__and2_1
X_5508_ _5508_/CLK _5508_/D vssd1 vssd1 vccd1 vccd1 _5508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5439_ _5439_/CLK _5439_/D vssd1 vssd1 vccd1 vccd1 _5439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput361 _5926_/X vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_12
Xoutput350 _5916_/X vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_12
XFILLER_102_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput372 _3777_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_12
Xoutput383 _3748_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput394 _3770_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643__228 _4658__243/A vssd1 vssd1 vccd1 vccd1 _5329_/CLK sky130_fd_sc_hd__inv_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4537__122 _4418__3/A vssd1 vssd1 vccd1 vccd1 _5179_/CLK sky130_fd_sc_hd__inv_2
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3623_ _3623_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3623_/X sky130_fd_sc_hd__and2_1
XFILLER_135_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3554_ _5065_/Q _3599_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5065_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2505_ _5103_/Q _5104_/Q _5105_/Q _5106_/Q vssd1 vssd1 vccd1 vccd1 _2512_/B sky130_fd_sc_hd__or4_4
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3485_ _3593_/A1 _5174_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5174_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5224_ _5224_/CLK _5224_/D vssd1 vssd1 vccd1 vccd1 _5224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2436_ _5738_/Q vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__inv_2
Xhold2404 hold2404/A vssd1 vssd1 vccd1 vccd1 hold903/A sky130_fd_sc_hd__buf_2
XFILLER_130_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2437 _3664_/A vssd1 vssd1 vccd1 vccd1 hold2437/X sky130_fd_sc_hd__buf_2
Xhold2426 hold2426/A vssd1 vssd1 vccd1 vccd1 input137/A sky130_fd_sc_hd__buf_2
Xhold2415 hold2415/A vssd1 vssd1 vccd1 vccd1 hold2415/X sky130_fd_sc_hd__buf_2
X_5155_ _5155_/CLK _5155_/D vssd1 vssd1 vccd1 vccd1 _5155_/Q sky130_fd_sc_hd__dfxtp_1
X_4487__72 _5262_/CLK vssd1 vssd1 vccd1 vccd1 _5129_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1703 hold2369/X vssd1 vssd1 vccd1 vccd1 hold2370/A sky130_fd_sc_hd__buf_2
Xhold2459 hold2459/A vssd1 vssd1 vccd1 vccd1 hold2459/X sky130_fd_sc_hd__buf_2
Xhold2448 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 hold2448/X sky130_fd_sc_hd__buf_2
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1736 hold2282/X vssd1 vssd1 vccd1 vccd1 hold2283/A sky130_fd_sc_hd__buf_2
XFILLER_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5086_ _5738_/CLK _5086_/D vssd1 vssd1 vccd1 vccd1 _5086_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1747 hold2555/X vssd1 vssd1 vccd1 vccd1 hold2556/A sky130_fd_sc_hd__buf_2
X_4106_ _5554_/Q _4153_/B vssd1 vssd1 vccd1 vccd1 _4107_/B sky130_fd_sc_hd__xor2_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4037_ _4041_/B _4041_/C _4253_/A vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__a21oi_1
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_40 _3185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_62 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 _3355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_717 vssd1 vssd1 vccd1 vccd1 CaravelHost_717/HI partID[13] sky130_fd_sc_hd__conb_1
XCaravelHost_728 vssd1 vssd1 vccd1 vccd1 partID[10] CaravelHost_728/LO sky130_fd_sc_hd__conb_1
XCaravelHost_706 vssd1 vssd1 vccd1 vccd1 CaravelHost_706/HI manufacturerID[6] sky130_fd_sc_hd__conb_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4771__356 _5697_/CLK vssd1 vssd1 vccd1 vccd1 _5462_/CLK sky130_fd_sc_hd__inv_2
XFILLER_125_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _3328_/A _3268_/X _3269_/X _3171_/A vssd1 vssd1 vccd1 vccd1 _3270_/X sky130_fd_sc_hd__o211a_1
XFILLER_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4812__397 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5503_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5911_ _5911_/A vssd1 vssd1 vccd1 vccd1 _5911_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4665__250 _4477__62/A vssd1 vssd1 vccd1 vccd1 _5353_/CLK sky130_fd_sc_hd__inv_2
X_5842_ _5842_/A vssd1 vssd1 vccd1 vccd1 _5842_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4706__291 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5397_/CLK sky130_fd_sc_hd__inv_2
X_2985_ _2863_/A _5378_/Q _3094_/A _2984_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _2985_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3606_ _4975_/Q _3606_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4975_/D sky130_fd_sc_hd__mux2_1
Xinput82 probe_out[51] vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__clkbuf_2
Xinput71 probe_out[41] vssd1 vssd1 vccd1 vccd1 _5878_/A sky130_fd_sc_hd__clkbuf_2
Xinput60 probe_out[31] vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__clkbuf_2
Xinput93 probe_out[61] vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__clkbuf_2
X_3537_ _3600_/A1 _5128_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5128_/D sky130_fd_sc_hd__mux2_1
Xhold833 hold833/A vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__buf_2
Xhold822 hold822/A vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__buf_2
XFILLER_143_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3468_ _5189_/Q _3612_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5189_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5207_ _5730_/CLK _5207_/D vssd1 vssd1 vccd1 vccd1 _5207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3399_ _5280_/Q _3564_/A1 _3405_/S vssd1 vssd1 vccd1 vccd1 _5280_/D sky130_fd_sc_hd__mux2_1
Xhold1500 hold2266/X vssd1 vssd1 vccd1 vccd1 hold2267/A sky130_fd_sc_hd__buf_2
Xhold2245 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 hold2245/X sky130_fd_sc_hd__buf_2
Xhold2234 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 hold2234/X sky130_fd_sc_hd__buf_2
X_5138_ _5138_/CLK _5138_/D vssd1 vssd1 vccd1 vccd1 _5138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1544 _3940_/X vssd1 vssd1 vccd1 vccd1 hold989/A sky130_fd_sc_hd__buf_2
Xhold1522 hold29/X vssd1 vssd1 vccd1 vccd1 hold984/A sky130_fd_sc_hd__buf_2
Xhold1533 hold995/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__buf_2
Xhold1511 hold978/X vssd1 vssd1 vccd1 vccd1 _5094_/D sky130_fd_sc_hd__buf_2
Xhold2267 hold2267/A vssd1 vssd1 vccd1 vccd1 hold973/A sky130_fd_sc_hd__buf_2
Xhold2256 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 hold2256/X sky130_fd_sc_hd__buf_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1555 hold1555/A vssd1 vssd1 vccd1 vccd1 _3941_/A0 sky130_fd_sc_hd__buf_2
Xhold1566 hold22/X vssd1 vssd1 vccd1 vccd1 hold1566/X sky130_fd_sc_hd__buf_2
Xhold2289 hold2289/A vssd1 vssd1 vccd1 vccd1 hold979/A sky130_fd_sc_hd__buf_2
Xhold1577 hold1577/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__buf_2
X_5069_ _5755_/CLK _5069_/D vssd1 vssd1 vccd1 vccd1 _5069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1599 hold2463/X vssd1 vssd1 vccd1 vccd1 hold2464/A sky130_fd_sc_hd__buf_2
Xhold1588 hold2447/X vssd1 vssd1 vccd1 vccd1 hold1588/X sky130_fd_sc_hd__buf_2
XFILLER_38_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2790 hold2790/A vssd1 vssd1 vccd1 vccd1 hold2790/X sky130_fd_sc_hd__buf_2
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4649__234 _5248_/CLK vssd1 vssd1 vccd1 vccd1 _5335_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2770_ _3409_/A1 _5462_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5462_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 hold131/X vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__buf_2
XFILLER_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__buf_2
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__buf_2
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4371_ _3649_/A _3778_/B _4370_/X vssd1 vssd1 vccd1 vccd1 _4371_/X sky130_fd_sc_hd__a21bo_1
XFILLER_125_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout609 _5322_/Q vssd1 vssd1 vccd1 vccd1 _3584_/A0 sky130_fd_sc_hd__buf_8
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3322_ _5700_/Q _2464_/Y _3326_/B2 _5716_/Q vssd1 vssd1 vccd1 vccd1 _3322_/X sky130_fd_sc_hd__o22a_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _5044_/Q _5633_/Q _3284_/S vssd1 vssd1 vccd1 vccd1 _3253_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_47_wb_clk_i clkbuf_4_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5001_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _5713_/Q _5462_/Q _5446_/Q _5478_/Q _3299_/S _3184_/S1 vssd1 vssd1 vccd1 vccd1
+ _3185_/B sky130_fd_sc_hd__mux4_2
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4457__42 _4457__42/A vssd1 vssd1 vccd1 vccd1 _5051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2968_ _4970_/Q _5181_/Q _3005_/S vssd1 vssd1 vccd1 vccd1 _2968_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5687_ _5691_/CLK _5687_/D vssd1 vssd1 vccd1 vccd1 _5687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2899_ _5144_/Q _5152_/Q _5216_/Q _5136_/Q _3036_/S _2944_/S0 vssd1 vssd1 vccd1 vccd1
+ _2899_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold641 hold641/A vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__buf_2
XFILLER_131_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold696 hold696/A vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__buf_2
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold674 _3929_/X vssd1 vssd1 vccd1 vccd1 _5088_/D sky130_fd_sc_hd__buf_2
XFILLER_131_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2053 hold2053/A vssd1 vssd1 vccd1 vccd1 _5112_/D sky130_fd_sc_hd__buf_2
XFILLER_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2042 hold2042/A vssd1 vssd1 vccd1 vccd1 _4991_/D sky130_fd_sc_hd__buf_2
Xhold1352 hold2655/X vssd1 vssd1 vccd1 vccd1 hold2656/A sky130_fd_sc_hd__buf_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2075 hold2075/A vssd1 vssd1 vccd1 vccd1 hold437/A sky130_fd_sc_hd__buf_2
Xhold2097 hold449/X vssd1 vssd1 vccd1 vccd1 hold2097/X sky130_fd_sc_hd__buf_2
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1374 hold2129/X vssd1 vssd1 vccd1 vccd1 hold2130/A sky130_fd_sc_hd__buf_2
XFILLER_45_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1396 hold561/X vssd1 vssd1 vccd1 vccd1 _5066_/D sky130_fd_sc_hd__buf_2
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4883__468 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5604_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _3940_/A0 _5097_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3940_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3871_ _5752_/Q _4401_/A _3897_/C _3887_/A vssd1 vssd1 vccd1 vccd1 _3871_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5610_ _5610_/CLK _5610_/D vssd1 vssd1 vccd1 vccd1 _5610_/Q sky130_fd_sc_hd__dfxtp_1
X_2822_ _3394_/A0 _5419_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5419_/D sky130_fd_sc_hd__mux2_1
X_5541_ _5542_/CLK _5541_/D vssd1 vssd1 vccd1 vccd1 _5541_/Q sky130_fd_sc_hd__dfxtp_2
X_2753_ _3392_/A0 _5477_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5477_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777__362 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5468_/CLK sky130_fd_sc_hd__inv_2
X_2684_ _3508_/A _3598_/B vssd1 vssd1 vccd1 vccd1 _2692_/S sky130_fd_sc_hd__or2_4
X_5472_ _5472_/CLK _5472_/D vssd1 vssd1 vccd1 vccd1 _5472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4354_ _4354_/A split5/X _4357_/C vssd1 vssd1 vccd1 vccd1 _4354_/X sky130_fd_sc_hd__and3_1
Xfanout417 _3622_/Y vssd1 vssd1 vccd1 vccd1 _3688_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout439 _4094_/C vssd1 vssd1 vccd1 vccd1 _4088_/B sky130_fd_sc_hd__buf_6
Xfanout406 _4278_/X vssd1 vssd1 vccd1 vccd1 _4308_/A2 sky130_fd_sc_hd__buf_4
Xfanout428 hold701/X vssd1 vssd1 vccd1 vccd1 hold702/A sky130_fd_sc_hd__buf_6
X_3305_ _3336_/A1 _3286_/X _3289_/X _3304_/X _3136_/X vssd1 vssd1 vccd1 vccd1 _3305_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4285_ _4318_/A2 _4286_/B _5663_/Q vssd1 vssd1 vccd1 vccd1 _4285_/X sky130_fd_sc_hd__a21o_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _5444_/Q _5460_/Q _3330_/S vssd1 vssd1 vccd1 vccd1 _3236_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3167_ _3320_/C1 _3166_/X _3334_/A1 vssd1 vssd1 vccd1 vccd1 _3167_/X sky130_fd_sc_hd__a21o_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3098_ _2867_/A _3099_/A _3097_/Y _4088_/B vssd1 vssd1 vccd1 vccd1 _5366_/D sky130_fd_sc_hd__o211a_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5739_ _5739_/CLK _5739_/D vssd1 vssd1 vccd1 vccd1 _5739_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold482 hold505/X vssd1 vssd1 vccd1 vccd1 hold506/A sky130_fd_sc_hd__buf_2
Xhold493 hold493/A vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__buf_2
X_4570__155 _4433__18/A vssd1 vssd1 vccd1 vccd1 _5220_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1171 hold1847/X vssd1 vssd1 vccd1 vccd1 hold1848/A sky130_fd_sc_hd__buf_2
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1193 hold2567/X vssd1 vssd1 vccd1 vccd1 hold2568/A sky130_fd_sc_hd__buf_2
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4611__196 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _4071_/B _4071_/C _5745_/Q vssd1 vssd1 vccd1 vccd1 _4070_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3021_ _5163_/Q _5348_/Q _3040_/S vssd1 vssd1 vccd1 vccd1 _3021_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4427__12 _4469__54/A vssd1 vssd1 vccd1 vccd1 _4978_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4972_ _4972_/CLK _4972_/D vssd1 vssd1 vccd1 vccd1 _4972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3923_ _5085_/Q _2490_/X _3923_/B1 _3922_/X _3901_/X vssd1 vssd1 vccd1 vccd1 _5085_/D
+ sky130_fd_sc_hd__a221o_1
X_3854_ _3888_/C _3855_/B vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2805_ _5434_/Q _2850_/A1 _2806_/S vssd1 vssd1 vccd1 vccd1 _5434_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3785_ _4403_/B1 _5017_/Q _3829_/A _3796_/B1 _4985_/Q vssd1 vssd1 vccd1 vccd1 _3785_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5524_ _5524_/CLK _5524_/D vssd1 vssd1 vccd1 vccd1 _5524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2736_ _3567_/A1 _5492_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5492_/D sky130_fd_sc_hd__mux2_1
X_5455_ _5455_/CLK _5455_/D vssd1 vssd1 vccd1 vccd1 _5455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2667_ _5580_/Q _3574_/A0 _2672_/S vssd1 vssd1 vccd1 vccd1 _5580_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4406_ _5750_/Q _4415_/A3 _4405_/X _4368_/A vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__o211a_1
X_4554__139 _4418__3/A vssd1 vssd1 vccd1 vccd1 _5196_/CLK sky130_fd_sc_hd__inv_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2598_ _3573_/A0 _5621_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5621_/D sky130_fd_sc_hd__mux2_1
X_5386_ _5386_/CLK _5386_/D vssd1 vssd1 vccd1 vccd1 _5386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _5686_/Q _4324_/X _4336_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5685_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4268_ _4268_/A _4268_/B _4268_/C _4268_/D vssd1 vssd1 vccd1 vccd1 _4269_/B sky130_fd_sc_hd__and4_2
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3219_ _5626_/Q _5516_/Q _5285_/Q _5468_/Q _3219_/S0 _3330_/S vssd1 vssd1 vccd1 vccd1
+ _3219_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4199_ _5546_/Q _4187_/B1 _4210_/C _4160_/B vssd1 vssd1 vccd1 vccd1 _4200_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4511__96 _4422__7/A vssd1 vssd1 vccd1 vccd1 _5153_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _5050_/Q _3579_/A0 _3570_/S vssd1 vssd1 vccd1 vccd1 _5050_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ _3577_/A0 _5718_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5718_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5240_ _5240_/CLK _5240_/D vssd1 vssd1 vccd1 vccd1 _5240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2452_ _5666_/Q vssd1 vssd1 vccd1 vccd1 _2452_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ _5171_/CLK _5171_/D vssd1 vssd1 vccd1 vccd1 _5171_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2619 hold2619/A vssd1 vssd1 vccd1 vccd1 hold2619/X sky130_fd_sc_hd__buf_2
Xhold2608 hold782/X vssd1 vssd1 vccd1 vccd1 hold2608/X sky130_fd_sc_hd__buf_2
XFILLER_110_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1907 hold1907/A vssd1 vssd1 vccd1 vccd1 _4392_/B1 sky130_fd_sc_hd__buf_2
Xhold1918 hold1918/A vssd1 vssd1 vccd1 vccd1 _4385_/B1 sky130_fd_sc_hd__buf_2
X_4122_ _5747_/Q _4122_/B _4122_/C vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__and3_1
X_4889__474 _4897__482/A vssd1 vssd1 vccd1 vccd1 _5610_/CLK sky130_fd_sc_hd__inv_2
Xhold1929 hold1929/A vssd1 vssd1 vccd1 vccd1 _4376_/B1 sky130_fd_sc_hd__buf_2
X_4053_ _5754_/Q _5665_/Q vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__xnor2_1
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
X_3004_ _2460_/A _5357_/Q _5124_/Q _3073_/B2 _3004_/C1 vssd1 vssd1 vccd1 vccd1 _3004_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3906_ _5744_/Q _3924_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3906_/X sky130_fd_sc_hd__and3_1
X_3837_ _5530_/Q _5529_/Q vssd1 vssd1 vccd1 vccd1 _4186_/A sky130_fd_sc_hd__nor2_8
XFILLER_146_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3768_ _5011_/Q _3774_/A2 _3774_/B1 _3767_/X _3774_/C1 vssd1 vssd1 vccd1 vccd1 _3768_/X
+ sky130_fd_sc_hd__o221a_4
X_2719_ _3277_/A1 _5507_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5507_/D sky130_fd_sc_hd__mux2_1
X_5507_ _5507_/CLK _5507_/D vssd1 vssd1 vccd1 vccd1 _5507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3699_ _4986_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3699_/X sky130_fd_sc_hd__or2_1
X_5438_ _5438_/CLK _5438_/D vssd1 vssd1 vccd1 vccd1 _5438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput362 _5845_/X vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_12
Xoutput351 _5844_/X vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_12
Xoutput340 _5843_/X vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_12
XFILLER_114_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5369_ _5369_/CLK _5369_/D vssd1 vssd1 vccd1 vccd1 _5369_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput384 _3694_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput395 _3697_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput373 _3691_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4682__267 _4425__10/A vssd1 vssd1 vccd1 vccd1 _5371_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4576__161 _4432__17/A vssd1 vssd1 vccd1 vccd1 _5226_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4923__508 _4453__38/A vssd1 vssd1 vccd1 vccd1 _5644_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3622_ _3659_/B vssd1 vssd1 vccd1 vccd1 _3622_/Y sky130_fd_sc_hd__inv_2
X_4817__402 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5508_/CLK sky130_fd_sc_hd__inv_2
X_3553_ _3589_/A _3598_/B vssd1 vssd1 vccd1 vccd1 _3561_/S sky130_fd_sc_hd__nor2_8
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3484_ _3592_/A1 _5175_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5175_/D sky130_fd_sc_hd__mux2_1
X_2504_ _5091_/Q _5092_/Q _3851_/B vssd1 vssd1 vccd1 vccd1 _4399_/C sky130_fd_sc_hd__or3_4
XFILLER_142_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2435_ _5739_/Q vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__inv_2
X_5223_ _5223_/CLK _5223_/D vssd1 vssd1 vccd1 vccd1 _5223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ _5154_/CLK _5154_/D vssd1 vssd1 vccd1 vccd1 _5154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2405 hold903/X vssd1 vssd1 vccd1 vccd1 hold2405/X sky130_fd_sc_hd__buf_2
Xhold2427 _3672_/A vssd1 vssd1 vccd1 vccd1 hold2427/X sky130_fd_sc_hd__buf_2
Xhold2416 hold2416/A vssd1 vssd1 vccd1 vccd1 input157/A sky130_fd_sc_hd__buf_2
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ _5553_/Q _5552_/Q _4210_/A vssd1 vssd1 vccd1 vccd1 _4153_/B sky130_fd_sc_hd__nand3_4
Xhold1704 hold2371/X vssd1 vssd1 vccd1 vccd1 hold2372/A sky130_fd_sc_hd__buf_2
Xhold2449 hold2449/A vssd1 vssd1 vccd1 vccd1 hold2449/X sky130_fd_sc_hd__buf_2
Xhold2438 hold2438/A vssd1 vssd1 vccd1 vccd1 hold2438/X sky130_fd_sc_hd__buf_2
X_5085_ _5684_/CLK _5085_/D vssd1 vssd1 vccd1 vccd1 _5085_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1737 hold2284/X vssd1 vssd1 vccd1 vccd1 hold2285/A sky130_fd_sc_hd__buf_2
X_4036_ _4041_/B _4041_/C vssd1 vssd1 vccd1 vccd1 _4264_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _3543_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _3213_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_74 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _2916_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_718 vssd1 vssd1 vccd1 vccd1 CaravelHost_718/HI versionID[0] sky130_fd_sc_hd__conb_1
XCaravelHost_729 vssd1 vssd1 vccd1 vccd1 partID[11] CaravelHost_729/LO sky130_fd_sc_hd__conb_1
XCaravelHost_707 vssd1 vssd1 vccd1 vccd1 CaravelHost_707/HI manufacturerID[7] sky130_fd_sc_hd__conb_1
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4909__494/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5910_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5841_ _5841_/A vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__clkbuf_4
X_2984_ _3094_/B _2980_/X _2981_/X _2983_/X vssd1 vssd1 vccd1 vccd1 _2984_/X sky130_fd_sc_hd__a31o_1
XFILLER_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput72 probe_out[42] vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__clkbuf_2
X_3605_ _4976_/Q _3605_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4976_/D sky130_fd_sc_hd__mux2_1
Xinput61 probe_out[32] vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__clkbuf_2
Xinput50 probe_out[22] vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__clkbuf_2
Xinput94 probe_out[62] vssd1 vssd1 vccd1 vccd1 _5899_/A sky130_fd_sc_hd__clkbuf_2
Xinput83 probe_out[52] vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__clkbuf_2
X_3536_ _3536_/A0 _5129_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5129_/D sky130_fd_sc_hd__mux2_1
Xhold823 hold823/A vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__buf_2
Xhold867 hold867/A vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__buf_2
X_3467_ _5190_/Q _3611_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5190_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2202 hold2825/X vssd1 vssd1 vccd1 vccd1 hold2826/A sky130_fd_sc_hd__buf_2
XFILLER_88_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5206_ _5730_/CLK _5206_/D vssd1 vssd1 vccd1 vccd1 _5206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3398_ _5281_/Q _3572_/A0 _3405_/S vssd1 vssd1 vccd1 vccd1 _5281_/D sky130_fd_sc_hd__mux2_1
Xhold1501 hold2268/X vssd1 vssd1 vccd1 vccd1 hold2269/A sky130_fd_sc_hd__buf_2
Xhold2235 hold2235/A vssd1 vssd1 vccd1 vccd1 hold955/A sky130_fd_sc_hd__buf_2
Xhold2246 hold2246/A vssd1 vssd1 vccd1 vccd1 hold961/A sky130_fd_sc_hd__buf_2
X_5137_ _5137_/CLK _5137_/D vssd1 vssd1 vccd1 vccd1 _5137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1523 hold984/X vssd1 vssd1 vccd1 vccd1 _5095_/D sky130_fd_sc_hd__buf_2
Xhold1534 hold38/X vssd1 vssd1 vccd1 vccd1 hold996/A sky130_fd_sc_hd__buf_2
Xhold2257 hold2257/A vssd1 vssd1 vccd1 vccd1 hold967/A sky130_fd_sc_hd__buf_2
Xhold1512 hold2288/X vssd1 vssd1 vccd1 vccd1 hold2289/A sky130_fd_sc_hd__buf_2
Xhold2268 hold973/X vssd1 vssd1 vccd1 vccd1 hold2268/X sky130_fd_sc_hd__buf_2
Xhold1545 hold989/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__buf_2
Xhold1556 _3941_/X vssd1 vssd1 vccd1 vccd1 hold1556/X sky130_fd_sc_hd__buf_2
Xhold1567 hold1567/A vssd1 vssd1 vccd1 vccd1 _3932_/A0 sky130_fd_sc_hd__buf_2
X_5068_ _5733_/CLK _5068_/D vssd1 vssd1 vccd1 vccd1 _5068_/Q sky130_fd_sc_hd__dfxtp_1
X_4945__530 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5703_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4019_ _4247_/B _4247_/C _4024_/A vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__a21oi_1
Xhold1578 hold40/X vssd1 vssd1 vccd1 vccd1 hold1578/X sky130_fd_sc_hd__buf_2
Xhold1589 hold1589/A vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__buf_2
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4794__379 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5485_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4688__273 _5384_/CLK vssd1 vssd1 vccd1 vccd1 _5377_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2791 hold2791/A vssd1 vssd1 vccd1 vccd1 hold2791/X sky130_fd_sc_hd__buf_2
XFILLER_75_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 hold117/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__buf_2
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold119 hold134/X vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__buf_2
X_4370_ _5292_/Q _4381_/B vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__and2_4
X_3321_ _5266_/Q _5293_/Q _3324_/S vssd1 vssd1 vccd1 vccd1 _3321_/X sky130_fd_sc_hd__mux2_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _5625_/Q _3237_/B _3171_/A _3251_/X vssd1 vssd1 vccd1 vccd1 _3252_/X sky130_fd_sc_hd__o211a_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3181_/X _3182_/X _3240_/S vssd1 vssd1 vccd1 vccd1 _3183_/X sky130_fd_sc_hd__mux2_1
X_4929__514 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5650_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_87_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4449__34/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4472__57 _4472__57/A vssd1 vssd1 vccd1 vccd1 _5114_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_16_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5384_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2967_ _5061_/Q _3073_/B2 _3029_/B1 _2966_/X vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__o211a_1
X_5755_ _5755_/CLK _5755_/D vssd1 vssd1 vccd1 vccd1 _5755_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2898_ _5120_/Q _5168_/Q _5353_/Q _5232_/Q _2944_/S0 _3040_/S vssd1 vssd1 vccd1 vccd1
+ _2898_/X sky130_fd_sc_hd__mux4_1
X_5686_ _5735_/CLK _5686_/D vssd1 vssd1 vccd1 vccd1 _5686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3519_ _5144_/Q _3609_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5144_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold675 hold675/A vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__buf_2
XFILLER_131_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2021 hold2654/X vssd1 vssd1 vccd1 vccd1 hold2655/A sky130_fd_sc_hd__buf_2
Xhold2010 hold2662/X vssd1 vssd1 vccd1 vccd1 hold2663/A sky130_fd_sc_hd__buf_2
XFILLER_131_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2043 wbs_stb_i vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__buf_2
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 hold2642/X vssd1 vssd1 vccd1 vccd1 hold2643/A sky130_fd_sc_hd__buf_2
Xhold2076 hold437/X vssd1 vssd1 vccd1 vccd1 hold2076/X sky130_fd_sc_hd__buf_2
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1375 hold494/X vssd1 vssd1 vccd1 vccd1 _5067_/D sky130_fd_sc_hd__buf_2
Xhold1386 hold2143/X vssd1 vssd1 vccd1 vccd1 hold2144/A sky130_fd_sc_hd__buf_2
Xhold1353 hold2659/X vssd1 vssd1 vccd1 vccd1 hold2024/A sky130_fd_sc_hd__buf_2
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2098 hold2098/A vssd1 vssd1 vccd1 vccd1 _4988_/D sky130_fd_sc_hd__buf_2
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4722__307 _4731__316/A vssd1 vssd1 vccd1 vccd1 _5413_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4616__201 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5293_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3870_ _5068_/Q _3959_/A _3870_/B1 vssd1 vssd1 vccd1 vccd1 _3870_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2821_ _3393_/A0 _5420_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5420_/D sky130_fd_sc_hd__mux2_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5540_ _5566_/CLK _5540_/D vssd1 vssd1 vccd1 vccd1 _5540_/Q sky130_fd_sc_hd__dfxtp_4
X_2752_ _3391_/A0 _5478_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5478_/D sky130_fd_sc_hd__mux2_1
X_5471_ _5471_/CLK _5471_/D vssd1 vssd1 vccd1 vccd1 _5471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2683_ _3443_/B _3453_/C _5373_/Q vssd1 vssd1 vccd1 vccd1 _3598_/B sky130_fd_sc_hd__or3b_4
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4353_ _4353_/A split5/X _4357_/C vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__and3_1
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout407 _4278_/X vssd1 vssd1 vccd1 vccd1 _4318_/A2 sky130_fd_sc_hd__clkbuf_4
X_4284_ _4281_/X _4322_/B _4283_/X _4279_/X vssd1 vssd1 vccd1 vccd1 _4286_/B sky130_fd_sc_hd__o211a_1
Xfanout429 hold741/X vssd1 vssd1 vccd1 vccd1 hold742/A sky130_fd_sc_hd__buf_4
Xfanout418 _3124_/Y vssd1 vssd1 vccd1 vccd1 _4360_/B sky130_fd_sc_hd__buf_6
X_3304_ _3294_/X _3295_/X _3353_/B _3292_/X vssd1 vssd1 vccd1 vccd1 _3304_/X sky130_fd_sc_hd__a211o_1
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3235_ _3328_/A _3233_/X _3234_/X vssd1 vssd1 vccd1 vccd1 _3235_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3166_ _5645_/Q _5637_/Q _5048_/Q _5653_/Q _3284_/S _3201_/S1 vssd1 vssd1 vccd1 vccd1
+ _3166_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3097_ _3099_/A _3097_/B vssd1 vssd1 vccd1 vccd1 _3097_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3999_ _3971_/A _3914_/C _3999_/S vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__mux2_1
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5738_ _5738_/CLK _5738_/D vssd1 vssd1 vccd1 vccd1 _5738_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5669_ _5731_/CLK _5669_/D vssd1 vssd1 vccd1 vccd1 _5669_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold483 hold483/A vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__buf_2
Xhold494 hold494/A vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__buf_2
XFILLER_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1172 hold1849/X vssd1 vssd1 vccd1 vccd1 hold1850/A sky130_fd_sc_hd__buf_2
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850__435 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5571_/CLK sky130_fd_sc_hd__inv_2
XFILLER_141_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3020_ _3041_/B1 _3018_/X _3019_/X vssd1 vssd1 vccd1 vccd1 _3043_/B sky130_fd_sc_hd__o21a_1
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4971_ _4971_/CLK _4971_/D vssd1 vssd1 vccd1 vccd1 _4971_/Q sky130_fd_sc_hd__dfxtp_1
X_4442__27 _5001_/CLK vssd1 vssd1 vccd1 vccd1 _5036_/CLK sky130_fd_sc_hd__inv_2
X_3922_ _5736_/Q _3924_/B _5292_/Q vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__and3_1
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _3844_/A _3955_/A _3927_/B _3857_/B vssd1 vssd1 vccd1 vccd1 _3887_/B sky130_fd_sc_hd__o31a_4
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2804_ _5435_/Q _2849_/A1 _2806_/S vssd1 vssd1 vccd1 vccd1 _5435_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3784_ _3789_/A1 _5016_/Q _3829_/A _3796_/B1 _4984_/Q vssd1 vssd1 vccd1 vccd1 _3784_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_145_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5523_ _5523_/CLK _5523_/D vssd1 vssd1 vccd1 vccd1 _5523_/Q sky130_fd_sc_hd__dfxtp_1
X_2735_ _3218_/A1 _5493_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5493_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5454_ _5454_/CLK _5454_/D vssd1 vssd1 vccd1 vccd1 _5454_/Q sky130_fd_sc_hd__dfxtp_1
X_2666_ _5581_/Q _3573_/A0 _2672_/S vssd1 vssd1 vccd1 vccd1 _5581_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4405_ _4355_/A split5/A _4415_/A3 vssd1 vssd1 vccd1 vccd1 _4405_/X sky130_fd_sc_hd__a21bo_1
X_5385_ _5385_/CLK _5385_/D vssd1 vssd1 vccd1 vccd1 _5385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4336_ _5685_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4336_/X sky130_fd_sc_hd__or2_1
X_2597_ _3159_/A _5622_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5622_/D sky130_fd_sc_hd__mux2_1
X_4593__178 _4449__34/A vssd1 vssd1 vccd1 vccd1 _5267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4267_ _5743_/Q _4023_/B _4266_/X vssd1 vssd1 vccd1 vccd1 _4268_/D sky130_fd_sc_hd__o21a_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4418__3/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4198_ _4204_/A _4198_/B vssd1 vssd1 vccd1 vccd1 _5545_/D sky130_fd_sc_hd__nor2_1
X_3218_ _3218_/A1 _3159_/B _3217_/X _3277_/C1 vssd1 vssd1 vccd1 vccd1 _5341_/D sky130_fd_sc_hd__o211a_1
X_3149_ _3133_/X _3137_/X _3171_/A vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4834__419 _4460__45/A vssd1 vssd1 vccd1 vccd1 _5525_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 hold352/X vssd1 vssd1 vccd1 vccd1 hold353/A sky130_fd_sc_hd__buf_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__buf_2
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4728__313 _5247_/CLK vssd1 vssd1 vccd1 vccd1 _5419_/CLK sky130_fd_sc_hd__inv_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2520_ _3576_/A0 _5719_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5719_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2451_ _5667_/Q vssd1 vssd1 vccd1 vccd1 _2451_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5170_ _5170_/CLK _5170_/D vssd1 vssd1 vccd1 vccd1 _5170_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2609 hold2609/A vssd1 vssd1 vccd1 vccd1 hold2609/X sky130_fd_sc_hd__buf_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1908 _4392_/X vssd1 vssd1 vccd1 vccd1 hold1908/X sky130_fd_sc_hd__buf_2
X_4121_ _4122_/B _4122_/C vssd1 vssd1 vccd1 vccd1 _4121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4052_ _5747_/Q _4052_/B _4052_/C vssd1 vssd1 vccd1 vccd1 _4275_/B sky130_fd_sc_hd__or3_1
Xhold1919 _4385_/X vssd1 vssd1 vccd1 vccd1 hold1919/X sky130_fd_sc_hd__buf_2
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _3034_/A _3003_/B vssd1 vssd1 vccd1 vccd1 _3003_/X sky130_fd_sc_hd__or2_1
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3905_ _5076_/Q _3926_/A2 _3923_/B1 _3904_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5076_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4521__106 _4433__18/A vssd1 vssd1 vccd1 vccd1 _5163_/CLK sky130_fd_sc_hd__inv_2
X_3836_ _3836_/A _5529_/Q vssd1 vssd1 vccd1 vccd1 _4226_/B sky130_fd_sc_hd__or2_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3767_ _3767_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3767_/X sky130_fd_sc_hd__and2_1
X_2718_ _3567_/A1 _5508_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5508_/D sky130_fd_sc_hd__mux2_1
X_5506_ _5506_/CLK _5506_/D vssd1 vssd1 vccd1 vccd1 _5506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3698_ _5069_/Q input28/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3698_/X sky130_fd_sc_hd__mux2_4
X_5437_ _5437_/CLK _5437_/D vssd1 vssd1 vccd1 vccd1 _5437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput341 _5907_/X vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_12
Xoutput352 _5917_/X vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_12
Xoutput330 _5897_/X vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_12
X_2649_ _5595_/Q _3575_/A0 _2653_/S vssd1 vssd1 vccd1 vccd1 _5595_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5368_ _5368_/CLK _5368_/D vssd1 vssd1 vccd1 vccd1 _5368_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput363 _5927_/X vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_12
Xoutput385 _3751_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput396 _3772_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__clkbuf_2
Xoutput374 _3721_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4319_ _4318_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _5679_/D sky130_fd_sc_hd__and2b_1
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5299_ _5299_/CLK _5299_/D vssd1 vssd1 vccd1 vccd1 _5299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout590 _3339_/A1 vssd1 vssd1 vccd1 vccd1 _3387_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962__547 _4962__547/A vssd1 vssd1 vccd1 vccd1 _5720_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3621_ _3621_/A _3778_/C vssd1 vssd1 vccd1 vccd1 _3621_/X sky130_fd_sc_hd__or2_4
X_3552_ _5114_/Q _3615_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5114_/D sky130_fd_sc_hd__mux2_1
X_4856__441 _4892__477/A vssd1 vssd1 vccd1 vccd1 _5577_/CLK sky130_fd_sc_hd__inv_2
X_2503_ _5093_/Q _5094_/Q _5095_/Q _5096_/Q vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__or4_2
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3483_ _3591_/A1 _5176_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5176_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _5222_/CLK _5222_/D vssd1 vssd1 vccd1 vccd1 _5222_/Q sky130_fd_sc_hd__dfxtp_1
X_2434_ _5741_/Q vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__inv_2
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5153_ _5153_/CLK _5153_/D vssd1 vssd1 vccd1 vccd1 _5153_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2406 hold2406/A vssd1 vssd1 vccd1 vccd1 hold2406/X sky130_fd_sc_hd__buf_2
Xhold2417 _3663_/A vssd1 vssd1 vccd1 vccd1 hold2417/X sky130_fd_sc_hd__buf_2
Xhold2428 hold2428/A vssd1 vssd1 vccd1 vccd1 hold999/A sky130_fd_sc_hd__buf_2
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4104_ _5551_/Q _4108_/B _4119_/C _4104_/D vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__and4_4
Xhold2439 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 hold2439/X sky130_fd_sc_hd__buf_2
X_5084_ _5084_/CLK _5084_/D vssd1 vssd1 vccd1 vccd1 _5084_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1738 hold2286/X vssd1 vssd1 vccd1 vccd1 hold2287/A sky130_fd_sc_hd__buf_2
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1727 hold2401/X vssd1 vssd1 vccd1 vccd1 hold2402/A sky130_fd_sc_hd__buf_2
X_4035_ _5671_/Q _4065_/B _4008_/B _5672_/Q vssd1 vssd1 vccd1 vccd1 _4041_/C sky130_fd_sc_hd__a31o_1
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_20 _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _4390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 _5726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 split2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3819_ _4353_/A _5018_/Q hold80/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__mux2_1
XANTENNA_64 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4599__184 _4965__550/A vssd1 vssd1 vccd1 vccd1 _5273_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4478__63 _4478__63/A vssd1 vssd1 vccd1 vccd1 _5120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XCaravelHost_719 vssd1 vssd1 vccd1 vccd1 CaravelHost_719/HI versionID[1] sky130_fd_sc_hd__conb_1
XCaravelHost_708 vssd1 vssd1 vccd1 vccd1 CaravelHost_708/HI manufacturerID[8] sky130_fd_sc_hd__conb_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2983_ _3045_/A1 _2964_/X _2967_/X _2982_/X _2883_/X vssd1 vssd1 vccd1 vccd1 _2983_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput40 probe_out[13] vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3604_ _4977_/Q _3604_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4977_/D sky130_fd_sc_hd__mux2_1
Xinput73 probe_out[43] vssd1 vssd1 vccd1 vccd1 _5880_/A sky130_fd_sc_hd__clkbuf_2
Xinput62 probe_out[33] vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__clkbuf_2
Xinput51 probe_out[23] vssd1 vssd1 vccd1 vccd1 _5860_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput95 probe_out[63] vssd1 vssd1 vccd1 vccd1 _5900_/A sky130_fd_sc_hd__clkbuf_2
Xinput84 probe_out[53] vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__clkbuf_2
X_3535_ _3589_/A _3535_/B vssd1 vssd1 vccd1 vccd1 _3543_/S sky130_fd_sc_hd__or2_4
Xhold824 hold824/A vssd1 vssd1 vccd1 vccd1 hold824/X sky130_fd_sc_hd__buf_2
X_3466_ _5191_/Q _3610_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5191_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold857 hold857/A vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__buf_2
Xhold868 hold868/A vssd1 vssd1 vccd1 vccd1 hold868/X sky130_fd_sc_hd__buf_2
Xhold879 _2467_/Y vssd1 vssd1 vccd1 vccd1 hold879/X sky130_fd_sc_hd__buf_2
XFILLER_131_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633__218 _5684_/CLK vssd1 vssd1 vccd1 vccd1 _5311_/CLK sky130_fd_sc_hd__inv_2
Xhold2203 hold2203/A vssd1 vssd1 vccd1 vccd1 hold2203/X sky130_fd_sc_hd__buf_2
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5205_ _5384_/CLK _5205_/D vssd1 vssd1 vccd1 vccd1 _5205_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2214 hold2819/X vssd1 vssd1 vccd1 vccd1 hold2820/A sky130_fd_sc_hd__buf_2
X_3397_ _3397_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3405_/S sky130_fd_sc_hd__nor2_8
Xhold2236 hold955/X vssd1 vssd1 vccd1 vccd1 hold2236/X sky130_fd_sc_hd__buf_2
XFILLER_130_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5136_ _5136_/CLK _5136_/D vssd1 vssd1 vccd1 vccd1 _5136_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1535 hold996/X vssd1 vssd1 vccd1 vccd1 _5096_/D sky130_fd_sc_hd__buf_2
Xhold1502 hold2270/X vssd1 vssd1 vccd1 vccd1 hold2271/A sky130_fd_sc_hd__buf_2
Xhold1524 hold2324/X vssd1 vssd1 vccd1 vccd1 hold2325/A sky130_fd_sc_hd__buf_2
Xhold2269 hold2269/A vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__buf_2
Xhold2247 hold961/X vssd1 vssd1 vccd1 vccd1 hold2247/X sky130_fd_sc_hd__buf_2
Xhold2258 hold967/X vssd1 vssd1 vccd1 vccd1 hold2258/X sky130_fd_sc_hd__buf_2
Xhold1513 hold2290/X vssd1 vssd1 vccd1 vccd1 hold2291/A sky130_fd_sc_hd__buf_2
XFILLER_123_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1557 hold1557/A vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__buf_2
Xhold1546 hold8/X vssd1 vssd1 vccd1 vccd1 hold990/A sky130_fd_sc_hd__buf_2
Xhold1568 _3932_/X vssd1 vssd1 vccd1 vccd1 hold1568/X sky130_fd_sc_hd__buf_2
X_5067_ _5733_/CLK _5067_/D vssd1 vssd1 vccd1 vccd1 _5067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4018_ _4247_/B _4247_/C vssd1 vssd1 vccd1 vccd1 _4018_/Y sky130_fd_sc_hd__nand2_1
Xhold1579 hold1579/A vssd1 vssd1 vccd1 vccd1 _3933_/A0 sky130_fd_sc_hd__buf_2
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4527__112 _4509__94/A vssd1 vssd1 vccd1 vccd1 _5169_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2792 hold2792/A vssd1 vssd1 vccd1 vccd1 hold2792/X sky130_fd_sc_hd__buf_2
XFILLER_90_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold109 hold135/X vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__buf_2
XFILLER_113_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3320_ _3325_/A _3318_/X _3319_/X _3320_/C1 vssd1 vssd1 vccd1 vccd1 _3320_/X sky130_fd_sc_hd__o211a_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _5467_/Q _3132_/A _3250_/X _3328_/A vssd1 vssd1 vccd1 vccd1 _3251_/X sky130_fd_sc_hd__o22a_1
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3182_ _5502_/Q _5494_/Q _5486_/Q _5510_/Q _3281_/S _3130_/B vssd1 vssd1 vccd1 vccd1
+ _3182_/X sky130_fd_sc_hd__mux4_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _4744__329/A sky130_fd_sc_hd__clkbuf_16
X_2966_ _4978_/Q _2870_/B _2965_/X _3034_/A vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__o22a_1
X_5754_ _5754_/CLK _5754_/D vssd1 vssd1 vccd1 vccd1 _5754_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2897_ _2897_/A1 _2895_/Y _2896_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5382_/D sky130_fd_sc_hd__o211a_1
X_5685_ _5735_/CLK _5685_/D vssd1 vssd1 vccd1 vccd1 _5685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3518_ _5145_/Q _3590_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5145_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold687 hold821/X vssd1 vssd1 vccd1 vccd1 hold822/A sky130_fd_sc_hd__buf_2
XFILLER_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3449_ _3612_/A1 _5213_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5213_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2000 hold2637/X vssd1 vssd1 vccd1 vccd1 hold2638/A sky130_fd_sc_hd__buf_2
Xhold2011 hold2664/X vssd1 vssd1 vccd1 vccd1 hold2665/A sky130_fd_sc_hd__buf_2
XFILLER_94_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2022 hold2656/X vssd1 vssd1 vccd1 vccd1 hold2657/A sky130_fd_sc_hd__buf_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2033 hold2678/X vssd1 vssd1 vccd1 vccd1 hold2679/A sky130_fd_sc_hd__buf_2
Xhold2044 hold292/X vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__buf_2
X_5119_ _5119_/CLK _5119_/D vssd1 vssd1 vccd1 vccd1 _5119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1332 hold2646/X vssd1 vssd1 vccd1 vccd1 hold2007/A sky130_fd_sc_hd__buf_2
Xhold2077 hold2077/A vssd1 vssd1 vccd1 vccd1 _4987_/D sky130_fd_sc_hd__buf_2
Xhold2088 _3789_/X vssd1 vssd1 vccd1 vccd1 hold2088/X sky130_fd_sc_hd__buf_2
Xhold1343 hold2679/X vssd1 vssd1 vccd1 vccd1 hold2680/A sky130_fd_sc_hd__buf_2
X_4448__33 _4449__34/A vssd1 vssd1 vccd1 vccd1 _5042_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1365 hold2116/X vssd1 vssd1 vccd1 vccd1 hold2117/A sky130_fd_sc_hd__buf_2
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1387 hold2145/X vssd1 vssd1 vccd1 vccd1 hold2146/A sky130_fd_sc_hd__buf_2
XFILLER_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761__346 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5452_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4802__387 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5493_/CLK sky130_fd_sc_hd__inv_2
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4655__240 _4459__44/A vssd1 vssd1 vccd1 vccd1 _5341_/CLK sky130_fd_sc_hd__inv_2
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2820_ _3392_/A0 _5421_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5421_/D sky130_fd_sc_hd__mux2_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2751_ _3390_/A0 _5479_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5479_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2682_ _3615_/A1 _5567_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5567_/D sky130_fd_sc_hd__mux2_1
X_5470_ _5470_/CLK _5470_/D vssd1 vssd1 vccd1 vccd1 _5470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ _4352_/A split5/X _4357_/C vssd1 vssd1 vccd1 vccd1 _4352_/X sky130_fd_sc_hd__and3_1
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout419 _4315_/B vssd1 vssd1 vccd1 vccd1 _4309_/B sky130_fd_sc_hd__clkbuf_4
X_4283_ _5664_/Q _5663_/Q _4283_/C vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__or3_1
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout408 _4186_/X vssd1 vssd1 vccd1 vccd1 _4210_/C sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_103_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5726_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3303_ _3334_/A1 _3280_/X _3283_/X _3302_/X _3169_/B vssd1 vssd1 vccd1 vccd1 _3303_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3234_ _5420_/Q _2482_/B _3237_/B _5412_/Q _3240_/S vssd1 vssd1 vccd1 vccd1 _3234_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3165_ _5613_/Q _5597_/Q _5581_/Q _5621_/Q _3284_/S _3201_/S1 vssd1 vssd1 vccd1 vccd1
+ _3165_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3096_ _5367_/Q _3094_/A _2919_/Y _4088_/B vssd1 vssd1 vccd1 vccd1 _5367_/D sky130_fd_sc_hd__o211a_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ hold97/X _3998_/A1 _3999_/S vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__mux2_1
XFILLER_13_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2949_ _3064_/C1 _2939_/X _3045_/A1 vssd1 vssd1 vccd1 vccd1 _2949_/X sky130_fd_sc_hd__a21o_1
X_5737_ _5738_/CLK _5737_/D vssd1 vssd1 vccd1 vccd1 _5737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4639__224 _4485__70/A vssd1 vssd1 vccd1 vccd1 _5317_/CLK sky130_fd_sc_hd__inv_2
X_5668_ _5731_/CLK _5668_/D vssd1 vssd1 vccd1 vccd1 _5668_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5599_ _5599_/CLK _5599_/D vssd1 vssd1 vccd1 vccd1 _5599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold484 _4323_/X vssd1 vssd1 vccd1 vccd1 _5680_/D sky130_fd_sc_hd__buf_2
XFILLER_131_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1151 hold2215/X vssd1 vssd1 vccd1 vccd1 hold2216/A sky130_fd_sc_hd__buf_2
Xhold1140 hold2406/X vssd1 vssd1 vccd1 vccd1 hold2407/A sky130_fd_sc_hd__buf_2
Xhold1162 hold2731/X vssd1 vssd1 vccd1 vccd1 hold1821/A sky130_fd_sc_hd__buf_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4786__371/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4970_ _4970_/CLK _4970_/D vssd1 vssd1 vccd1 vccd1 _4970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3921_ _5084_/Q _3926_/A2 _3923_/B1 _3920_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5084_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3852_ _3852_/A _3855_/B vssd1 vssd1 vccd1 vccd1 _3927_/B sky130_fd_sc_hd__or2_1
X_2803_ _5436_/Q _2848_/A1 _2806_/S vssd1 vssd1 vccd1 vccd1 _5436_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5522_ _5522_/CLK _5522_/D vssd1 vssd1 vccd1 vccd1 _5522_/Q sky130_fd_sc_hd__dfxtp_1
X_3783_ _3789_/A1 _5015_/Q _3829_/A _3796_/B1 _4983_/Q vssd1 vssd1 vccd1 vccd1 _3783_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2734_ _2743_/A0 _5494_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5494_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5453_ _5453_/CLK _5453_/D vssd1 vssd1 vccd1 vccd1 _5453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2665_ _5582_/Q _3159_/A _2672_/S vssd1 vssd1 vccd1 vccd1 _5582_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5384_ _5384_/CLK _5384_/D vssd1 vssd1 vccd1 vccd1 _5384_/Q sky130_fd_sc_hd__dfxtp_1
X_4404_ _5749_/Q _4401_/Y hold469/X vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__a21o_1
X_2596_ _3370_/A _2664_/B vssd1 vssd1 vccd1 vccd1 _2604_/S sky130_fd_sc_hd__or2_4
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4335_ _5685_/Q _4324_/X _4334_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5684_/D sky130_fd_sc_hd__o211a_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4266_ _5742_/Q _4266_/B vssd1 vssd1 vccd1 vccd1 _4266_/X sky130_fd_sc_hd__xor2_1
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4197_ _5545_/Q _4187_/B1 _4210_/C _4127_/Y vssd1 vssd1 vccd1 vccd1 _4198_/B sky130_fd_sc_hd__o2bb2a_1
X_3217_ _5341_/Q _3125_/A _3353_/A _3216_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3217_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3148_ _3240_/S _3143_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3079_ _3597_/A1 _2895_/Y _3078_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5375_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_71_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5735_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4873__458 _4875__460/A vssd1 vssd1 vccd1 vccd1 _5594_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold270 hold367/X vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__buf_2
Xhold281 hold356/X vssd1 vssd1 vccd1 vccd1 hold357/A sky130_fd_sc_hd__buf_2
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4914__499 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5635_/CLK sky130_fd_sc_hd__inv_2
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__buf_2
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4767__352 _5024_/CLK vssd1 vssd1 vccd1 vccd1 _5458_/CLK sky130_fd_sc_hd__inv_2
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4808__393 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5499_/CLK sky130_fd_sc_hd__inv_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2450_ _5668_/Q vssd1 vssd1 vccd1 vccd1 _2450_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1909 hold1909/A vssd1 vssd1 vccd1 vccd1 hold858/A sky130_fd_sc_hd__buf_2
X_4120_ _4132_/B _4119_/C _5547_/Q vssd1 vssd1 vccd1 vccd1 _4122_/C sky130_fd_sc_hd__a21o_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _4049_/Y _4050_/X _4271_/A _4271_/B vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__o211a_1
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_4502__87 _4510__95/A vssd1 vssd1 vccd1 vccd1 _5144_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3002_ _5156_/Q _5312_/Q _3002_/S vssd1 vssd1 vccd1 vccd1 _3003_/B sky130_fd_sc_hd__mux2_1
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3904_ _5745_/Q _3924_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3904_/X sky130_fd_sc_hd__and3_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4560__145 _4504__89/A vssd1 vssd1 vccd1 vccd1 _5210_/CLK sky130_fd_sc_hd__inv_2
X_3835_ _5562_/Q _5563_/Q _5564_/Q _5565_/Q _5555_/Q _5556_/Q vssd1 vssd1 vccd1 vccd1
+ _3835_/X sky130_fd_sc_hd__mux4_2
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3766_ _5010_/Q _3774_/A2 _3774_/B1 _3765_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3766_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4601__186 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5275_/CLK sky130_fd_sc_hd__inv_2
X_2717_ _3218_/A1 _5509_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5509_/D sky130_fd_sc_hd__mux2_1
X_5505_ _5505_/CLK _5505_/D vssd1 vssd1 vccd1 vccd1 _5505_/Q sky130_fd_sc_hd__dfxtp_1
X_5436_ _5436_/CLK _5436_/D vssd1 vssd1 vccd1 vccd1 _5436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3697_ _3718_/A1 _3695_/X _3696_/X split2/X vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__o211a_2
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput353 _5918_/X vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_12
Xoutput342 _5908_/X vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_12
Xoutput331 _5898_/X vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_12
Xoutput320 _5888_/X vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_12
X_2648_ _5596_/Q _2743_/A0 _2653_/S vssd1 vssd1 vccd1 vccd1 _5596_/D sky130_fd_sc_hd__mux2_1
X_5367_ _5367_/CLK _5367_/D vssd1 vssd1 vccd1 vccd1 _5367_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput364 _5928_/X vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_12
Xoutput375 _3724_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput386 _3754_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__clkbuf_2
X_2579_ _2743_/A0 _5636_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5636_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _4018_/Y _4318_/A2 _4322_/B _4013_/A vssd1 vssd1 vccd1 vccd1 _4318_/X sky130_fd_sc_hd__o22a_1
X_5298_ _5298_/CLK _5298_/D vssd1 vssd1 vccd1 vccd1 _5298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput397 _3774_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4249_ _5745_/Q _4249_/B vssd1 vssd1 vccd1 vccd1 _4249_/X sky130_fd_sc_hd__xor2_1
XFILLER_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout591 _5692_/Q vssd1 vssd1 vccd1 vccd1 _3339_/A1 sky130_fd_sc_hd__buf_4
Xfanout580 _5694_/Q vssd1 vssd1 vccd1 vccd1 _3394_/A0 sky130_fd_sc_hd__buf_4
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4544__129 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5186_/CLK sky130_fd_sc_hd__inv_2
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3620_ _4389_/B _3617_/B _3618_/X _4966_/Q vssd1 vssd1 vccd1 vccd1 _3778_/C sky130_fd_sc_hd__a31o_4
X_4895__480 _4901__486/A vssd1 vssd1 vccd1 vccd1 _5616_/CLK sky130_fd_sc_hd__inv_2
X_3551_ _5115_/Q _3596_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5115_/D sky130_fd_sc_hd__mux2_1
X_2502_ _4401_/A _3897_/C vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__nand2_4
X_3482_ _3590_/A1 _5177_/Q _3489_/S vssd1 vssd1 vccd1 vccd1 _5177_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5221_ _5221_/CLK _5221_/D vssd1 vssd1 vccd1 vccd1 _5221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2433_ _5748_/Q vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__clkinv_4
X_5152_ _5152_/CLK _5152_/D vssd1 vssd1 vccd1 vccd1 _5152_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2407 hold2407/A vssd1 vssd1 vccd1 vccd1 hold2407/X sky130_fd_sc_hd__buf_2
Xhold2418 hold2418/A vssd1 vssd1 vccd1 vccd1 hold2418/X sky130_fd_sc_hd__buf_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4103_ _5550_/Q _5549_/Q _5548_/Q _5547_/Q vssd1 vssd1 vccd1 vccd1 _4104_/D sky130_fd_sc_hd__and4_2
Xhold2429 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 hold2429/X sky130_fd_sc_hd__buf_2
X_5083_ _5739_/CLK _5083_/D vssd1 vssd1 vccd1 vccd1 _5083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1728 hold2403/X vssd1 vssd1 vccd1 vccd1 hold2404/A sky130_fd_sc_hd__buf_2
X_4034_ _4034_/A _4063_/A _4008_/B vssd1 vssd1 vccd1 vccd1 _4046_/B sky130_fd_sc_hd__or3b_2
XFILLER_65_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_21 _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 hold236/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _5291_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _4352_/A _5017_/Q hold80/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__mux2_1
XANTENNA_65 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 hold980/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3749_ _5086_/Q input15/X _3763_/B vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5419_ _5419_/CLK _5419_/D vssd1 vssd1 vccd1 vccd1 _5419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4493__78 _4509__94/A vssd1 vssd1 vccd1 vccd1 _5135_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4879__464 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5600_/CLK sky130_fd_sc_hd__inv_2
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_709 vssd1 vssd1 vccd1 vccd1 CaravelHost_709/HI manufacturerID[9] sky130_fd_sc_hd__conb_1
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2982_ _2978_/X _2979_/X _3075_/B1 _2976_/X vssd1 vssd1 vccd1 vccd1 _2982_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
X_3603_ _4978_/Q _3603_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4978_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput63 probe_out[34] vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__clkbuf_2
Xinput52 probe_out[24] vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__clkbuf_2
Xinput41 probe_out[14] vssd1 vssd1 vccd1 vccd1 _5851_/A sky130_fd_sc_hd__clkbuf_2
Xhold803 hold803/A vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__buf_2
X_3534_ _5130_/Q _3615_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5130_/D sky130_fd_sc_hd__mux2_1
Xinput96 probe_out[64] vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput85 probe_out[54] vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__clkbuf_2
Xinput74 probe_out[44] vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__clkbuf_2
Xhold825 hold825/A vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3465_ _5192_/Q _3609_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5192_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4672__257 _4485__70/A vssd1 vssd1 vccd1 vccd1 _5360_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold858 hold858/A vssd1 vssd1 vccd1 vccd1 hold858/X sky130_fd_sc_hd__buf_2
XFILLER_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5204_ _5384_/CLK _5204_/D vssd1 vssd1 vccd1 vccd1 _5204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2204 hold2204/A vssd1 vssd1 vccd1 vccd1 hold2204/X sky130_fd_sc_hd__buf_2
Xhold2215 hold2821/X vssd1 vssd1 vccd1 vccd1 hold2215/X sky130_fd_sc_hd__buf_2
Xhold2226 hold2812/X vssd1 vssd1 vccd1 vccd1 hold2813/A sky130_fd_sc_hd__buf_2
Xhold2237 hold2237/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__buf_2
X_3396_ _3396_/A0 _5282_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5282_/D sky130_fd_sc_hd__mux2_1
X_4713__298 _5259_/CLK vssd1 vssd1 vccd1 vccd1 _5404_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5135_ _5135_/CLK _5135_/D vssd1 vssd1 vccd1 vccd1 _5135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1514 hold2292/X vssd1 vssd1 vccd1 vccd1 hold2293/A sky130_fd_sc_hd__buf_2
Xhold1525 hold2326/X vssd1 vssd1 vccd1 vccd1 hold2327/A sky130_fd_sc_hd__buf_2
Xhold2259 hold2259/A vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__buf_2
Xhold1503 hold2272/X vssd1 vssd1 vccd1 vccd1 hold2273/A sky130_fd_sc_hd__buf_2
Xhold2248 hold2248/A vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__buf_2
Xhold1558 hold17/X vssd1 vssd1 vccd1 vccd1 hold1558/X sky130_fd_sc_hd__buf_2
Xhold1547 hold990/X vssd1 vssd1 vccd1 vccd1 _5097_/D sky130_fd_sc_hd__buf_2
X_5066_ _5733_/CLK _5066_/D vssd1 vssd1 vccd1 vccd1 _5066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1536 hold2386/X vssd1 vssd1 vccd1 vccd1 hold2387/A sky130_fd_sc_hd__buf_2
Xhold1569 hold1569/A vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__buf_2
X_4017_ _5678_/Q _4032_/B _5679_/Q vssd1 vssd1 vccd1 vccd1 _4247_/C sky130_fd_sc_hd__a21o_1
X_4566__151 _4508__93/A vssd1 vssd1 vccd1 vccd1 _5216_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5899_ _5899_/A vssd1 vssd1 vccd1 vccd1 _5899_/X sky130_fd_sc_hd__clkbuf_4
X_4607__192 _4463__48/A vssd1 vssd1 vccd1 vccd1 _5281_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2760 _4384_/X vssd1 vssd1 vccd1 vccd1 hold2760/X sky130_fd_sc_hd__buf_2
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2793 hold2793/A vssd1 vssd1 vccd1 vccd1 hold2793/X sky130_fd_sc_hd__buf_2
XFILLER_113_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _5515_/Q _5284_/Q _3299_/S vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _5628_/Q _5518_/Q _5287_/Q _5470_/Q _3219_/S0 _3330_/S vssd1 vssd1 vccd1 vccd1
+ _3181_/X sky130_fd_sc_hd__mux4_2
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5753_ _5755_/CLK _5753_/D vssd1 vssd1 vccd1 vccd1 _5753_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2965_ _5037_/Q _5534_/Q _3072_/S vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2896_ _2863_/A _5382_/Q _3094_/A _2893_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _2896_/X
+ sky130_fd_sc_hd__a221o_1
X_5684_ _5684_/CLK _5684_/D vssd1 vssd1 vccd1 vccd1 _5684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_96_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4898__483/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4510__95/A
+ sky130_fd_sc_hd__clkbuf_16
X_3517_ _3589_/A _3526_/B vssd1 vssd1 vccd1 vccd1 _3525_/S sky130_fd_sc_hd__nor2_8
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold666 hold733/X vssd1 vssd1 vccd1 vccd1 hold734/A sky130_fd_sc_hd__buf_2
Xhold688 hold823/X vssd1 vssd1 vccd1 vccd1 hold824/A sky130_fd_sc_hd__buf_2
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3448_ _3611_/A1 _5214_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5214_/D sky130_fd_sc_hd__mux2_1
Xhold2012 hold2666/X vssd1 vssd1 vccd1 vccd1 hold2667/A sky130_fd_sc_hd__buf_2
Xhold2001 hold2001/A vssd1 vssd1 vccd1 vccd1 _4993_/D sky130_fd_sc_hd__buf_2
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2023 hold2658/X vssd1 vssd1 vccd1 vccd1 hold2659/A sky130_fd_sc_hd__buf_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _3406_/A _3397_/A vssd1 vssd1 vccd1 vccd1 _3387_/S sky130_fd_sc_hd__nor2_8
Xhold2034 hold2680/X vssd1 vssd1 vccd1 vccd1 hold2681/A sky130_fd_sc_hd__buf_2
Xhold2045 hold187/X vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__buf_2
X_5118_ _5118_/CLK _5118_/D vssd1 vssd1 vccd1 vccd1 _5118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2067 hold2706/X vssd1 vssd1 vccd1 vccd1 hold2707/A sky130_fd_sc_hd__buf_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2056 hold2694/X vssd1 vssd1 vccd1 vccd1 hold2695/A sky130_fd_sc_hd__buf_2
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1366 hold2118/X vssd1 vssd1 vccd1 vccd1 hold2119/A sky130_fd_sc_hd__buf_2
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1344 hold2683/X vssd1 vssd1 vccd1 vccd1 hold2036/A sky130_fd_sc_hd__buf_2
Xhold2089 hold2089/A vssd1 vssd1 vccd1 vccd1 hold441/A sky130_fd_sc_hd__buf_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1388 hold2147/X vssd1 vssd1 vccd1 vccd1 hold2148/A sky130_fd_sc_hd__buf_2
X_5049_ _5049_/CLK _5049_/D vssd1 vssd1 vccd1 vccd1 _5049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4463__48 _4463__48/A vssd1 vssd1 vccd1 vccd1 _5057_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2590 _4413_/X vssd1 vssd1 vccd1 vccd1 hold2590/X sky130_fd_sc_hd__buf_2
XFILLER_36_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2750_ _3389_/A0 _5480_/Q _2757_/S vssd1 vssd1 vccd1 vccd1 _5480_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2681_ _2850_/A1 _5568_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5568_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4935__520 _4937__522/A vssd1 vssd1 vccd1 vccd1 _5656_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4351_ _4351_/A _4351_/B split4/A _4357_/C vssd1 vssd1 vccd1 vccd1 _4351_/X sky130_fd_sc_hd__and4_1
XFILLER_140_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4282_ _5664_/Q _5663_/Q vssd1 vssd1 vccd1 vccd1 _4282_/Y sky130_fd_sc_hd__nand2_2
Xfanout409 _4182_/X vssd1 vssd1 vccd1 vccd1 _4187_/B1 sky130_fd_sc_hd__buf_4
X_3302_ _3297_/X _3298_/X _3301_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3302_/X sky130_fd_sc_hd__a211o_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3233_ _5658_/Q _5388_/Q _3327_/S vssd1 vssd1 vccd1 vccd1 _3233_/X sky130_fd_sc_hd__mux2_1
X_4419__4 _4419__4/A vssd1 vssd1 vccd1 vccd1 _4970_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3164_ _3326_/C1 _3161_/X _3163_/X vssd1 vssd1 vccd1 vccd1 _3164_/X sky130_fd_sc_hd__a21o_1
X_3095_ _5368_/Q _3099_/A _3094_/Y _4088_/B vssd1 vssd1 vccd1 vccd1 _5368_/D sky130_fd_sc_hd__o211a_1
XFILLER_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4784__369 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5475_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3997_ _5265_/Q _3660_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _5265_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2948_ _2945_/X _2946_/X _2947_/X _3043_/A _3094_/B vssd1 vssd1 vccd1 vccd1 _2948_/X
+ sky130_fd_sc_hd__o221a_2
X_5736_ _5738_/CLK _5736_/D vssd1 vssd1 vccd1 vccd1 _5736_/Q sky130_fd_sc_hd__dfxtp_1
X_5667_ _5731_/CLK _5667_/D vssd1 vssd1 vccd1 vccd1 _5667_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4678__263 _4425__10/A vssd1 vssd1 vccd1 vccd1 _5367_/CLK sky130_fd_sc_hd__inv_2
X_2879_ _5033_/Q _5177_/Q _5241_/Q _5225_/Q _2944_/S0 _3040_/S vssd1 vssd1 vccd1 vccd1
+ _2879_/X sky130_fd_sc_hd__mux4_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5598_ _5598_/CLK _5598_/D vssd1 vssd1 vccd1 vccd1 _5598_/Q sky130_fd_sc_hd__dfxtp_1
X_4508__93 _4508__93/A vssd1 vssd1 vccd1 vccd1 _5150_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold441 hold441/A vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__buf_2
Xhold463 hold463/A vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__buf_2
Xhold452 hold452/A vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__buf_2
Xhold474 hold474/A vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__buf_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1152 hold2219/X vssd1 vssd1 vccd1 vccd1 hold2220/A sky130_fd_sc_hd__buf_2
XFILLER_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1163 hold1822/X vssd1 vssd1 vccd1 vccd1 hold1823/A sky130_fd_sc_hd__buf_2
Xhold1185 hold2550/X vssd1 vssd1 vccd1 vccd1 hold2551/A sky130_fd_sc_hd__buf_2
XFILLER_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919__504 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5640_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _5737_/Q _3920_/B _5292_/Q vssd1 vssd1 vccd1 vccd1 _3920_/X sky130_fd_sc_hd__and3_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3851_ _5092_/Q _3851_/B _5091_/Q vssd1 vssd1 vccd1 vccd1 _3855_/B sky130_fd_sc_hd__or3b_4
X_2802_ _5437_/Q _3584_/A0 _2806_/S vssd1 vssd1 vccd1 vccd1 _5437_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3782_ _3782_/A _3829_/B vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__or2_4
X_5521_ _5521_/CLK _5521_/D vssd1 vssd1 vccd1 vccd1 _5521_/Q sky130_fd_sc_hd__dfxtp_1
X_2733_ _2790_/A0 _5495_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5495_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5452_ _5452_/CLK _5452_/D vssd1 vssd1 vccd1 vccd1 _5452_/Q sky130_fd_sc_hd__dfxtp_1
X_2664_ _3571_/A _2664_/B vssd1 vssd1 vccd1 vccd1 _2672_/S sky130_fd_sc_hd__nor2_8
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5383_ _5383_/CLK _5383_/D vssd1 vssd1 vccd1 vccd1 _5383_/Q sky130_fd_sc_hd__dfxtp_4
X_4403_ _4356_/A _4357_/B _4415_/A3 _4403_/B1 vssd1 vssd1 vccd1 vccd1 _4403_/X sky130_fd_sc_hd__a31o_1
X_2595_ _5335_/Q _3344_/A _3346_/A vssd1 vssd1 vccd1 vccd1 _2664_/B sky130_fd_sc_hd__nand3_4
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4334_ _5684_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4334_/X sky130_fd_sc_hd__or2_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4265_ _4263_/X _4265_/B _4265_/C _4265_/D vssd1 vssd1 vccd1 vccd1 _4268_/C sky130_fd_sc_hd__and4b_1
X_4196_ _4204_/A _4196_/B vssd1 vssd1 vccd1 vccd1 _5544_/D sky130_fd_sc_hd__nor2_1
X_3216_ _3136_/X _3203_/X _3207_/X _3215_/X vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__a31o_1
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3147_ _5723_/Q _5300_/Q _5273_/Q _5707_/Q _3324_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3147_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4433__18 _4433__18/A vssd1 vssd1 vccd1 vccd1 _5027_/CLK sky130_fd_sc_hd__inv_2
X_3078_ _2863_/A _5375_/Q _3094_/A _3077_/Y _2894_/X vssd1 vssd1 vccd1 vccd1 _3078_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4472__57/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5719_ _5719_/CLK _5719_/D vssd1 vssd1 vccd1 vccd1 _5719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__buf_2
XFILLER_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold282 _3808_/X vssd1 vssd1 vccd1 vccd1 _5008_/D sky130_fd_sc_hd__buf_2
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__buf_2
XFILLER_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4499__84 _4504__89/A vssd1 vssd1 vccd1 vccd1 _5141_/CLK sky130_fd_sc_hd__inv_2
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4050_ _5750_/Q _4254_/B _4254_/C vssd1 vssd1 vccd1 vccd1 _4050_/X sky130_fd_sc_hd__and3_1
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_3001_ _3074_/A1 _2999_/X _3000_/X _3097_/B vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__o211a_1
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3903_ _5075_/Q _3926_/A2 _3925_/B1 _3902_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5075_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3834_ _5557_/Q _3834_/B vssd1 vssd1 vccd1 vccd1 _3834_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3765_ _3765_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__and2_1
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3696_ _4985_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3696_/X sky130_fd_sc_hd__or2_1
X_2716_ _2743_/A0 _5510_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5510_/D sky130_fd_sc_hd__mux2_1
X_5504_ _5504_/CLK _5504_/D vssd1 vssd1 vccd1 vccd1 _5504_/Q sky130_fd_sc_hd__dfxtp_1
X_5435_ _5435_/CLK _5435_/D vssd1 vssd1 vccd1 vccd1 _5435_/Q sky130_fd_sc_hd__dfxtp_1
X_2647_ _5597_/Q _3573_/A0 _2653_/S vssd1 vssd1 vccd1 vccd1 _5597_/D sky130_fd_sc_hd__mux2_1
Xoutput310 _5879_/X vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_12
Xoutput343 _5909_/X vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_12
Xoutput332 _5899_/X vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_12
Xoutput321 _5889_/X vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_12
X_5366_ _5366_/CLK _5366_/D vssd1 vssd1 vccd1 vccd1 _5366_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput365 _5929_/X vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_12
Xoutput354 _5919_/X vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_12
Xoutput387 _3756_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput376 _3727_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__clkbuf_2
X_2578_ _3573_/A0 _5637_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5637_/D sky130_fd_sc_hd__mux2_4
XFILLER_141_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4317_ _4316_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _5678_/D sky130_fd_sc_hd__and2b_1
X_5297_ _5297_/CLK _5297_/D vssd1 vssd1 vccd1 vccd1 _5297_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput398 _3700_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__clkbuf_2
X_4248_ _5744_/Q _4248_/B vssd1 vssd1 vccd1 vccd1 _4248_/X sky130_fd_sc_hd__xor2_1
XFILLER_59_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4179_ _5530_/Q _5529_/Q _4186_/B _4217_/A vssd1 vssd1 vccd1 vccd1 _4179_/X sky130_fd_sc_hd__a31o_1
XFILLER_55_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4840__425 _5001_/CLK vssd1 vssd1 vccd1 vccd1 _5533_/CLK sky130_fd_sc_hd__inv_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout592 _2897_/A1 vssd1 vssd1 vccd1 vccd1 _3590_/A1 sky130_fd_sc_hd__buf_4
XFILLER_76_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout581 _3277_/A1 vssd1 vssd1 vccd1 vccd1 _3577_/A0 sky130_fd_sc_hd__buf_4
Xfanout570 _3409_/A1 vssd1 vssd1 vccd1 vccd1 _3574_/A0 sky130_fd_sc_hd__buf_8
XFILLER_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4583__168 _4509__94/A vssd1 vssd1 vccd1 vccd1 _5233_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _5116_/Q _3595_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5116_/D sky130_fd_sc_hd__mux2_1
X_2501_ _3920_/B _3955_/A vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__or2_2
X_5220_ _5220_/CLK _5220_/D vssd1 vssd1 vccd1 vccd1 _5220_/Q sky130_fd_sc_hd__dfxtp_1
X_3481_ _3607_/A _3589_/B vssd1 vssd1 vccd1 vccd1 _3489_/S sky130_fd_sc_hd__or2_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5151_ _5151_/CLK _5151_/D vssd1 vssd1 vccd1 vccd1 _5151_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2408 hold2408/A vssd1 vssd1 vccd1 vccd1 _5751_/D sky130_fd_sc_hd__buf_2
Xhold2419 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 hold2419/X sky130_fd_sc_hd__buf_2
XFILLER_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5082_ _5739_/CLK _5082_/D vssd1 vssd1 vccd1 vccd1 _5082_/Q sky130_fd_sc_hd__dfxtp_1
X_4102_ _5548_/Q _5547_/Q vssd1 vssd1 vccd1 vccd1 _4108_/D sky130_fd_sc_hd__and2_2
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4033_ _5742_/Q _4270_/B _4031_/X _4028_/X vssd1 vssd1 vccd1 vccd1 _4075_/B sky130_fd_sc_hd__o211ai_4
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1729 hold2405/X vssd1 vssd1 vccd1 vccd1 hold2406/A sky130_fd_sc_hd__buf_2
Xhold1718 hold2378/X vssd1 vssd1 vccd1 vccd1 hold2379/A sky130_fd_sc_hd__buf_2
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824__409 _4909__494/A vssd1 vssd1 vccd1 vccd1 _5515_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_22 _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_66 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _4351_/B _5016_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _5016_/D sky130_fd_sc_hd__mux2_1
XANTENNA_55 hold956/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 hold2295/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3748_ _3824_/A1 _3746_/X _3747_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3748_/X sky130_fd_sc_hd__o211a_4
XANTENNA_77 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4718__303 _4731__316/A vssd1 vssd1 vccd1 vccd1 _5409_/CLK sky130_fd_sc_hd__inv_2
X_3679_ _5252_/Q _3682_/B vssd1 vssd1 vccd1 vccd1 _3679_/X sky130_fd_sc_hd__and2_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5418_ _5418_/CLK _5418_/D vssd1 vssd1 vccd1 vccd1 _5418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5349_ _5349_/CLK _5349_/D vssd1 vssd1 vccd1 vccd1 _5349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4469__54 _4469__54/A vssd1 vssd1 vccd1 vccd1 _5063_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2981_ _3043_/A _2981_/B _2981_/C vssd1 vssd1 vccd1 vccd1 _2981_/X sky130_fd_sc_hd__or3_1
XFILLER_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_2
X_3602_ _4979_/Q _3602_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4979_/D sky130_fd_sc_hd__mux2_1
Xinput64 probe_out[35] vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__clkbuf_2
Xinput53 probe_out[25] vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__clkbuf_2
Xinput42 probe_out[15] vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3533_ _5131_/Q _3614_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5131_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput97 probe_out[65] vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__clkbuf_2
Xinput86 probe_out[55] vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__clkbuf_2
Xinput75 probe_out[45] vssd1 vssd1 vccd1 vccd1 _5882_/A sky130_fd_sc_hd__clkbuf_2
Xhold804 hold804/A vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__buf_2
Xhold826 hold826/A vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__buf_2
X_3464_ _5193_/Q _3608_/A1 _3471_/S vssd1 vssd1 vccd1 vccd1 _5193_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold848 hold848/A vssd1 vssd1 vccd1 vccd1 hold848/X sky130_fd_sc_hd__buf_2
XFILLER_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5203_ _5730_/CLK _5203_/D vssd1 vssd1 vccd1 vccd1 _5203_/Q sky130_fd_sc_hd__dfxtp_1
X_5134_ _5134_/CLK _5134_/D vssd1 vssd1 vccd1 vccd1 _5134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2205 hold2205/A vssd1 vssd1 vccd1 vccd1 hold696/A sky130_fd_sc_hd__buf_2
Xhold2216 hold2216/A vssd1 vssd1 vccd1 vccd1 hold2216/X sky130_fd_sc_hd__buf_2
Xhold2227 hold2814/X vssd1 vssd1 vccd1 vccd1 hold2227/X sky130_fd_sc_hd__buf_2
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3395_ _3395_/A0 _5283_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5283_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1515 hold2294/X vssd1 vssd1 vccd1 vccd1 hold2295/A sky130_fd_sc_hd__buf_2
Xhold2249 hold18/X vssd1 vssd1 vccd1 vccd1 hold2249/X sky130_fd_sc_hd__buf_2
Xhold2238 hold12/X vssd1 vssd1 vccd1 vccd1 hold2238/X sky130_fd_sc_hd__buf_2
Xhold1526 hold2328/X vssd1 vssd1 vccd1 vccd1 hold2329/A sky130_fd_sc_hd__buf_2
Xhold1504 hold2274/X vssd1 vssd1 vccd1 vccd1 hold2275/A sky130_fd_sc_hd__buf_2
X_5065_ _5065_/CLK _5065_/D vssd1 vssd1 vccd1 vccd1 _5065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1559 hold1559/A vssd1 vssd1 vccd1 vccd1 _5098_/D sky130_fd_sc_hd__buf_2
Xhold1548 hold2419/X vssd1 vssd1 vccd1 vccd1 hold2420/A sky130_fd_sc_hd__buf_2
Xhold1537 hold2388/X vssd1 vssd1 vccd1 vccd1 hold2389/A sky130_fd_sc_hd__buf_2
XFILLER_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4016_ _5740_/Q _4016_/B vssd1 vssd1 vccd1 vccd1 _4074_/D sky130_fd_sc_hd__xor2_2
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5898_ _5898_/A vssd1 vssd1 vccd1 vccd1 _5898_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4952__537 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5710_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2772 _4382_/X vssd1 vssd1 vccd1 vccd1 hold2772/X sky130_fd_sc_hd__buf_2
X_4846__431 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5567_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2794 hold2794/A vssd1 vssd1 vccd1 vccd1 _5693_/D sky130_fd_sc_hd__buf_2
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3180_ _3573_/A0 _3159_/B _3179_/X _3277_/C1 vssd1 vssd1 vccd1 vccd1 _5343_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4589__174 _5111_/CLK vssd1 vssd1 vccd1 vccd1 _5239_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2964_ _3034_/A _2962_/X _2963_/X vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__o21a_1
X_5752_ _5752_/CLK _5752_/D vssd1 vssd1 vccd1 vccd1 _5752_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2895_ _5383_/Q _3962_/B vssd1 vssd1 vccd1 vccd1 _2895_/Y sky130_fd_sc_hd__nand2_4
X_5683_ _5683_/CLK _5683_/D vssd1 vssd1 vccd1 vccd1 _5683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3516_ _3615_/A1 _5146_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5146_/D sky130_fd_sc_hd__mux2_1
Xhold667 hold702/X vssd1 vssd1 vccd1 vccd1 hold703/A sky130_fd_sc_hd__buf_2
X_3447_ _3592_/A1 _5215_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5215_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_65_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5262_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold689 hold825/X vssd1 vssd1 vccd1 vccd1 hold826/A sky130_fd_sc_hd__buf_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2024 hold2024/A vssd1 vssd1 vccd1 vccd1 _5345_/D sky130_fd_sc_hd__buf_2
X_3378_ _3579_/A0 _5301_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5301_/D sky130_fd_sc_hd__mux2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2013 hold2013/A vssd1 vssd1 vccd1 vccd1 _4994_/D sky130_fd_sc_hd__buf_2
Xhold2035 hold2682/X vssd1 vssd1 vccd1 vccd1 hold2683/A sky130_fd_sc_hd__buf_2
X_5117_ _5117_/CLK _5117_/D vssd1 vssd1 vccd1 vccd1 _5117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1323 hold2618/X vssd1 vssd1 vccd1 vccd1 hold2619/A sky130_fd_sc_hd__buf_2
Xhold2068 hold2708/X vssd1 vssd1 vccd1 vccd1 hold2709/A sky130_fd_sc_hd__buf_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2057 hold2696/X vssd1 vssd1 vccd1 vccd1 hold2697/A sky130_fd_sc_hd__buf_2
Xhold2046 hold293/X vssd1 vssd1 vccd1 vccd1 hold178/A sky130_fd_sc_hd__buf_2
Xhold1367 hold2120/X vssd1 vssd1 vccd1 vccd1 hold2121/A sky130_fd_sc_hd__buf_2
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1356 hold2687/X vssd1 vssd1 vccd1 vccd1 hold2688/A sky130_fd_sc_hd__buf_2
X_5048_ _5048_/CLK _5048_/D vssd1 vssd1 vccd1 vccd1 _5048_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1389 hold542/X vssd1 vssd1 vccd1 vccd1 _5071_/D sky130_fd_sc_hd__buf_2
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4439__24 _4439__24/A vssd1 vssd1 vccd1 vccd1 _5033_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2591 hold2591/A vssd1 vssd1 vccd1 vccd1 hold2591/X sky130_fd_sc_hd__buf_2
XFILLER_91_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4623__208 _4965__550/A vssd1 vssd1 vccd1 vccd1 _5300_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2680_ _2849_/A1 _5569_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5569_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ _4350_/A split5/X _4357_/C vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__and3_1
XFILLER_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4517__102 _4485__70/A vssd1 vssd1 vccd1 vccd1 _5159_/CLK sky130_fd_sc_hd__inv_2
X_3301_ _3301_/A1 _3299_/X _3300_/X _3171_/A vssd1 vssd1 vccd1 vccd1 _3301_/X sky130_fd_sc_hd__o211a_1
X_4281_ _4281_/A input1/X vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__or2_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3232_ _5719_/Q _3326_/B2 _3323_/C1 _3231_/X vssd1 vssd1 vccd1 vccd1 _3242_/C sky130_fd_sc_hd__o211a_1
X_3163_ _3320_/C1 _3162_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3163_/X sky130_fd_sc_hd__a21o_1
X_3094_ _3094_/A _3094_/B vssd1 vssd1 vccd1 vccd1 _3094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_112_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5247_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3996_ _5264_/Q _3659_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _5264_/D sky130_fd_sc_hd__mux2_1
X_2947_ _2937_/X _2938_/X _2947_/S vssd1 vssd1 vccd1 vccd1 _2947_/X sky130_fd_sc_hd__mux2_1
X_5735_ _5735_/CLK _5735_/D vssd1 vssd1 vccd1 vccd1 _5735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5666_ _5731_/CLK _5666_/D vssd1 vssd1 vccd1 vccd1 _5666_/Q sky130_fd_sc_hd__dfxtp_4
X_2878_ _5201_/Q _5185_/Q _4974_/Q _5193_/Q _3036_/S _2943_/S1 vssd1 vssd1 vccd1 vccd1
+ _2878_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5597_ _5597_/CLK _5597_/D vssd1 vssd1 vccd1 vccd1 _5597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold431 hold500/X vssd1 vssd1 vccd1 vccd1 hold501/A sky130_fd_sc_hd__buf_2
XFILLER_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold453 hold453/A vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__buf_2
XFILLER_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1120 hold1120/A vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__buf_2
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 hold1824/X vssd1 vssd1 vccd1 vccd1 hold1825/A sky130_fd_sc_hd__buf_2
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1197 hold1904/X vssd1 vssd1 vccd1 vccd1 hold1905/A sky130_fd_sc_hd__buf_2
Xhold1186 hold2554/X vssd1 vssd1 vccd1 vccd1 hold2555/A sky130_fd_sc_hd__buf_2
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958__543 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5716_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _4399_/C _3850_/B _3850_/C _3850_/D vssd1 vssd1 vccd1 vccd1 _3857_/B sky130_fd_sc_hd__or4_4
X_2801_ _5438_/Q _3601_/A1 _2806_/S vssd1 vssd1 vccd1 vccd1 _5438_/D sky130_fd_sc_hd__mux2_1
X_3781_ _3782_/A _3829_/B vssd1 vssd1 vccd1 vccd1 _3781_/Y sky130_fd_sc_hd__nor2_8
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2732_ _3159_/A _5496_/Q _2739_/S vssd1 vssd1 vccd1 vccd1 _5496_/D sky130_fd_sc_hd__mux2_1
X_5520_ _5520_/CLK _5520_/D vssd1 vssd1 vccd1 vccd1 _5520_/Q sky130_fd_sc_hd__dfxtp_1
X_4421__6 _4421__6/A vssd1 vssd1 vccd1 vccd1 _4972_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2663_ _3606_/A1 _5583_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5583_/D sky130_fd_sc_hd__mux2_1
X_5451_ _5451_/CLK _5451_/D vssd1 vssd1 vccd1 vccd1 _5451_/Q sky130_fd_sc_hd__dfxtp_1
X_5382_ _5382_/CLK _5382_/D vssd1 vssd1 vccd1 vccd1 _5382_/Q sky130_fd_sc_hd__dfxtp_1
X_4402_ _5748_/Q _4415_/A3 hold691/X hold711/A vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__o211a_1
X_2594_ _3396_/A0 _5623_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5623_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4333_ _4325_/Y _4331_/X _4332_/X vssd1 vssd1 vccd1 vccd1 _5683_/D sky130_fd_sc_hd__a21oi_1
X_4751__336 _5024_/CLK vssd1 vssd1 vccd1 vccd1 _5442_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4264_ _5747_/Q _4264_/B vssd1 vssd1 vccd1 vccd1 _4265_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3215_ _3334_/A1 _3210_/X _3213_/X _3214_/X _3169_/B vssd1 vssd1 vccd1 vccd1 _3215_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4195_ _5544_/Q _4187_/B1 _4210_/C _4130_/Y vssd1 vssd1 vccd1 vccd1 _4196_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3146_ _5057_/Q _5281_/Q _5528_/Q _5308_/Q _3324_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3146_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3077_ _3077_/A _3077_/B vssd1 vssd1 vccd1 vccd1 _3077_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4645__230 _5553_/CLK vssd1 vssd1 vccd1 vccd1 _5331_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3979_ _3644_/A _5249_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _5249_/D sky130_fd_sc_hd__mux2_1
X_5718_ _5718_/CLK _5718_/D vssd1 vssd1 vccd1 vccd1 _5718_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_80_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4965__550/A sky130_fd_sc_hd__clkbuf_16
X_5649_ _5649_/CLK _5649_/D vssd1 vssd1 vccd1 vccd1 _5649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold250 _3805_/X vssd1 vssd1 vccd1 vccd1 _5005_/D sky130_fd_sc_hd__buf_2
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XCaravelHost_690 vssd1 vssd1 vccd1 vccd1 CaravelHost_690/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__buf_2
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__buf_2
XFILLER_104_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
X_3000_ _5435_/Q _2460_/Y _3031_/B1 _5427_/Q vssd1 vssd1 vccd1 vccd1 _3000_/X sky130_fd_sc_hd__o22a_1
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4629__214 _5683_/CLK vssd1 vssd1 vccd1 vccd1 _5306_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3902_ _5746_/Q _3924_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3902_/X sky130_fd_sc_hd__and3_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3833_ _5558_/Q _5559_/Q _5560_/Q _5561_/Q _5555_/Q _5556_/Q vssd1 vssd1 vccd1 vccd1
+ _3834_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3764_ _5009_/Q _3774_/A2 _3774_/B1 _3763_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3764_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3695_ _5068_/Q input25/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__mux2_1
X_2715_ _2790_/A0 _5511_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5511_/D sky130_fd_sc_hd__mux2_1
X_5503_ _5503_/CLK _5503_/D vssd1 vssd1 vccd1 vccd1 _5503_/Q sky130_fd_sc_hd__dfxtp_1
X_5434_ _5434_/CLK _5434_/D vssd1 vssd1 vccd1 vccd1 _5434_/Q sky130_fd_sc_hd__dfxtp_1
X_2646_ _5598_/Q _3159_/A _2653_/S vssd1 vssd1 vccd1 vccd1 _5598_/D sky130_fd_sc_hd__mux2_1
Xoutput300 _5870_/X vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_12
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput344 _5910_/X vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_12
Xoutput322 _5890_/X vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_12
Xoutput333 _5900_/X vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_12
Xoutput311 _5880_/X vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_12
XFILLER_102_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5365_ _5365_/CLK _5365_/D vssd1 vssd1 vccd1 vccd1 _5365_/Q sky130_fd_sc_hd__dfxtp_4
Xoutput366 _5930_/X vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_12
Xoutput355 _5920_/X vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_12
Xoutput377 _3730_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__clkbuf_2
X_2577_ _3159_/A _5638_/Q _2584_/S vssd1 vssd1 vccd1 vccd1 _5638_/D sky130_fd_sc_hd__mux2_4
X_4316_ _4270_/B _4318_/A2 _4322_/B _4013_/B vssd1 vssd1 vccd1 vccd1 _4316_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput399 _3703_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput388 _3758_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__clkbuf_2
X_5296_ _5296_/CLK _5296_/D vssd1 vssd1 vccd1 vccd1 _5296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4247_ _5740_/Q _4247_/B _4247_/C vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__and3_1
XFILLER_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4178_ _4244_/S _4178_/B _4178_/C vssd1 vssd1 vccd1 vccd1 _5529_/D sky130_fd_sc_hd__and3_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3129_ _3130_/B _3281_/S _2464_/A vssd1 vssd1 vccd1 vccd1 _3132_/A sky130_fd_sc_hd__a21oi_4
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout560 _2853_/A1 vssd1 vssd1 vccd1 vccd1 _3389_/A0 sky130_fd_sc_hd__buf_4
Xfanout593 _2897_/A1 vssd1 vssd1 vccd1 vccd1 _3608_/A1 sky130_fd_sc_hd__buf_2
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout582 _3277_/A1 vssd1 vssd1 vccd1 vccd1 _3568_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout571 _5697_/Q vssd1 vssd1 vccd1 vccd1 _3409_/A1 sky130_fd_sc_hd__buf_6
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3480_ _3615_/A1 _5178_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5178_/D sky130_fd_sc_hd__mux2_1
X_2500_ _3920_/B _3955_/A vssd1 vssd1 vccd1 vccd1 _3930_/C sky130_fd_sc_hd__nor2_2
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5150_ _5150_/CLK _5150_/D vssd1 vssd1 vccd1 vccd1 _5150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2409 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 hold2409/X sky130_fd_sc_hd__buf_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5081_ _5677_/CLK _5081_/D vssd1 vssd1 vccd1 vccd1 _5081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4101_ _4132_/B _4119_/C vssd1 vssd1 vccd1 vccd1 _4167_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _5678_/Q _4032_/B vssd1 vssd1 vccd1 vccd1 _4270_/B sky130_fd_sc_hd__xnor2_4
Xhold1719 hold2380/X vssd1 vssd1 vccd1 vccd1 hold2381/A sky130_fd_sc_hd__buf_2
XFILLER_2_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4863__448 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5584_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5111_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4904__489 _4937__522/A vssd1 vssd1 vccd1 vccd1 _5625_/CLK sky130_fd_sc_hd__inv_2
XANTENNA_23 _3637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_12 wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 hold973/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ _4350_/A _5015_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _5015_/D sky130_fd_sc_hd__mux2_1
XANTENNA_34 hold2430/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_67 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3747_ _5002_/Q _3750_/B vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__or2_1
XANTENNA_78 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4757__342 _5697_/CLK vssd1 vssd1 vccd1 vccd1 _5448_/CLK sky130_fd_sc_hd__inv_2
X_3678_ _5251_/Q _3682_/B vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__and2_1
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2629_ _2776_/A _3066_/S _2617_/X vssd1 vssd1 vccd1 vccd1 _2862_/C sky130_fd_sc_hd__a21oi_1
X_5417_ _5417_/CLK _5417_/D vssd1 vssd1 vccd1 vccd1 _5417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5348_ _5348_/CLK _5348_/D vssd1 vssd1 vccd1 vccd1 _5348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5279_ _5279_/CLK _5279_/D vssd1 vssd1 vccd1 vccd1 _5279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550__135 _4422__7/A vssd1 vssd1 vccd1 vccd1 _5192_/CLK sky130_fd_sc_hd__inv_2
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4484__69 _5007_/CLK vssd1 vssd1 vccd1 vccd1 _5126_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ _2971_/X _2973_/X _2919_/B _2970_/X vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__a211o_1
XFILLER_61_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__clkbuf_2
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
X_3601_ _4980_/Q _3601_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4980_/D sky130_fd_sc_hd__mux2_1
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_2
Xinput54 probe_out[26] vssd1 vssd1 vccd1 vccd1 _5863_/A sky130_fd_sc_hd__clkbuf_2
Xinput43 probe_out[16] vssd1 vssd1 vccd1 vccd1 _5853_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3532_ _5132_/Q _3613_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5132_/D sky130_fd_sc_hd__mux2_1
Xinput98 probe_out[66] vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput87 probe_out[56] vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__clkbuf_2
Xinput76 probe_out[46] vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__clkbuf_2
Xinput65 probe_out[36] vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__clkbuf_2
Xhold816 hold816/A vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__buf_2
Xhold827 _4396_/X vssd1 vssd1 vccd1 vccd1 _5746_/D sky130_fd_sc_hd__buf_2
X_3463_ _3526_/A _3607_/B vssd1 vssd1 vccd1 vccd1 _3471_/S sky130_fd_sc_hd__nor2_8
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5202_ _5730_/CLK _5202_/D vssd1 vssd1 vccd1 vccd1 _5202_/Q sky130_fd_sc_hd__dfxtp_1
X_5133_ _5133_/CLK _5133_/D vssd1 vssd1 vccd1 vccd1 _5133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2206 hold696/X vssd1 vssd1 vccd1 vccd1 hold2206/X sky130_fd_sc_hd__buf_2
Xhold2228 hold2228/A vssd1 vssd1 vccd1 vccd1 hold2228/X sky130_fd_sc_hd__buf_2
Xhold2217 hold2217/A vssd1 vssd1 vccd1 vccd1 hold628/A sky130_fd_sc_hd__buf_2
X_3394_ _3394_/A0 _5284_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5284_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1516 hold2296/X vssd1 vssd1 vccd1 vccd1 hold2297/A sky130_fd_sc_hd__buf_2
Xhold2239 hold2239/A vssd1 vssd1 vccd1 vccd1 hold956/A sky130_fd_sc_hd__buf_2
Xhold1505 hold975/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__buf_2
X_5064_ _5064_/CLK _5064_/D vssd1 vssd1 vccd1 vccd1 _5064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1549 hold2421/X vssd1 vssd1 vccd1 vccd1 hold2422/A sky130_fd_sc_hd__buf_2
Xhold1527 hold2330/X vssd1 vssd1 vccd1 vccd1 hold2331/A sky130_fd_sc_hd__buf_2
Xhold1538 hold2390/X vssd1 vssd1 vccd1 vccd1 hold2391/A sky130_fd_sc_hd__buf_2
X_4015_ _5680_/Q _4247_/B _4014_/X vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__a21oi_4
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5897_ _5897_/A vssd1 vssd1 vccd1 vccd1 _5897_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_40_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4534__119 _4438__23/A vssd1 vssd1 vccd1 vccd1 _5176_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2740 hold2740/A vssd1 vssd1 vccd1 vccd1 hold2740/X sky130_fd_sc_hd__buf_2
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4885__470 _5252_/CLK vssd1 vssd1 vccd1 vccd1 _5606_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2963_ _5602_/Q _2460_/A _3073_/B2 _5586_/Q _3073_/C1 vssd1 vssd1 vccd1 vccd1 _2963_/X
+ sky130_fd_sc_hd__o221a_1
X_5751_ _5751_/CLK _5751_/D vssd1 vssd1 vccd1 vccd1 _5751_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2894_ _5383_/Q _3962_/B vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__and2_4
X_5682_ _5691_/CLK _5682_/D vssd1 vssd1 vccd1 vccd1 _5682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3515_ _3596_/A1 _5147_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5147_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold668 _4190_/Y vssd1 vssd1 vccd1 vccd1 _5541_/D sky130_fd_sc_hd__buf_2
X_3446_ _3591_/A1 _5216_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5216_/D sky130_fd_sc_hd__mux2_1
X_4869__454 _5106_/CLK vssd1 vssd1 vccd1 vccd1 _5590_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _3569_/A1 _5302_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5302_/D sky130_fd_sc_hd__mux2_1
Xhold2036 hold2036/A vssd1 vssd1 vccd1 vccd1 _4992_/D sky130_fd_sc_hd__buf_2
X_5116_ _5116_/CLK _5116_/D vssd1 vssd1 vccd1 vccd1 _5116_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2047 _3956_/X vssd1 vssd1 vccd1 vccd1 hold2047/X sky130_fd_sc_hd__buf_2
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 hold929/X vssd1 vssd1 vccd1 vccd1 hold2069/X sky130_fd_sc_hd__buf_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 hold2622/X vssd1 vssd1 vccd1 vccd1 hold1989/A sky130_fd_sc_hd__buf_2
Xhold2058 hold2698/X vssd1 vssd1 vccd1 vccd1 hold2058/X sky130_fd_sc_hd__buf_2
XFILLER_85_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1368 hold489/X vssd1 vssd1 vccd1 vccd1 _5068_/D sky130_fd_sc_hd__buf_2
Xhold1357 hold2691/X vssd1 vssd1 vccd1 vccd1 hold2042/A sky130_fd_sc_hd__buf_2
Xhold1335 hold2663/X vssd1 vssd1 vccd1 vccd1 hold2664/A sky130_fd_sc_hd__buf_2
X_5047_ _5047_/CLK _5047_/D vssd1 vssd1 vccd1 vccd1 _5047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4504__89/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1379 hold2134/X vssd1 vssd1 vccd1 vccd1 hold2135/A sky130_fd_sc_hd__buf_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput200 hold89/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__buf_8
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2592 hold2592/A vssd1 vssd1 vccd1 vccd1 hold2592/X sky130_fd_sc_hd__buf_2
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4454__39 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5048_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4662__247 _4435__20/A vssd1 vssd1 vccd1 vccd1 _5350_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4703__288 _5106_/CLK vssd1 vssd1 vccd1 vccd1 _5394_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4556__141 _4418__3/A vssd1 vssd1 vccd1 vccd1 _5198_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3300_ _5474_/Q _3331_/A2 _3237_/B _5709_/Q vssd1 vssd1 vccd1 vccd1 _3300_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4280_ _4281_/A input1/X vssd1 vssd1 vccd1 vccd1 _4283_/C sky130_fd_sc_hd__nor2_1
XFILLER_100_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3231_ _5703_/Q _3132_/A _3230_/X _3325_/A vssd1 vssd1 vccd1 vccd1 _3231_/X sky130_fd_sc_hd__o22a_1
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3162_ _5722_/Q _5299_/Q _5272_/Q _5706_/Q _3324_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3162_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _3093_/A _3093_/B vssd1 vssd1 vccd1 vccd1 _5369_/D sky130_fd_sc_hd__nor2_1
XFILLER_82_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3995_ _5263_/Q _3658_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _5263_/D sky130_fd_sc_hd__mux2_1
X_2946_ _2947_/S _2943_/X _2919_/B vssd1 vssd1 vccd1 vccd1 _2946_/X sky130_fd_sc_hd__a21o_1
X_5734_ _5734_/CLK _5734_/D vssd1 vssd1 vccd1 vccd1 _5734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2877_ _2871_/X _2876_/X _2945_/A vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__mux2_1
X_5665_ _5731_/CLK _5665_/D vssd1 vssd1 vccd1 vccd1 _5665_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5596_ _5596_/CLK _5596_/D vssd1 vssd1 vccd1 vccd1 _5596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold432 hold504/X vssd1 vssd1 vccd1 vccd1 hold505/A sky130_fd_sc_hd__buf_2
Xhold454 _3785_/X vssd1 vssd1 vccd1 vccd1 _4985_/D sky130_fd_sc_hd__buf_2
XFILLER_131_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3429_ _5230_/Q _3593_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5230_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 hold198/X vssd1 vssd1 vccd1 vccd1 hold1121/X sky130_fd_sc_hd__buf_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1132 hold2379/X vssd1 vssd1 vccd1 vccd1 hold2380/A sky130_fd_sc_hd__buf_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1176 hold1871/X vssd1 vssd1 vccd1 vccd1 hold1872/A sky130_fd_sc_hd__buf_2
XFILLER_85_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1165 hold1826/X vssd1 vssd1 vccd1 vccd1 hold1827/A sky130_fd_sc_hd__buf_2
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1198 hold1906/X vssd1 vssd1 vccd1 vccd1 hold1907/A sky130_fd_sc_hd__buf_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2800_ _5439_/Q _3501_/A1 _2806_/S vssd1 vssd1 vccd1 vccd1 _5439_/D sky130_fd_sc_hd__mux2_1
X_3780_ _5024_/Q _5023_/Q vssd1 vssd1 vccd1 vccd1 _3829_/B sky130_fd_sc_hd__nand2b_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2731_ _3397_/A _2740_/B vssd1 vssd1 vccd1 vccd1 _2739_/S sky130_fd_sc_hd__or2_4
X_5450_ _5450_/CLK _5450_/D vssd1 vssd1 vccd1 vccd1 _5450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2662_ _3605_/A1 _5584_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5584_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4401_ _4401_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _4401_/Y sky130_fd_sc_hd__nand2_2
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5381_ _5381_/CLK _5381_/D vssd1 vssd1 vccd1 vccd1 _5381_/Q sky130_fd_sc_hd__dfxtp_1
X_2593_ _3395_/A0 _5624_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5624_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4332_ _4080_/A _4325_/B _4082_/A vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__a21bo_1
X_4790__375 _4897__482/A vssd1 vssd1 vccd1 vccd1 _5481_/CLK sky130_fd_sc_hd__inv_2
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4263_ _5746_/Q _4039_/X _4260_/X _4261_/Y _4262_/Y vssd1 vssd1 vccd1 vccd1 _4263_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3214_ _3282_/C1 _3211_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3214_/X sky130_fd_sc_hd__a21o_1
X_4194_ _4204_/A _4194_/B vssd1 vssd1 vccd1 vccd1 _5543_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145_ _3171_/A _3145_/B vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__and2_1
X_3076_ _3094_/B _3065_/Y _3068_/Y _3075_/X vssd1 vssd1 vccd1 vccd1 _3077_/B sky130_fd_sc_hd__a31o_1
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3978_ _3643_/A _5248_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _3978_/X sky130_fd_sc_hd__mux2_1
X_2929_ _2924_/X _2927_/X _2928_/X _3043_/A _3094_/B vssd1 vssd1 vccd1 vccd1 _2929_/X
+ sky130_fd_sc_hd__o221a_2
X_5717_ _5717_/CLK _5717_/D vssd1 vssd1 vccd1 vccd1 _5717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _5648_/CLK _5648_/D vssd1 vssd1 vccd1 vccd1 _5648_/Q sky130_fd_sc_hd__dfxtp_1
X_5579_ _5579_/CLK _5579_/D vssd1 vssd1 vccd1 vccd1 _5579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XCaravelHost_691 vssd1 vssd1 vccd1 vccd1 CaravelHost_691/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XCaravelHost_680 vssd1 vssd1 vccd1 vccd1 CaravelHost_680/HI la_data_out[108] sky130_fd_sc_hd__conb_1
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__buf_2
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__buf_2
XFILLER_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__buf_2
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold284 hold351/X vssd1 vssd1 vccd1 vccd1 hold352/A sky130_fd_sc_hd__buf_2
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__buf_2
XFILLER_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4925__510 _4455__40/A vssd1 vssd1 vccd1 vccd1 _5646_/CLK sky130_fd_sc_hd__inv_2
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774__359 _5243_/CLK vssd1 vssd1 vccd1 vccd1 _5465_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
X_4668__253 _5004_/CLK vssd1 vssd1 vccd1 vccd1 _5356_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4709__294 _5010_/CLK vssd1 vssd1 vccd1 vccd1 _5400_/CLK sky130_fd_sc_hd__inv_2
X_3901_ _4369_/A _3855_/X _3887_/X hold554/X vssd1 vssd1 vccd1 vccd1 _3901_/X sky130_fd_sc_hd__a31o_4
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _4351_/B _4357_/B _3832_/A3 _4361_/A vssd1 vssd1 vccd1 vccd1 _3832_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3763_ _3763_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3763_/X sky130_fd_sc_hd__and2_1
X_5502_ _5502_/CLK _5502_/D vssd1 vssd1 vccd1 vccd1 _5502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _3718_/A1 _3692_/X _3693_/X split4/X vssd1 vssd1 vccd1 vccd1 _3694_/X sky130_fd_sc_hd__o211a_1
X_2714_ _3389_/A0 _5512_/Q _2721_/S vssd1 vssd1 vccd1 vccd1 _5512_/D sky130_fd_sc_hd__mux2_1
X_5433_ _5433_/CLK _5433_/D vssd1 vssd1 vccd1 vccd1 _5433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2645_ _3397_/A _2664_/B vssd1 vssd1 vccd1 vccd1 _2653_/S sky130_fd_sc_hd__nor2_8
Xoutput301 _5871_/X vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_12
X_5364_ _5364_/CLK _5364_/D vssd1 vssd1 vccd1 vccd1 _5364_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput334 _5901_/X vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput312 _5881_/X vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_12
Xoutput323 _5891_/X vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_12
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4315_ _4314_/X _4315_/B vssd1 vssd1 vccd1 vccd1 _4315_/X sky130_fd_sc_hd__and2b_1
Xoutput367 _5931_/X vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_12
Xoutput356 _5921_/X vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_12
Xoutput345 _5911_/X vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_12
Xoutput378 _3733_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__clkbuf_2
X_2576_ _3571_/B _3397_/A vssd1 vssd1 vccd1 vccd1 _2584_/S sky130_fd_sc_hd__or2_4
XFILLER_141_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5295_ _5295_/CLK _5295_/D vssd1 vssd1 vccd1 vccd1 _5295_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput389 _3760_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4246_ _4247_/B _4247_/C _5740_/Q vssd1 vssd1 vccd1 vccd1 _4246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4177_ _5529_/Q _4177_/B _4177_/C _4177_/D vssd1 vssd1 vccd1 vccd1 _4177_/X sky130_fd_sc_hd__and4_1
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3128_ _3128_/A _3128_/B vssd1 vssd1 vccd1 vccd1 _3128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3059_ _5599_/Q _2867_/A _2866_/B _5583_/Q _3064_/C1 vssd1 vssd1 vccd1 vccd1 _3059_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout550 _4099_/X vssd1 vssd1 vccd1 vccd1 _4132_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout583 _5694_/Q vssd1 vssd1 vccd1 vccd1 _3277_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout561 _5699_/Q vssd1 vssd1 vccd1 vccd1 _2853_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout572 _5696_/Q vssd1 vssd1 vccd1 vccd1 _3392_/A0 sky130_fd_sc_hd__buf_4
Xfanout594 _2897_/A1 vssd1 vssd1 vccd1 vccd1 _3599_/A1 sky130_fd_sc_hd__buf_4
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5080_ _5742_/CLK _5080_/D vssd1 vssd1 vccd1 vccd1 _5080_/Q sky130_fd_sc_hd__dfxtp_1
X_4100_ _5546_/Q _5545_/Q _5544_/Q _5543_/Q vssd1 vssd1 vccd1 vccd1 _4119_/C sky130_fd_sc_hd__and4_4
Xhold1709 hold2813/X vssd1 vssd1 vccd1 vccd1 hold2814/A sky130_fd_sc_hd__buf_2
X_4031_ _5746_/Q _4249_/B vssd1 vssd1 vccd1 vccd1 _4031_/X sky130_fd_sc_hd__xor2_4
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 _3671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _4746__331/A sky130_fd_sc_hd__clkbuf_16
X_3815_ hold97/A hold76/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__nand2_8
XANTENNA_24 _3770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 hold2249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 hold986/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_68 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3746_ _5085_/Q input13/X _3763_/B vssd1 vssd1 vccd1 vccd1 _3746_/X sky130_fd_sc_hd__mux2_1
X_4796__381 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5487_/CLK sky130_fd_sc_hd__inv_2
XANTENNA_79 _3661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3677_ _5250_/Q _3682_/B vssd1 vssd1 vccd1 vccd1 _3677_/X sky130_fd_sc_hd__and2_1
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5416_ _5416_/CLK _5416_/D vssd1 vssd1 vccd1 vccd1 _5416_/Q sky130_fd_sc_hd__dfxtp_1
X_2628_ _3443_/B _5367_/Q vssd1 vssd1 vccd1 vccd1 _2861_/B sky130_fd_sc_hd__xor2_1
XFILLER_142_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5347_ _5347_/CLK _5347_/D vssd1 vssd1 vccd1 vccd1 _5347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2559_ _3573_/A0 _5653_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5653_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _5278_/CLK _5278_/D vssd1 vssd1 vccd1 vccd1 _5278_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2900 hold2900/A vssd1 vssd1 vccd1 vccd1 _5752_/D sky130_fd_sc_hd__buf_2
X_4229_ _5337_/Q _4360_/B _4164_/B _4228_/X _4244_/S vssd1 vssd1 vccd1 vccd1 _5558_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__clkbuf_2
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3600_ _4981_/Q _3600_/A1 _3606_/S vssd1 vssd1 vccd1 vccd1 _4981_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_2
X_3531_ _5133_/Q _3612_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5133_/D sky130_fd_sc_hd__mux2_1
Xinput55 probe_out[27] vssd1 vssd1 vccd1 vccd1 _5864_/A sky130_fd_sc_hd__clkbuf_2
Xinput44 probe_out[17] vssd1 vssd1 vccd1 vccd1 _5854_/A sky130_fd_sc_hd__clkbuf_2
Xinput88 probe_out[57] vssd1 vssd1 vccd1 vccd1 _5894_/A sky130_fd_sc_hd__clkbuf_2
Xinput77 probe_out[47] vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__clkbuf_2
Xinput66 probe_out[37] vssd1 vssd1 vccd1 vccd1 _5874_/A sky130_fd_sc_hd__clkbuf_2
X_3462_ _3615_/A1 _5194_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5194_/D sky130_fd_sc_hd__mux2_1
Xinput99 probe_out[67] vssd1 vssd1 vccd1 vccd1 _5904_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5201_ _5201_/CLK _5201_/D vssd1 vssd1 vccd1 vccd1 _5201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4830__415 _4460__45/A vssd1 vssd1 vccd1 vccd1 _5521_/CLK sky130_fd_sc_hd__inv_2
X_3393_ _3393_/A0 _5285_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5285_/D sky130_fd_sc_hd__mux2_1
X_5132_ _5132_/CLK _5132_/D vssd1 vssd1 vccd1 vccd1 _5132_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2207 hold2207/A vssd1 vssd1 vccd1 vccd1 hold2207/X sky130_fd_sc_hd__buf_2
Xhold2218 hold628/X vssd1 vssd1 vccd1 vccd1 hold2218/X sky130_fd_sc_hd__buf_2
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2229 hold2229/A vssd1 vssd1 vccd1 vccd1 hold641/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_106_wb_clk_i _5743_/CLK vssd1 vssd1 vccd1 vccd1 _5742_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1517 hold981/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__buf_2
Xhold1506 hold31/X vssd1 vssd1 vccd1 vccd1 hold976/A sky130_fd_sc_hd__buf_2
X_5063_ _5063_/CLK _5063_/D vssd1 vssd1 vccd1 vccd1 _5063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1528 hold2332/X vssd1 vssd1 vccd1 vccd1 hold2333/A sky130_fd_sc_hd__buf_2
Xhold1539 hold2392/X vssd1 vssd1 vccd1 vccd1 hold2393/A sky130_fd_sc_hd__buf_2
XFILLER_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4014_ _5680_/Q _5679_/Q _5678_/Q _4032_/B vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__and4b_2
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5896_ _5896_/A vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3729_ _4996_/Q _3729_/B vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__or2_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4573__158 _5111_/CLK vssd1 vssd1 vccd1 vccd1 _5223_/CLK sky130_fd_sc_hd__inv_2
XFILLER_130_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2730 _4371_/X vssd1 vssd1 vccd1 vccd1 hold2730/X sky130_fd_sc_hd__buf_2
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2752 _4386_/X vssd1 vssd1 vccd1 vccd1 hold2752/X sky130_fd_sc_hd__buf_2
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4614__199 _5022_/CLK vssd1 vssd1 vccd1 vccd1 _5288_/CLK sky130_fd_sc_hd__inv_2
Xhold2796 _4360_/Y vssd1 vssd1 vccd1 vccd1 hold2796/X sky130_fd_sc_hd__buf_2
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5024_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2962_ _5452_/Q _5570_/Q _3024_/S vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5750_ _5751_/CLK _5750_/D vssd1 vssd1 vccd1 vccd1 _5750_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5681_ _5735_/CLK _5681_/D vssd1 vssd1 vccd1 vccd1 _5681_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2893_ _2883_/X _2888_/X _2892_/X _2884_/X vssd1 vssd1 vccd1 vccd1 _2893_/X sky130_fd_sc_hd__a31o_2
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3514_ _3595_/A1 _5148_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5148_/D sky130_fd_sc_hd__mux2_1
X_3445_ _3590_/A1 _5217_/Q _3452_/S vssd1 vssd1 vccd1 vccd1 _5217_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3376_ _3568_/A1 _5303_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5303_/D sky130_fd_sc_hd__mux2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2004 hold2641/X vssd1 vssd1 vccd1 vccd1 hold2642/A sky130_fd_sc_hd__buf_2
X_5115_ _5115_/CLK _5115_/D vssd1 vssd1 vccd1 vccd1 _5115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2048 hold2048/A vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__buf_2
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1303 _4389_/X vssd1 vssd1 vccd1 vccd1 hold458/A sky130_fd_sc_hd__buf_2
XFILLER_58_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 hold2605/X vssd1 vssd1 vccd1 vccd1 hold2606/A sky130_fd_sc_hd__buf_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2059 hold2059/A vssd1 vssd1 vccd1 vccd1 _4996_/D sky130_fd_sc_hd__buf_2
XFILLER_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1336 hold2667/X vssd1 vssd1 vccd1 vccd1 hold2013/A sky130_fd_sc_hd__buf_2
X_5046_ _5046_/CLK _5046_/D vssd1 vssd1 vccd1 vccd1 _5046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_74_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5683_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5879_/A vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput201 hold170/X vssd1 vssd1 vccd1 vccd1 _3626_/A sky130_fd_sc_hd__buf_8
XFILLER_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2582 _3931_/A vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__buf_2
XFILLER_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2593 hold2593/A vssd1 vssd1 vccd1 vccd1 hold205/A sky130_fd_sc_hd__buf_2
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_90_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4595__180 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5269_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3230_ _5269_/Q _5296_/Q _3290_/S vssd1 vssd1 vccd1 vccd1 _3230_/X sky130_fd_sc_hd__mux2_1
X_3161_ _5056_/Q _5280_/Q _5527_/Q _5307_/Q _3324_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3161_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3092_ _5369_/Q _2634_/B _2778_/A vssd1 vssd1 vccd1 vccd1 _3093_/B sky130_fd_sc_hd__o21ai_1
XFILLER_82_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942__527 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5700_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3994_ _5262_/Q _3657_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _5262_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2945_/A _2945_/B vssd1 vssd1 vccd1 vccd1 _2945_/X sky130_fd_sc_hd__and2_1
X_5733_ _5733_/CLK _5733_/D vssd1 vssd1 vccd1 vccd1 _5733_/Q sky130_fd_sc_hd__dfxtp_1
X_2876_ _5121_/Q _5169_/Q _5354_/Q _5233_/Q _2944_/S0 _3040_/S vssd1 vssd1 vccd1 vccd1
+ _2876_/X sky130_fd_sc_hd__mux4_1
X_5664_ _5735_/CLK _5664_/D vssd1 vssd1 vccd1 vccd1 _5664_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4836__421 _4463__48/A vssd1 vssd1 vccd1 vccd1 _5527_/CLK sky130_fd_sc_hd__inv_2
X_5595_ _5595_/CLK _5595_/D vssd1 vssd1 vccd1 vccd1 _5595_/Q sky130_fd_sc_hd__dfxtp_1
Xhold400 hold400/A vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__buf_2
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold433 _4315_/X vssd1 vssd1 vccd1 vccd1 _5677_/D sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_121_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5019_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3428_ _5231_/Q _3592_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5231_/D sky130_fd_sc_hd__mux2_1
Xhold499 hold517/X vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__buf_2
Xhold488 hold488/A vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__buf_2
X_3359_ _3281_/S _3353_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _3359_/Y sky130_fd_sc_hd__o21ai_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 hold2370/X vssd1 vssd1 vccd1 vccd1 hold2371/A sky130_fd_sc_hd__buf_2
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1122 hold1122/A vssd1 vssd1 vccd1 vccd1 _3959_/C sky130_fd_sc_hd__buf_2
Xhold1133 hold2383/X vssd1 vssd1 vccd1 vccd1 hold2384/A sky130_fd_sc_hd__buf_2
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5029_ _5029_/CLK _5029_/D vssd1 vssd1 vccd1 vccd1 _5029_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1177 hold1873/X vssd1 vssd1 vccd1 vccd1 hold1874/A sky130_fd_sc_hd__buf_2
XFILLER_73_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1199 hold1908/X vssd1 vssd1 vccd1 vccd1 hold1909/A sky130_fd_sc_hd__buf_2
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579__164 _4507__92/A vssd1 vssd1 vccd1 vccd1 _5229_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4514__99 _4514__99/A vssd1 vssd1 vccd1 vccd1 _5156_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2390 hold6/X vssd1 vssd1 vccd1 vccd1 hold2390/X sky130_fd_sc_hd__buf_2
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ _3339_/A1 _5497_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5497_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2661_ _3604_/A1 _5585_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5585_/D sky130_fd_sc_hd__mux2_1
X_4400_ _4357_/A _4357_/B _4415_/A3 vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__a21bo_1
XFILLER_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5380_ _5380_/CLK _5380_/D vssd1 vssd1 vccd1 vccd1 _5380_/Q sky130_fd_sc_hd__dfxtp_1
X_2592_ _5694_/Q _5625_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5625_/D sky130_fd_sc_hd__mux2_1
X_4331_ _4080_/A _4080_/B _4279_/X vssd1 vssd1 vccd1 vccd1 _4331_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4262_ _5750_/Q _4262_/B vssd1 vssd1 vccd1 vccd1 _4262_/Y sky130_fd_sc_hd__xnor2_1
X_3213_ _3355_/B _3213_/B vssd1 vssd1 vccd1 vccd1 _3213_/X sky130_fd_sc_hd__and2_1
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _5543_/Q _4187_/B1 _4210_/C _4133_/B vssd1 vssd1 vccd1 vccd1 _4194_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3144_ _5715_/Q _5464_/Q _5448_/Q _5480_/Q _3299_/S _3184_/S1 vssd1 vssd1 vccd1 vccd1
+ _3145_/B sky130_fd_sc_hd__mux4_2
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3075_ _2883_/X _3071_/Y _3074_/Y _3075_/B1 vssd1 vssd1 vccd1 vccd1 _3075_/X sky130_fd_sc_hd__a31o_2
XFILLER_95_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3977_ _3642_/A _5247_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _5247_/D sky130_fd_sc_hd__mux2_1
X_2928_ _2917_/X _2918_/X _2947_/S vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__mux2_1
X_5716_ _5716_/CLK _5716_/D vssd1 vssd1 vccd1 vccd1 _5716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2859_ _5386_/Q _3395_/A0 _2860_/S vssd1 vssd1 vccd1 vccd1 _5386_/D sky130_fd_sc_hd__mux2_1
X_5647_ _5647_/CLK _5647_/D vssd1 vssd1 vccd1 vccd1 _5647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5578_ _5578_/CLK _5578_/D vssd1 vssd1 vccd1 vccd1 _5578_/Q sky130_fd_sc_hd__dfxtp_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__buf_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XCaravelHost_692 vssd1 vssd1 vccd1 vccd1 CaravelHost_692/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XCaravelHost_681 vssd1 vssd1 vccd1 vccd1 CaravelHost_681/HI la_data_out[109] sky130_fd_sc_hd__conb_1
XCaravelHost_670 vssd1 vssd1 vccd1 vccd1 CaravelHost_670/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__buf_2
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold285 hold353/X vssd1 vssd1 vccd1 vccd1 hold354/A sky130_fd_sc_hd__buf_2
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold296 _3623_/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__buf_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3900_ _4399_/B _3898_/X _3899_/X vssd1 vssd1 vccd1 vccd1 _5074_/D sky130_fd_sc_hd__a21o_1
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _4351_/B _4357_/B _3832_/A3 _4361_/A vssd1 vssd1 vccd1 vccd1 _3831_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3762_ _5008_/Q _3774_/A2 _3753_/X _3761_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3762_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5501_ _5501_/CLK _5501_/D vssd1 vssd1 vccd1 vccd1 _5501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3693_ _4984_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__or2_1
X_2713_ _3370_/A _2740_/B vssd1 vssd1 vccd1 vccd1 _2721_/S sky130_fd_sc_hd__or2_4
XFILLER_145_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2644_ _5599_/Q _3606_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5599_/D sky130_fd_sc_hd__mux2_1
X_5432_ _5432_/CLK _5432_/D vssd1 vssd1 vccd1 vccd1 _5432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5363_ _5730_/CLK _5363_/D vssd1 vssd1 vccd1 vccd1 _5363_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput335 _5902_/X vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_12
Xoutput302 _5872_/X vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_12
Xoutput313 _5882_/X vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_12
X_2575_ _5331_/Q _3350_/B split3/A _5332_/Q vssd1 vssd1 vccd1 vccd1 _3397_/A sky130_fd_sc_hd__or4bb_4
Xoutput324 _5892_/X vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_12
XFILLER_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _4266_/B _4318_/A2 _4322_/B _4027_/A vssd1 vssd1 vccd1 vccd1 _4314_/X sky130_fd_sc_hd__o22a_1
Xoutput368 _5932_/X vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_12
Xoutput357 _5922_/X vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_12
Xoutput346 _5912_/X vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_12
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput379 _3736_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__clkbuf_2
X_5294_ _5294_/CLK _5294_/D vssd1 vssd1 vccd1 vccd1 _5294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4245_ _5664_/Q _5663_/Q vssd1 vssd1 vccd1 vccd1 _4269_/A sky130_fd_sc_hd__nand2b_1
X_4948__533 _4964__549/A vssd1 vssd1 vccd1 vccd1 _5706_/CLK sky130_fd_sc_hd__inv_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4176_ _5529_/Q _4186_/B vssd1 vssd1 vccd1 vccd1 _4178_/C sky130_fd_sc_hd__nand2_1
XFILLER_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3127_ _3127_/A _3290_/S vssd1 vssd1 vccd1 vccd1 _3127_/X sky130_fd_sc_hd__or2_1
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3058_ _5449_/Q _5567_/Q _3063_/S vssd1 vssd1 vccd1 vccd1 _3058_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout551 _4099_/X vssd1 vssd1 vccd1 vccd1 _4108_/B sky130_fd_sc_hd__clkbuf_4
Xfanout540 _5326_/Q vssd1 vssd1 vccd1 vccd1 _3327_/S sky130_fd_sc_hd__clkbuf_16
Xfanout573 _3218_/A1 vssd1 vssd1 vccd1 vccd1 _3575_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout562 _3572_/A0 vssd1 vssd1 vccd1 vccd1 _3159_/A sky130_fd_sc_hd__clkbuf_8
Xfanout584 _5693_/Q vssd1 vssd1 vccd1 vccd1 _3395_/A0 sky130_fd_sc_hd__buf_6
Xfanout595 _2897_/A1 vssd1 vssd1 vccd1 vccd1 _3536_/A0 sky130_fd_sc_hd__buf_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741__326 _5010_/CLK vssd1 vssd1 vccd1 vccd1 _5432_/CLK sky130_fd_sc_hd__inv_2
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4635__220 _5684_/CLK vssd1 vssd1 vccd1 vccd1 _5313_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4030_ _5674_/Q _4052_/B _4020_/X vssd1 vssd1 vccd1 vccd1 _4249_/B sky130_fd_sc_hd__o21bai_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_14 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_47 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _5265_/Q hold358/X _3814_/A3 _3814_/B1 _5014_/Q vssd1 vssd1 vccd1 vccd1 _5014_/D
+ sky130_fd_sc_hd__o32a_1
XANTENNA_25 _3772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 hold968/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_69 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ _3824_/A1 _3743_/X _3744_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3745_/X sky130_fd_sc_hd__o211a_4
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _5249_/Q _3682_/B vssd1 vssd1 vccd1 vccd1 _3676_/X sky130_fd_sc_hd__and2_1
X_5415_ _5415_/CLK _5415_/D vssd1 vssd1 vccd1 vccd1 _5415_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_99_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4816__401/A
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_28_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4422__7/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2627_ _2625_/X _2626_/Y _2862_/B vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5346_ _5726_/CLK _5346_/D vssd1 vssd1 vccd1 vccd1 _5346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2558_ _3159_/A _5654_/Q _2565_/S vssd1 vssd1 vccd1 vccd1 _5654_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _5277_/CLK _5277_/D vssd1 vssd1 vccd1 vccd1 _5277_/Q sky130_fd_sc_hd__dfxtp_1
X_2489_ _3350_/A _3350_/B vssd1 vssd1 vccd1 vccd1 _2489_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4228_ _5558_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__or2_1
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4159_ _4167_/B _4167_/C vssd1 vssd1 vccd1 vccd1 _4160_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4619__204 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5296_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_2
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _3767_/A sky130_fd_sc_hd__clkbuf_2
X_3530_ _5134_/Q _3611_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5134_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput45 probe_out[18] vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__clkbuf_2
Xinput89 probe_out[58] vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__clkbuf_2
Xinput78 probe_out[48] vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__clkbuf_2
Xinput67 probe_out[38] vssd1 vssd1 vccd1 vccd1 _5875_/A sky130_fd_sc_hd__clkbuf_2
Xinput56 probe_out[28] vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__clkbuf_2
X_3461_ _3614_/A1 _5195_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5195_/D sky130_fd_sc_hd__mux2_1
X_5200_ _5200_/CLK _5200_/D vssd1 vssd1 vccd1 vccd1 _5200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3392_ _3392_/A0 _5286_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5286_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5131_ _5131_/CLK _5131_/D vssd1 vssd1 vccd1 vccd1 _5131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2208 hold2208/A vssd1 vssd1 vccd1 vccd1 hold2208/X sky130_fd_sc_hd__buf_2
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2219 hold2219/A vssd1 vssd1 vccd1 vccd1 hold2219/X sky130_fd_sc_hd__buf_2
X_5062_ _5062_/CLK _5062_/D vssd1 vssd1 vccd1 vccd1 _5062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1507 hold976/X vssd1 vssd1 vccd1 vccd1 _3937_/A0 sky130_fd_sc_hd__buf_2
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4013_ _4013_/A _4013_/B _4032_/B vssd1 vssd1 vccd1 vccd1 _4247_/B sky130_fd_sc_hd__or3b_4
Xhold1529 hold993/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__buf_2
Xhold1518 hold28/X vssd1 vssd1 vccd1 vccd1 hold982/A sky130_fd_sc_hd__buf_2
X_4910__495 _4449__34/A vssd1 vssd1 vccd1 vccd1 _5631_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5895_ _5895_/A vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3728_ _5079_/Q input7/X _3728_/S vssd1 vssd1 vccd1 vccd1 _3728_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3659_ _3659_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__or2_1
XFILLER_121_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5329_ _5329_/CLK _5329_/D vssd1 vssd1 vccd1 vccd1 _5329_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2731 hold2731/A vssd1 vssd1 vccd1 vccd1 hold2731/X sky130_fd_sc_hd__buf_2
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2720 _3782_/A vssd1 vssd1 vccd1 vccd1 hold2720/X sky130_fd_sc_hd__buf_2
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2764 _4373_/X vssd1 vssd1 vccd1 vccd1 hold2764/X sky130_fd_sc_hd__buf_2
Xhold2797 hold2797/A vssd1 vssd1 vccd1 vccd1 hold2797/X sky130_fd_sc_hd__buf_2
XFILLER_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4853__438 _5106_/CLK vssd1 vssd1 vccd1 vccd1 _5574_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4747__332 _5006_/CLK vssd1 vssd1 vccd1 vccd1 _5438_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2961_ _5117_/Q _3041_/A2 _2945_/A _2960_/X vssd1 vssd1 vccd1 vccd1 _2981_/C sky130_fd_sc_hd__o211a_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5680_ _5683_/CLK _5680_/D vssd1 vssd1 vccd1 vccd1 _5680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2892_ _3073_/C1 _2889_/X _2891_/X vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__a21o_2
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3513_ _3594_/A1 _5149_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5149_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3444_ _3607_/A _3526_/B vssd1 vssd1 vccd1 vccd1 _3452_/S sky130_fd_sc_hd__or2_4
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 hold2670/X vssd1 vssd1 vccd1 vccd1 hold2671/A sky130_fd_sc_hd__buf_2
Xhold2005 hold2643/X vssd1 vssd1 vccd1 vccd1 hold2644/A sky130_fd_sc_hd__buf_2
X_3375_ _3567_/A1 _5304_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5304_/D sky130_fd_sc_hd__mux2_1
X_5114_ _5114_/CLK _5114_/D vssd1 vssd1 vccd1 vccd1 _5114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2049 hold180/X vssd1 vssd1 vccd1 vccd1 hold2049/X sky130_fd_sc_hd__buf_2
Xhold1304 hold458/X vssd1 vssd1 vccd1 vccd1 _4390_/C sky130_fd_sc_hd__buf_2
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 hold2609/X vssd1 vssd1 vccd1 vccd1 hold1978/A sky130_fd_sc_hd__buf_2
XFILLER_73_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/CLK _5045_/D vssd1 vssd1 vccd1 vccd1 _5045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540__125 _4423__8/A vssd1 vssd1 vccd1 vccd1 _5182_/CLK sky130_fd_sc_hd__inv_2
X_5878_ _5878_/A vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_43_wb_clk_i _4676__261/A vssd1 vssd1 vccd1 vccd1 _4425__10/A sky130_fd_sc_hd__clkbuf_16
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput202 hold129/X vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2572 _4358_/Y vssd1 vssd1 vccd1 vccd1 hold2572/X sky130_fd_sc_hd__buf_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2583 _4361_/Y vssd1 vssd1 vccd1 vccd1 hold2583/X sky130_fd_sc_hd__buf_2
Xhold2550 hold2550/A vssd1 vssd1 vccd1 vccd1 hold2550/X sky130_fd_sc_hd__buf_2
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1871 hold2744/X vssd1 vssd1 vccd1 vccd1 hold1871/X sky130_fd_sc_hd__buf_2
Xhold2594 hold205/X vssd1 vssd1 vccd1 vccd1 hold2594/X sky130_fd_sc_hd__buf_2
Xhold1860 hold194/X vssd1 vssd1 vccd1 vccd1 hold1860/X sky130_fd_sc_hd__buf_2
XFILLER_91_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1882 hold2748/X vssd1 vssd1 vccd1 vccd1 hold1882/X sky130_fd_sc_hd__buf_2
Xhold1893 hold2752/X vssd1 vssd1 vccd1 vccd1 hold1893/X sky130_fd_sc_hd__buf_2
XFILLER_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3160_ _3156_/X _3158_/X _3159_/X _4093_/B vssd1 vssd1 vccd1 vccd1 _5344_/D sky130_fd_sc_hd__o211a_1
X_3091_ _3091_/A _3091_/B vssd1 vssd1 vccd1 vccd1 _5370_/D sky130_fd_sc_hd__nor2_1
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3993_ _5261_/Q _3656_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _3993_/X sky130_fd_sc_hd__mux2_1
X_4524__109 _4478__63/A vssd1 vssd1 vccd1 vccd1 _5166_/CLK sky130_fd_sc_hd__inv_2
X_5732_ _5751_/CLK _5732_/D vssd1 vssd1 vccd1 vccd1 _5732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2944_ _5030_/Q _5174_/Q _5238_/Q _5222_/Q _2944_/S0 _3040_/S vssd1 vssd1 vccd1 vccd1
+ _2945_/B sky130_fd_sc_hd__mux4_2
X_2875_ _2883_/B _2875_/B vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__or2_4
X_5663_ _5683_/CLK _5663_/D vssd1 vssd1 vccd1 vccd1 _5663_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4875__460 _4875__460/A vssd1 vssd1 vccd1 vccd1 _5596_/CLK sky130_fd_sc_hd__inv_2
X_5594_ _5594_/CLK _5594_/D vssd1 vssd1 vccd1 vccd1 _5594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold401 hold401/A vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__buf_2
XFILLER_144_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold445 hold445/A vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__buf_2
XFILLER_143_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3427_ _5232_/Q _3591_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5232_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold489 hold489/A vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__buf_2
XFILLER_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3358_ _3130_/B _3357_/A _3357_/Y _4093_/B vssd1 vssd1 vccd1 vccd1 _5327_/D sky130_fd_sc_hd__o211a_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1123 _3959_/X vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__buf_2
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3289_ _3325_/A _3287_/X _3288_/X vssd1 vssd1 vccd1 vccd1 _3289_/X sky130_fd_sc_hd__o21a_1
X_5028_ _5028_/CLK _5028_/D vssd1 vssd1 vccd1 vccd1 _5028_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1178 hold1875/X vssd1 vssd1 vccd1 vccd1 hold1876/A sky130_fd_sc_hd__buf_2
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold990 hold990/A vssd1 vssd1 vccd1 vccd1 hold990/X sky130_fd_sc_hd__buf_2
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2380 hold2380/A vssd1 vssd1 vccd1 vccd1 hold2380/X sky130_fd_sc_hd__buf_2
Xhold2391 hold2391/A vssd1 vssd1 vccd1 vccd1 hold986/A sky130_fd_sc_hd__buf_2
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859__444 _4875__460/A vssd1 vssd1 vccd1 vccd1 _5580_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2660_ _3603_/A1 _5586_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5586_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2591_ _3393_/A0 _5626_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5626_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4330_ _5682_/Q _4325_/Y _4329_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _5682_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4261_ _5751_/Q _4261_/B vssd1 vssd1 vccd1 vccd1 _4261_/Y sky130_fd_sc_hd__xnor2_1
X_3212_ _5712_/Q _5461_/Q _5445_/Q _5477_/Q _3330_/S _3219_/S0 vssd1 vssd1 vccd1 vccd1
+ _3213_/B sky130_fd_sc_hd__mux4_2
X_4192_ _4204_/A _4192_/B vssd1 vssd1 vccd1 vccd1 _4192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3143_ _5416_/Q _5392_/Q _5662_/Q _5424_/Q _3327_/S _3184_/S1 vssd1 vssd1 vccd1 vccd1
+ _3143_/X sky130_fd_sc_hd__mux4_1
X_3074_ _3074_/A1 _3072_/X _3073_/X vssd1 vssd1 vccd1 vccd1 _3074_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3976_ _4389_/A _5246_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _3976_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2927_ _2947_/S _2922_/X _2919_/B vssd1 vssd1 vccd1 vccd1 _2927_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5715_ _5715_/CLK _5715_/D vssd1 vssd1 vccd1 vccd1 _5715_/Q sky130_fd_sc_hd__dfxtp_1
X_5646_ _5646_/CLK _5646_/D vssd1 vssd1 vccd1 vccd1 _5646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2858_ _5387_/Q _3394_/A0 _2860_/S vssd1 vssd1 vccd1 vccd1 _5387_/D sky130_fd_sc_hd__mux2_1
Xhold220 _3993_/X vssd1 vssd1 vccd1 vccd1 _5261_/D sky130_fd_sc_hd__buf_2
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5577_ _5577_/CLK _5577_/D vssd1 vssd1 vccd1 vccd1 _5577_/Q sky130_fd_sc_hd__dfxtp_1
X_2789_ _2853_/A1 _5448_/Q _2796_/S vssd1 vssd1 vccd1 vccd1 _5448_/D sky130_fd_sc_hd__mux2_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__buf_2
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XCaravelHost_682 vssd1 vssd1 vccd1 vccd1 CaravelHost_682/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XCaravelHost_671 vssd1 vssd1 vccd1 vccd1 CaravelHost_671/HI la_data_out[99] sky130_fd_sc_hd__conb_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__buf_2
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XCaravelHost_660 vssd1 vssd1 vccd1 vccd1 CaravelHost_660/HI core0Index[5] sky130_fd_sc_hd__conb_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__buf_2
Xhold286 hold355/X vssd1 vssd1 vccd1 vccd1 hold356/A sky130_fd_sc_hd__buf_2
XCaravelHost_693 vssd1 vssd1 vccd1 vccd1 CaravelHost_693/HI la_data_out[121] sky130_fd_sc_hd__conb_1
X_4652__237 _4459__44/A vssd1 vssd1 vccd1 vccd1 _5338_/CLK sky130_fd_sc_hd__inv_2
XFILLER_131_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__buf_2
XFILLER_86_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4546__131 _4418__3/A vssd1 vssd1 vccd1 vccd1 _5188_/CLK sky130_fd_sc_hd__inv_2
XFILLER_121_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3830_ _3829_/X _3830_/B vssd1 vssd1 vccd1 vccd1 _3830_/X sky130_fd_sc_hd__and2b_1
X_3761_ _3761_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3761_/X sky130_fd_sc_hd__and2_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5500_ _5500_/CLK _5500_/D vssd1 vssd1 vccd1 vccd1 _5500_/Q sky130_fd_sc_hd__dfxtp_1
X_2712_ _5335_/Q _5334_/Q _3346_/A vssd1 vssd1 vccd1 vccd1 _2740_/B sky130_fd_sc_hd__or3b_4
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3692_ _5067_/Q input14/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3692_/X sky130_fd_sc_hd__mux2_4
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2643_ _5600_/Q _3605_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5600_/D sky130_fd_sc_hd__mux2_1
X_5431_ _5431_/CLK _5431_/D vssd1 vssd1 vccd1 vccd1 _5431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5362_ _5362_/CLK _5362_/D vssd1 vssd1 vccd1 vccd1 _5362_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput325 _5893_/X vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_12
Xoutput314 _5883_/X vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_12
X_2574_ _3579_/A0 _5639_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5639_/D sky130_fd_sc_hd__mux2_1
Xoutput303 _5873_/X vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_12
XFILLER_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4313_ _4312_/X _4315_/B vssd1 vssd1 vccd1 vccd1 _4313_/X sky130_fd_sc_hd__and2b_1
Xoutput369 _5933_/X vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_12
Xoutput358 _5923_/X vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_12
Xoutput336 _5903_/X vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_12
Xoutput347 _5913_/X vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_12
X_5293_ _5293_/CLK _5293_/D vssd1 vssd1 vccd1 vccd1 _5293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4244_ _5566_/Q _4164_/B _4244_/S vssd1 vssd1 vccd1 vccd1 _5566_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4175_ _4165_/B _4186_/B _4242_/B _5529_/Q vssd1 vssd1 vccd1 vccd1 _4178_/B sky130_fd_sc_hd__a211o_1
XFILLER_68_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3126_ _3126_/A _3290_/S vssd1 vssd1 vccd1 vccd1 _3128_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3057_ _3099_/B _3055_/X _3056_/X vssd1 vssd1 vccd1 vccd1 _3057_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3959_ _3959_/A _3959_/B _3959_/C vssd1 vssd1 vccd1 vccd1 _3959_/X sky130_fd_sc_hd__or3_1
XFILLER_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5629_ _5629_/CLK _5629_/D vssd1 vssd1 vccd1 vccd1 _5629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout541 _3312_/S vssd1 vssd1 vccd1 vccd1 _3281_/S sky130_fd_sc_hd__clkbuf_16
Xfanout530 _2482_/B vssd1 vssd1 vccd1 vccd1 _2464_/A sky130_fd_sc_hd__buf_6
Xfanout552 _4021_/C vssd1 vssd1 vccd1 vccd1 _4065_/B sky130_fd_sc_hd__buf_6
XFILLER_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout574 _3218_/A1 vssd1 vssd1 vccd1 vccd1 _3566_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout563 _5699_/Q vssd1 vssd1 vccd1 vccd1 _3572_/A0 sky130_fd_sc_hd__buf_4
XFILLER_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout596 _5325_/Q vssd1 vssd1 vccd1 vccd1 _2897_/A1 sky130_fd_sc_hd__buf_6
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout585 _3308_/A1 vssd1 vssd1 vccd1 vccd1 _3569_/A1 sky130_fd_sc_hd__buf_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4780__365 _5022_/CLK vssd1 vssd1 vccd1 vccd1 _5471_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4495__80 _4422__7/A vssd1 vssd1 vccd1 vccd1 _5137_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _5264_/Q hold358/X _3814_/A3 _3814_/B1 _5013_/Q vssd1 vssd1 vccd1 vccd1 _3813_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_48 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 _3639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _3774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 hold30/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_59 _3662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3744_ _5001_/Q _3750_/B vssd1 vssd1 vccd1 vccd1 _3744_/X sky130_fd_sc_hd__or2_1
XFILLER_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3675_ _3675_/A _3682_/B vssd1 vssd1 vccd1 vccd1 _3675_/X sky130_fd_sc_hd__and2_1
XFILLER_118_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4915__500 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5636_/CLK sky130_fd_sc_hd__inv_2
XFILLER_146_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2626_ _2625_/A _5367_/Q _3081_/A vssd1 vssd1 vccd1 vccd1 _2626_/Y sky130_fd_sc_hd__a21oi_1
X_5414_ _5414_/CLK _5414_/D vssd1 vssd1 vccd1 vccd1 _5414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5345_ _5751_/CLK _5345_/D vssd1 vssd1 vccd1 vccd1 _5345_/Q sky130_fd_sc_hd__dfxtp_4
X_2557_ _3370_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _2565_/S sky130_fd_sc_hd__or2_4
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5276_ _5276_/CLK _5276_/D vssd1 vssd1 vccd1 vccd1 _5276_/Q sky130_fd_sc_hd__dfxtp_1
X_2488_ _5345_/Q _4361_/B vssd1 vssd1 vccd1 vccd1 _3350_/B sky130_fd_sc_hd__nand2_8
Xclkbuf_leaf_68_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4485__70/A
+ sky130_fd_sc_hd__clkbuf_16
X_4227_ _4225_/X _4226_/X _4217_/A vssd1 vssd1 vccd1 vccd1 _5557_/D sky130_fd_sc_hd__a21oi_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4158_ _5545_/Q _5544_/Q _5543_/Q _4132_/B _5546_/Q vssd1 vssd1 vccd1 vccd1 _4167_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4764__349 _5252_/CLK vssd1 vssd1 vccd1 vccd1 _5455_/CLK sky130_fd_sc_hd__inv_2
X_3109_ _5357_/Q _3604_/A1 _3111_/S vssd1 vssd1 vccd1 vccd1 _5357_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4089_ _5690_/Q _4094_/C vssd1 vssd1 vccd1 vccd1 _4089_/X sky130_fd_sc_hd__and2_1
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4658__243 _4658__243/A vssd1 vssd1 vccd1 vccd1 _5344_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__clkbuf_2
Xinput35 caravel_wb_error_i vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput46 probe_out[19] vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput79 probe_out[49] vssd1 vssd1 vccd1 vccd1 _5886_/A sky130_fd_sc_hd__clkbuf_2
Xinput68 probe_out[39] vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__clkbuf_2
Xinput57 probe_out[29] vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3460_ _3613_/A1 _5196_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5196_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3391_ _3391_/A0 _5287_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5287_/D sky130_fd_sc_hd__mux2_4
X_5130_ _5130_/CLK _5130_/D vssd1 vssd1 vccd1 vccd1 _5130_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2209 hold2209/A vssd1 vssd1 vccd1 vccd1 _4966_/D sky130_fd_sc_hd__buf_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5061_ _5061_/CLK _5061_/D vssd1 vssd1 vccd1 vccd1 _5061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1508 _3937_/X vssd1 vssd1 vccd1 vccd1 hold977/A sky130_fd_sc_hd__buf_2
XFILLER_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4012_ _4027_/A _4011_/A _4065_/B _4029_/C vssd1 vssd1 vccd1 vccd1 _4032_/B sky130_fd_sc_hd__and4bb_4
Xhold1519 hold982/X vssd1 vssd1 vccd1 vccd1 _3938_/A0 sky130_fd_sc_hd__buf_2
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5894_ _5894_/A vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_115_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5244_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3727_ _3733_/A1 _3725_/X _3726_/X split2/A vssd1 vssd1 vccd1 vccd1 _3727_/X sky130_fd_sc_hd__o211a_1
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3658_ _3658_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__or2_1
X_3589_ _3589_/A _3589_/B vssd1 vssd1 vccd1 vccd1 _3597_/S sky130_fd_sc_hd__nor2_8
X_2609_ _3575_/A0 _5611_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5611_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5328_ _5328_/CLK _5328_/D vssd1 vssd1 vccd1 vccd1 _5328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5259_ _5259_/CLK _5259_/D vssd1 vssd1 vccd1 vccd1 _5259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2798 hold2798/A vssd1 vssd1 vccd1 vccd1 hold2798/X sky130_fd_sc_hd__buf_2
Xhold2787 hold2884/X vssd1 vssd1 vccd1 vccd1 hold2885/A sky130_fd_sc_hd__buf_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4892__477 _4892__477/A vssd1 vssd1 vccd1 vccd1 _5613_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4786__371 _4786__371/A vssd1 vssd1 vccd1 vccd1 _5477_/CLK sky130_fd_sc_hd__inv_2
X_4465__50 _4424__9/A vssd1 vssd1 vccd1 vccd1 _5059_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4424__9 _4424__9/A vssd1 vssd1 vccd1 vccd1 _4975_/CLK sky130_fd_sc_hd__inv_2
X_2960_ _5229_/Q _2870_/B _2959_/X _3041_/B1 vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__o22a_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2891_ _3029_/B1 _2890_/X _2919_/B vssd1 vssd1 vccd1 vccd1 _2891_/X sky130_fd_sc_hd__a21o_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3512_ _3611_/A1 _5150_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5150_/D sky130_fd_sc_hd__mux2_1
X_3443_ _5373_/Q _3443_/B _3453_/C vssd1 vssd1 vccd1 vccd1 _3526_/B sky130_fd_sc_hd__or3b_4
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3374_ _3575_/A0 _5305_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5305_/D sky130_fd_sc_hd__mux2_1
X_5113_ _5754_/CLK _5113_/D vssd1 vssd1 vccd1 vccd1 _5113_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 hold2645/X vssd1 vssd1 vccd1 vccd1 hold2646/A sky130_fd_sc_hd__buf_2
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1305 hold2626/X vssd1 vssd1 vccd1 vccd1 hold2627/A sky130_fd_sc_hd__buf_2
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 hold2686/X vssd1 vssd1 vccd1 vccd1 hold2687/A sky130_fd_sc_hd__buf_2
Xhold2028 hold2672/X vssd1 vssd1 vccd1 vccd1 hold2673/A sky130_fd_sc_hd__buf_2
XFILLER_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1327 hold2634/X vssd1 vssd1 vccd1 vccd1 hold2635/A sky130_fd_sc_hd__buf_2
X_5044_ _5044_/CLK _5044_/D vssd1 vssd1 vccd1 vccd1 _5044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5877_ _5877_/A vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4961__546/A sky130_fd_sc_hd__clkbuf_16
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_wb_clk_i _4676__261/A vssd1 vssd1 vccd1 vccd1 _5725_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2540 hold848/X vssd1 vssd1 vccd1 vccd1 hold2540/X sky130_fd_sc_hd__buf_2
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput203 hold224/X vssd1 vssd1 vccd1 vccd1 _3628_/A sky130_fd_sc_hd__buf_4
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2573 hold2573/A vssd1 vssd1 vccd1 vccd1 hold2573/X sky130_fd_sc_hd__buf_2
XFILLER_84_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2551 hold2551/A vssd1 vssd1 vccd1 vccd1 hold2551/X sky130_fd_sc_hd__buf_2
Xhold2562 _4412_/X vssd1 vssd1 vccd1 vccd1 hold2562/X sky130_fd_sc_hd__buf_2
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1850 hold1850/A vssd1 vssd1 vccd1 vccd1 _5738_/D sky130_fd_sc_hd__buf_2
Xhold1872 hold1872/A vssd1 vssd1 vccd1 vccd1 hold584/A sky130_fd_sc_hd__buf_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2584 hold2584/A vssd1 vssd1 vccd1 vccd1 hold2584/X sky130_fd_sc_hd__buf_2
Xhold2595 hold2595/A vssd1 vssd1 vccd1 vccd1 hold2595/X sky130_fd_sc_hd__buf_2
Xhold1861 hold1861/A vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__buf_2
Xhold1883 hold1883/A vssd1 vssd1 vccd1 vccd1 hold867/A sky130_fd_sc_hd__buf_2
Xhold1894 hold1894/A vssd1 vssd1 vccd1 vccd1 hold841/A sky130_fd_sc_hd__buf_2
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820__405 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5511_/CLK sky130_fd_sc_hd__inv_2
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3090_ _5370_/Q _3093_/A _2778_/A vssd1 vssd1 vccd1 vccd1 _3091_/B sky130_fd_sc_hd__o21ai_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _5260_/Q _3655_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2943_ _5198_/Q _5182_/Q _4971_/Q _5190_/Q _3036_/S _2943_/S1 vssd1 vssd1 vccd1 vccd1
+ _2943_/X sky130_fd_sc_hd__mux4_2
X_4563__148 _4507__92/A vssd1 vssd1 vccd1 vccd1 _5213_/CLK sky130_fd_sc_hd__inv_2
X_5731_ _5731_/CLK _5731_/D vssd1 vssd1 vccd1 vccd1 _5731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2874_ _2883_/B _2875_/B vssd1 vssd1 vccd1 vccd1 _2874_/Y sky130_fd_sc_hd__nor2_2
X_5662_ _5662_/CLK _5662_/D vssd1 vssd1 vccd1 vccd1 _5662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4604__189 _5565_/CLK vssd1 vssd1 vccd1 vccd1 _5278_/CLK sky130_fd_sc_hd__inv_2
X_5593_ _5593_/CLK _5593_/D vssd1 vssd1 vccd1 vccd1 _5593_/Q sky130_fd_sc_hd__dfxtp_1
Xhold402 hold402/A vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__buf_2
XFILLER_143_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold468 hold824/X vssd1 vssd1 vccd1 vccd1 hold825/A sky130_fd_sc_hd__buf_2
X_3426_ _5233_/Q _3608_/A1 _3433_/S vssd1 vssd1 vccd1 vccd1 _5233_/D sky130_fd_sc_hd__mux2_1
Xhold479 hold499/X vssd1 vssd1 vccd1 vccd1 hold500/A sky130_fd_sc_hd__buf_2
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3357_ _3357_/A _3357_/B vssd1 vssd1 vccd1 vccd1 _3357_/Y sky130_fd_sc_hd__nand2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1124 hold199/X vssd1 vssd1 vccd1 vccd1 _3960_/C sky130_fd_sc_hd__buf_2
Xhold1113 hold2353/X vssd1 vssd1 vccd1 vccd1 hold2354/A sky130_fd_sc_hd__buf_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5027_/CLK _5027_/D vssd1 vssd1 vccd1 vccd1 _5027_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1157 hold2227/X vssd1 vssd1 vccd1 vccd1 hold2228/A sky130_fd_sc_hd__buf_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3288_ _5616_/Q _2464_/A _3326_/B2 _5608_/Q _3316_/C1 vssd1 vssd1 vccd1 vccd1 _3288_/X
+ sky130_fd_sc_hd__o221a_1
Xhold1179 hold1877/X vssd1 vssd1 vccd1 vccd1 hold1878/A sky130_fd_sc_hd__buf_2
XFILLER_54_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5929_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_126_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold991 hold991/A vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__buf_2
Xhold980 hold980/A vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__buf_2
XFILLER_122_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2381 hold2381/A vssd1 vssd1 vccd1 vccd1 hold909/A sky130_fd_sc_hd__buf_2
XFILLER_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2370 hold2370/A vssd1 vssd1 vccd1 vccd1 hold2370/X sky130_fd_sc_hd__buf_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2392 hold986/X vssd1 vssd1 vccd1 vccd1 hold2392/X sky130_fd_sc_hd__buf_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4435__20 _4435__20/A vssd1 vssd1 vccd1 vccd1 _5029_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4898__483 _4898__483/A vssd1 vssd1 vccd1 vccd1 _5619_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _3392_/A0 _5627_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5627_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _4260_/A _4260_/B _4260_/C _4260_/D vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__or4_1
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4191_ _5542_/Q _4187_/B1 _4210_/C _4135_/B vssd1 vssd1 vccd1 vccd1 _4192_/B sky130_fd_sc_hd__o2bb2a_1
X_3211_ _5413_/Q _5389_/Q _5659_/Q _5421_/Q _3327_/S _3219_/S0 vssd1 vssd1 vccd1 vccd1
+ _3211_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3142_ _5614_/Q _5598_/Q _5582_/Q _5622_/Q _3284_/S _3201_/S1 vssd1 vssd1 vccd1 vccd1
+ _3142_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3073_ _2460_/A _5355_/Q _5122_/Q _3073_/B2 _3073_/C1 vssd1 vssd1 vccd1 vccd1 _3073_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3975_ _3640_/A _5245_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _5245_/D sky130_fd_sc_hd__mux2_1
X_2926_ _5430_/Q _5406_/Q _5398_/Q _5438_/Q _3069_/S _2942_/S1 vssd1 vssd1 vccd1 vccd1
+ _2926_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5714_ _5714_/CLK _5714_/D vssd1 vssd1 vccd1 vccd1 _5714_/Q sky130_fd_sc_hd__dfxtp_1
X_2857_ _5388_/Q _3402_/A1 _2860_/S vssd1 vssd1 vccd1 vccd1 _5388_/D sky130_fd_sc_hd__mux2_1
X_5645_ _5645_/CLK _5645_/D vssd1 vssd1 vccd1 vccd1 _5645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold210 hold237/X vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__buf_2
X_5576_ _5576_/CLK _5576_/D vssd1 vssd1 vccd1 vccd1 _5576_/Q sky130_fd_sc_hd__dfxtp_1
X_2788_ _2788_/A _3571_/A vssd1 vssd1 vccd1 vccd1 _2796_/S sky130_fd_sc_hd__or2_4
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 _3997_/S sky130_fd_sc_hd__buf_2
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XCaravelHost_683 vssd1 vssd1 vccd1 vccd1 CaravelHost_683/HI la_data_out[111] sky130_fd_sc_hd__conb_1
XCaravelHost_672 vssd1 vssd1 vccd1 vccd1 CaravelHost_672/HI la_data_out[100] sky130_fd_sc_hd__conb_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__buf_2
Xhold221 hold234/X vssd1 vssd1 vccd1 vccd1 hold235/A sky130_fd_sc_hd__buf_2
XCaravelHost_661 vssd1 vssd1 vccd1 vccd1 CaravelHost_661/HI core0Index[6] sky130_fd_sc_hd__conb_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__buf_2
Xhold287 hold357/X vssd1 vssd1 vccd1 vccd1 hold358/A sky130_fd_sc_hd__buf_2
X_4691__276 _5384_/CLK vssd1 vssd1 vccd1 vccd1 _5380_/CLK sky130_fd_sc_hd__inv_2
XCaravelHost_694 vssd1 vssd1 vccd1 vccd1 CaravelHost_694/HI la_data_out[122] sky130_fd_sc_hd__conb_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__buf_2
XFILLER_131_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3409_ _5271_/Q _3409_/A1 _3414_/S vssd1 vssd1 vccd1 vccd1 _5271_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__buf_2
XFILLER_112_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4389_ _4389_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4389_/X sky130_fd_sc_hd__and3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4585__170 _4435__20/A vssd1 vssd1 vccd1 vccd1 _5235_/CLK sky130_fd_sc_hd__inv_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4932__517 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5653_/CLK sky130_fd_sc_hd__inv_2
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4826__411 _5019_/CLK vssd1 vssd1 vccd1 vccd1 _5517_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _5007_/Q _3750_/B _3774_/B1 _3759_/X _3774_/C1 vssd1 vssd1 vccd1 vccd1 _3760_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_60_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2711_ _3396_/A0 _5513_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5513_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5430_ _5430_/CLK _5430_/D vssd1 vssd1 vccd1 vccd1 _5430_/Q sky130_fd_sc_hd__dfxtp_1
X_3691_ _3718_/A1 _3689_/X _3690_/X split4/X vssd1 vssd1 vccd1 vccd1 _3691_/X sky130_fd_sc_hd__o211a_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2642_ _5601_/Q _3604_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5601_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5361_ _5361_/CLK _5361_/D vssd1 vssd1 vccd1 vccd1 _5361_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput326 _5894_/X vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_12
X_2573_ _3578_/A0 _5640_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5640_/D sky130_fd_sc_hd__mux2_1
Xoutput304 _5874_/X vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_12
Xoutput315 _5884_/X vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_12
XFILLER_141_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5292_ _5677_/CLK hold53/X vssd1 vssd1 vccd1 vccd1 _5292_/Q sky130_fd_sc_hd__dfxtp_2
X_4312_ _4023_/B _4318_/A2 _4322_/B _2442_/Y vssd1 vssd1 vccd1 vccd1 _4312_/X sky130_fd_sc_hd__o22a_1
Xoutput359 _5924_/X vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_12
Xoutput348 _5914_/X vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_12
Xoutput337 _5904_/X vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_12
X_4243_ _5344_/Q _3124_/Y _4164_/B _4242_/X hold741/X vssd1 vssd1 vccd1 vccd1 _4243_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _4152_/Y _4153_/X _4171_/X _4172_/X _4173_/Y vssd1 vssd1 vccd1 vccd1 _4177_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _3125_/A _4360_/B vssd1 vssd1 vccd1 vccd1 _3125_/Y sky130_fd_sc_hd__nor2_1
X_3056_ _4975_/Q _2866_/A _2866_/B _5058_/Q _3097_/B vssd1 vssd1 vccd1 vccd1 _3056_/X
+ sky130_fd_sc_hd__o221a_1
X_4569__154 _4433__18/A vssd1 vssd1 vccd1 vccd1 _5219_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3958_ _3959_/A _3958_/A2 _3960_/B vssd1 vssd1 vccd1 vccd1 _3958_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2909_ _3029_/B1 _2907_/X _2908_/X vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3889_ _3886_/X _3887_/X _3888_/Y _5749_/Q vssd1 vssd1 vccd1 vccd1 _3889_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5628_ _5628_/CLK _5628_/D vssd1 vssd1 vccd1 vccd1 _5628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5559_ _5564_/CLK _5559_/D vssd1 vssd1 vccd1 vccd1 _5559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout520 _3066_/S vssd1 vssd1 vccd1 vccd1 _3040_/S sky130_fd_sc_hd__buf_6
Xfanout542 fanout547/X vssd1 vssd1 vccd1 vccd1 _3312_/S sky130_fd_sc_hd__buf_6
Xfanout531 _5328_/Q vssd1 vssd1 vccd1 vccd1 _2482_/B sky130_fd_sc_hd__buf_8
Xfanout553 _3797_/A3 vssd1 vssd1 vccd1 vccd1 _3829_/A sky130_fd_sc_hd__buf_6
Xfanout575 _5696_/Q vssd1 vssd1 vccd1 vccd1 _3218_/A1 sky130_fd_sc_hd__buf_4
Xfanout564 _2790_/A0 vssd1 vssd1 vccd1 vccd1 _3390_/A0 sky130_fd_sc_hd__buf_4
XFILLER_132_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout597 _2916_/A1 vssd1 vssd1 vccd1 vccd1 _3591_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout586 _3308_/A1 vssd1 vssd1 vccd1 vccd1 _3578_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3812_ _5263_/Q hold358/X _3814_/A3 _3814_/B1 _5012_/Q vssd1 vssd1 vccd1 vccd1 _5012_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_119_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 _3639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _3796_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 hold39/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_49 _4356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3743_ _5084_/Q input12/X _3763_/B vssd1 vssd1 vccd1 vccd1 _3743_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3674_ _3674_/A _3682_/B vssd1 vssd1 vccd1 vccd1 _3674_/X sky130_fd_sc_hd__and2_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2625_ _2625_/A _5367_/Q _3081_/A vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__or3_1
X_5413_ _5413_/CLK _5413_/D vssd1 vssd1 vccd1 vccd1 _5413_/Q sky130_fd_sc_hd__dfxtp_1
X_5344_ _5344_/CLK _5344_/D vssd1 vssd1 vccd1 vccd1 _5344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2556_ _5334_/Q _3346_/A _5335_/Q vssd1 vssd1 vccd1 vccd1 _3571_/B sky130_fd_sc_hd__or3b_4
XFILLER_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2903 _4410_/X vssd1 vssd1 vccd1 vccd1 hold2903/X sky130_fd_sc_hd__buf_2
X_5275_ _5275_/CLK _5275_/D vssd1 vssd1 vccd1 vccd1 _5275_/Q sky130_fd_sc_hd__dfxtp_1
X_2487_ _2487_/A _2487_/B _2487_/C _2487_/D vssd1 vssd1 vccd1 vccd1 _4361_/B sky130_fd_sc_hd__or4_4
XFILLER_141_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4226_ _5557_/Q _4226_/B _4222_/B _4220_/B vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__or4bb_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4157_ _5746_/Q _4157_/B vssd1 vssd1 vccd1 vccd1 _4157_/X sky130_fd_sc_hd__xor2_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3108_ _5358_/Q _3603_/A1 _3111_/S vssd1 vssd1 vccd1 vccd1 _5358_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4088_ _5689_/Q _4088_/B vssd1 vssd1 vccd1 vccd1 _4088_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4883__468/A
+ sky130_fd_sc_hd__clkbuf_16
X_3039_ _5219_/Q _2873_/B _2870_/B vssd1 vssd1 vccd1 vccd1 _3039_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4697__282 _5244_/CLK vssd1 vssd1 vccd1 vccd1 _5388_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4938__523 _5246_/CLK vssd1 vssd1 vccd1 vccd1 _5659_/CLK sky130_fd_sc_hd__inv_2
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_2
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_2
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput36 probe_out[0] vssd1 vssd1 vccd1 vccd1 _5837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput58 probe_out[2] vssd1 vssd1 vccd1 vccd1 _5839_/A sky130_fd_sc_hd__clkbuf_2
Xinput47 probe_out[1] vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__clkbuf_2
Xinput69 probe_out[3] vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3390_ _3390_/A0 _5288_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5288_/D sky130_fd_sc_hd__mux2_4
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5060_ _5060_/CLK _5060_/D vssd1 vssd1 vccd1 vccd1 _5060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4011_ _4011_/A _4063_/A _4029_/C vssd1 vssd1 vccd1 vccd1 _4027_/B sky130_fd_sc_hd__or3b_4
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1509 hold977/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__buf_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5893_ _5893_/A vssd1 vssd1 vccd1 vccd1 _5893_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3726_ _4995_/Q _3729_/B vssd1 vssd1 vccd1 vccd1 _3726_/X sky130_fd_sc_hd__or2_1
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3657_ _3657_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3657_/X sky130_fd_sc_hd__or2_1
XFILLER_106_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3588_ _3597_/A1 _5034_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5034_/D sky130_fd_sc_hd__mux2_1
X_2608_ _2743_/A0 _5612_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5612_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2539_ _3566_/A1 _5704_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5704_/D sky130_fd_sc_hd__mux2_1
X_4731__316 _4731__316/A vssd1 vssd1 vccd1 vccd1 _5422_/CLK sky130_fd_sc_hd__inv_2
X_5327_ _5327_/CLK _5327_/D vssd1 vssd1 vccd1 vccd1 _5327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5258_ _5259_/CLK _5258_/D vssd1 vssd1 vccd1 vccd1 _5258_/Q sky130_fd_sc_hd__dfxtp_2
Xhold2744 _4379_/X vssd1 vssd1 vccd1 vccd1 hold2744/X sky130_fd_sc_hd__buf_2
XFILLER_75_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5189_ _5189_/CLK _5189_/D vssd1 vssd1 vccd1 vccd1 _5189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2799 hold2799/A vssd1 vssd1 vccd1 vccd1 hold2799/X sky130_fd_sc_hd__buf_2
X_4209_ _5551_/Q _4209_/B vssd1 vssd1 vccd1 vccd1 _4209_/Y sky130_fd_sc_hd__nand2_1
Xhold2788 hold2886/X vssd1 vssd1 vccd1 vccd1 hold2887/A sky130_fd_sc_hd__buf_2
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4625__210 _4457__42/A vssd1 vssd1 vccd1 vccd1 _5302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480__65 _5084_/CLK vssd1 vssd1 vccd1 vccd1 _5122_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2890_ _5432_/Q _5408_/Q _5400_/Q _5440_/Q _3024_/S _2942_/S1 vssd1 vssd1 vccd1 vccd1
+ _2890_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3511_ _3610_/A1 _5151_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5151_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3442_ _5218_/Q _3597_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5218_/D sky130_fd_sc_hd__mux2_1
Xhold628 hold628/A vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__buf_2
XFILLER_143_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3373_ _3574_/A0 _5306_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5306_/D sky130_fd_sc_hd__mux2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5733_/CLK _5112_/D vssd1 vssd1 vccd1 vccd1 _5112_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 hold2007/A vssd1 vssd1 vccd1 vccd1 _4995_/D sky130_fd_sc_hd__buf_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1306 hold2630/X vssd1 vssd1 vccd1 vccd1 hold1995/A sky130_fd_sc_hd__buf_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 hold2674/X vssd1 vssd1 vccd1 vccd1 hold2675/A sky130_fd_sc_hd__buf_2
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 hold2638/X vssd1 vssd1 vccd1 vccd1 hold2001/A sky130_fd_sc_hd__buf_2
Xhold1339 hold2671/X vssd1 vssd1 vccd1 vccd1 hold2672/A sky130_fd_sc_hd__buf_2
X_5043_ _5043_/CLK _5043_/D vssd1 vssd1 vccd1 vccd1 _5043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5876_ _5876_/A vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3709_ _3718_/A1 _3707_/X _3708_/X split4/A vssd1 vssd1 vccd1 vccd1 _3709_/X sky130_fd_sc_hd__o211a_1
XFILLER_108_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2530 hold2530/A vssd1 vssd1 vccd1 vccd1 _5322_/D sky130_fd_sc_hd__buf_2
Xinput204 hold295/X vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__buf_6
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4470__55/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2541 hold2541/A vssd1 vssd1 vccd1 vccd1 hold2541/X sky130_fd_sc_hd__buf_2
Xhold2574 hold2574/A vssd1 vssd1 vccd1 vccd1 hold2574/X sky130_fd_sc_hd__buf_2
XFILLER_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2552 hold2552/A vssd1 vssd1 vccd1 vccd1 hold512/A sky130_fd_sc_hd__buf_2
Xhold2563 hold2563/A vssd1 vssd1 vccd1 vccd1 hold2563/X sky130_fd_sc_hd__buf_2
XFILLER_48_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2585 hold2585/A vssd1 vssd1 vccd1 vccd1 hold2585/X sky130_fd_sc_hd__buf_2
Xhold2596 hold2596/A vssd1 vssd1 vccd1 vccd1 hold2596/X sky130_fd_sc_hd__buf_2
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1862 hold148/X vssd1 vssd1 vccd1 vccd1 hold1862/X sky130_fd_sc_hd__buf_2
Xhold1873 hold584/X vssd1 vssd1 vccd1 vccd1 hold1873/X sky130_fd_sc_hd__buf_2
XFILLER_72_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1884 hold867/X vssd1 vssd1 vccd1 vccd1 hold1884/X sky130_fd_sc_hd__buf_2
Xhold1895 hold841/X vssd1 vssd1 vccd1 vccd1 hold1895/X sky130_fd_sc_hd__buf_2
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4900__485 _4901__486/A vssd1 vssd1 vccd1 vccd1 _5621_/CLK sky130_fd_sc_hd__inv_2
XFILLER_138_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _5259_/Q _3654_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _3991_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2942_ _5429_/Q _5405_/Q _5397_/Q _5437_/Q _3069_/S _2942_/S1 vssd1 vssd1 vccd1 vccd1
+ _2942_/X sky130_fd_sc_hd__mux4_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5730_ _5730_/CLK _5730_/D vssd1 vssd1 vccd1 vccd1 _5730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2873_ _5367_/Q _2873_/B vssd1 vssd1 vccd1 vccd1 _2875_/B sky130_fd_sc_hd__nor2_1
X_5661_ _5661_/CLK _5661_/D vssd1 vssd1 vccd1 vccd1 _5661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5592_ _5592_/CLK _5592_/D vssd1 vssd1 vccd1 vccd1 _5592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold403 hold403/A vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__buf_2
Xhold425 hold502/X vssd1 vssd1 vccd1 vccd1 hold503/A sky130_fd_sc_hd__buf_2
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold458 hold458/A vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__buf_2
Xhold469 _4403_/X vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__buf_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3425_ _3526_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3433_/S sky130_fd_sc_hd__nor2_8
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _2464_/A _3357_/A _3355_/Y _4093_/B vssd1 vssd1 vccd1 vccd1 _5328_/D sky130_fd_sc_hd__o211a_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1114 hold2357/X vssd1 vssd1 vccd1 vccd1 hold2358/A sky130_fd_sc_hd__buf_2
X_3287_ _5576_/Q _5592_/Q _3318_/S vssd1 vssd1 vccd1 vccd1 _3287_/X sky130_fd_sc_hd__mux2_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5026_ _5026_/CLK _5026_/D vssd1 vssd1 vccd1 vccd1 _5026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1158 hold2231/X vssd1 vssd1 vccd1 vccd1 hold2232/A sky130_fd_sc_hd__buf_2
Xhold1125 hold2050/X vssd1 vssd1 vccd1 vccd1 hold2051/A sky130_fd_sc_hd__buf_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1169 hold2736/X vssd1 vssd1 vccd1 vccd1 hold1844/A sky130_fd_sc_hd__buf_2
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4843__428 _4468__53/A vssd1 vssd1 vccd1 vccd1 _5536_/CLK sky130_fd_sc_hd__inv_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5928_ _5928_/A vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5859_ _5859_/A vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__clkbuf_4
X_4737__322 _5005_/CLK vssd1 vssd1 vccd1 vccd1 _5428_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold981 hold981/A vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__buf_2
Xhold970 hold970/A vssd1 vssd1 vccd1 vccd1 hold970/X sky130_fd_sc_hd__buf_2
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold992 hold992/A vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__buf_2
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2382 hold909/X vssd1 vssd1 vccd1 vccd1 hold2382/X sky130_fd_sc_hd__buf_2
Xhold2371 hold2371/A vssd1 vssd1 vccd1 vccd1 hold2371/X sky130_fd_sc_hd__buf_2
Xhold2393 hold2393/A vssd1 vssd1 vccd1 vccd1 input136/A sky130_fd_sc_hd__buf_2
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1692 hold2339/X vssd1 vssd1 vccd1 vccd1 hold2340/A sky130_fd_sc_hd__buf_2
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4450__35 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5044_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4190_ _4204_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4190_/Y sky130_fd_sc_hd__nor2_1
X_3210_ _3208_/X _3209_/X _3240_/S vssd1 vssd1 vccd1 vccd1 _3210_/X sky130_fd_sc_hd__mux2_1
X_3141_ _5646_/Q _5638_/Q _5049_/Q _5654_/Q _3284_/S _3130_/B vssd1 vssd1 vccd1 vccd1
+ _3141_/X sky130_fd_sc_hd__mux4_1
X_4530__115 _4439__24/A vssd1 vssd1 vccd1 vccd1 _5172_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3072_ _5154_/Q _5310_/Q _3072_/S vssd1 vssd1 vccd1 vccd1 _3072_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3974_ _3639_/A _5244_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _5244_/D sky130_fd_sc_hd__mux2_1
X_2925_ _5127_/Q _5159_/Q _5315_/Q _5360_/Q _2941_/S0 _3072_/S vssd1 vssd1 vccd1 vccd1
+ _2925_/X sky130_fd_sc_hd__mux4_2
X_5713_ _5713_/CLK _5713_/D vssd1 vssd1 vccd1 vccd1 _5713_/Q sky130_fd_sc_hd__dfxtp_1
X_5644_ _5644_/CLK _5644_/D vssd1 vssd1 vccd1 vccd1 _5644_/Q sky130_fd_sc_hd__dfxtp_1
X_2856_ _5389_/Q _5696_/Q _2860_/S vssd1 vssd1 vccd1 vccd1 _5389_/D sky130_fd_sc_hd__mux2_1
X_2787_ _5449_/Q _3606_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5449_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__buf_2
Xhold211 hold226/X vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__buf_2
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5743_/CLK sky130_fd_sc_hd__clkbuf_8
X_5575_ _5575_/CLK _5575_/D vssd1 vssd1 vccd1 vccd1 _5575_/Q sky130_fd_sc_hd__dfxtp_1
XCaravelHost_651 vssd1 vssd1 vccd1 vccd1 CaravelHost_651/HI caravel_irq[0] sky130_fd_sc_hd__conb_1
XFILLER_144_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold233 _3991_/X vssd1 vssd1 vccd1 vccd1 _5259_/D sky130_fd_sc_hd__buf_2
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XCaravelHost_673 vssd1 vssd1 vccd1 vccd1 CaravelHost_673/HI la_data_out[101] sky130_fd_sc_hd__conb_1
Xhold222 hold236/X vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__buf_2
XCaravelHost_662 vssd1 vssd1 vccd1 vccd1 CaravelHost_662/HI core0Index[7] sky130_fd_sc_hd__conb_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__buf_2
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold255 hold270/X vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__buf_2
XCaravelHost_695 vssd1 vssd1 vccd1 vccd1 CaravelHost_695/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XCaravelHost_684 vssd1 vssd1 vccd1 vccd1 CaravelHost_684/HI la_data_out[112] sky130_fd_sc_hd__conb_1
Xhold288 _3809_/X vssd1 vssd1 vccd1 vccd1 _5009_/D sky130_fd_sc_hd__buf_2
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 _3930_/A sky130_fd_sc_hd__buf_2
X_3408_ _5272_/Q _3564_/A1 _3414_/S vssd1 vssd1 vccd1 vccd1 _5272_/D sky130_fd_sc_hd__mux2_1
X_4388_ _4389_/C _5743_/Q vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__and2b_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3339_/A1 _3159_/B _3338_/X _4093_/B vssd1 vssd1 vccd1 vccd1 _5337_/D sky130_fd_sc_hd__o211a_1
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _5010_/CLK _5009_/D vssd1 vssd1 vccd1 vccd1 _5009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4865__450 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5586_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4906__491 _5019_/CLK vssd1 vssd1 vccd1 vccd1 _5627_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2710_ _3395_/A0 _5514_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5514_/D sky130_fd_sc_hd__mux2_1
X_3690_ _4983_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3690_/X sky130_fd_sc_hd__or2_1
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2641_ _5602_/Q _3603_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5602_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5360_ _5360_/CLK _5360_/D vssd1 vssd1 vccd1 vccd1 _5360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2572_ _3577_/A0 _5641_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5641_/D sky130_fd_sc_hd__mux2_1
Xoutput316 _5885_/X vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_12
Xoutput305 _5875_/X vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_12
XFILLER_126_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5291_ _5291_/CLK hold35/X vssd1 vssd1 vccd1 vccd1 _5291_/Q sky130_fd_sc_hd__dfxtp_2
X_4311_ _4310_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _5675_/D sky130_fd_sc_hd__and2b_1
Xoutput349 _5915_/X vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_12
Xoutput338 _5905_/X vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_12
Xoutput327 _5895_/X vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_12
X_4242_ _5565_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__or2_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _5746_/Q _4157_/B _4118_/B vssd1 vssd1 vccd1 vccd1 _4173_/Y sky130_fd_sc_hd__a21boi_1
Xclkbuf_leaf_109_wb_clk_i _5743_/CLK vssd1 vssd1 vccd1 vccd1 _5546_/CLK sky130_fd_sc_hd__clkbuf_16
X_3124_ _4093_/C vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3055_ _5034_/Q _5531_/Q _3063_/S vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ _4368_/A _3957_/B vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__and2_1
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2908_ _3073_/C1 _2906_/X _3043_/A vssd1 vssd1 vccd1 vccd1 _2908_/X sky130_fd_sc_hd__a21o_1
X_3888_ _3888_/A _4399_/C _3888_/C vssd1 vssd1 vccd1 vccd1 _3888_/Y sky130_fd_sc_hd__nor3_1
X_2839_ _2848_/A1 _5404_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5404_/D sky130_fd_sc_hd__mux2_1
X_5627_ _5627_/CLK _5627_/D vssd1 vssd1 vccd1 vccd1 _5627_/Q sky130_fd_sc_hd__dfxtp_1
X_5558_ _5564_/CLK _5558_/D vssd1 vssd1 vccd1 vccd1 _5558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5489_ _5489_/CLK _5489_/D vssd1 vssd1 vccd1 vccd1 _5489_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout521 _3005_/S vssd1 vssd1 vccd1 vccd1 _3066_/S sky130_fd_sc_hd__buf_6
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout532 _3184_/S1 vssd1 vssd1 vccd1 vccd1 _3219_/S0 sky130_fd_sc_hd__clkbuf_16
Xfanout510 _2464_/Y vssd1 vssd1 vccd1 vccd1 _3331_/A2 sky130_fd_sc_hd__buf_8
X_4849__434 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5570_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout543 fanout547/X vssd1 vssd1 vccd1 vccd1 _3284_/S sky130_fd_sc_hd__clkbuf_16
Xfanout565 _5698_/Q vssd1 vssd1 vccd1 vccd1 _2790_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout554 _3797_/A3 vssd1 vssd1 vccd1 vccd1 _3796_/A3 sky130_fd_sc_hd__buf_4
Xfanout598 _2916_/A1 vssd1 vssd1 vccd1 vccd1 _3609_/A1 sky130_fd_sc_hd__buf_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout576 _3402_/A1 vssd1 vssd1 vccd1 vccd1 _3393_/A0 sky130_fd_sc_hd__buf_4
Xfanout587 _5693_/Q vssd1 vssd1 vccd1 vccd1 _3308_/A1 sky130_fd_sc_hd__buf_4
XFILLER_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_7_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5755_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3811_ _5262_/Q hold358/X _3814_/A3 _3814_/B1 _5011_/Q vssd1 vssd1 vccd1 vccd1 _3811_/X
+ sky130_fd_sc_hd__o32a_1
X_4642__227 _4921__506/A vssd1 vssd1 vccd1 vccd1 _5328_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_39 _5025_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 _4389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 _3389_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3742_ _3824_/A1 _3740_/X _3741_/X _3766_/C1 vssd1 vssd1 vccd1 vccd1 _3742_/X sky130_fd_sc_hd__o211a_4
XFILLER_146_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3673_ _3673_/A _3682_/B vssd1 vssd1 vccd1 vccd1 _3673_/X sky130_fd_sc_hd__and2_1
X_2624_ _3453_/C _5370_/Q _5369_/Q vssd1 vssd1 vccd1 vccd1 _3081_/A sky130_fd_sc_hd__nand3_2
X_5412_ _5412_/CLK _5412_/D vssd1 vssd1 vccd1 vccd1 _5412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _5343_/CLK _5343_/D vssd1 vssd1 vccd1 vccd1 _5343_/Q sky130_fd_sc_hd__dfxtp_1
X_4536__121 _4419__4/A vssd1 vssd1 vccd1 vccd1 _5178_/CLK sky130_fd_sc_hd__inv_2
X_2555_ _5655_/Q _3396_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _5655_/D sky130_fd_sc_hd__mux2_1
Xhold2904 hold2904/A vssd1 vssd1 vccd1 vccd1 hold2904/X sky130_fd_sc_hd__buf_2
X_5274_ _5274_/CLK _5274_/D vssd1 vssd1 vccd1 vccd1 _5274_/Q sky130_fd_sc_hd__dfxtp_1
X_2486_ _2486_/A _2486_/B vssd1 vssd1 vccd1 vccd1 _2487_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4225_ _4220_/B _4222_/X _5557_/Q vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__a21bo_1
X_4156_ _4108_/B _4119_/C _4108_/D _4122_/B _2456_/Y vssd1 vssd1 vccd1 vccd1 _4157_/B
+ sky130_fd_sc_hd__a32o_2
XFILLER_110_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3107_ _5359_/Q _3584_/A0 _3111_/S vssd1 vssd1 vccd1 vccd1 _5359_/D sky130_fd_sc_hd__mux2_1
X_4486__71 _5007_/CLK vssd1 vssd1 vccd1 vccd1 _5128_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _5688_/Q _4088_/B vssd1 vssd1 vccd1 vccd1 _4087_/X sky130_fd_sc_hd__and2_1
XFILLER_83_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3038_ _3099_/B _3036_/X _3037_/X vssd1 vssd1 vccd1 vccd1 _3038_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_77_wb_clk_i _4962__547/A vssd1 vssd1 vccd1 vccd1 _4456__41/A sky130_fd_sc_hd__clkbuf_16
X_4989_ _5022_/CLK _4989_/D vssd1 vssd1 vccd1 vccd1 _4989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _3771_/A sky130_fd_sc_hd__clkbuf_2
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
Xinput37 probe_out[10] vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput59 probe_out[30] vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__clkbuf_2
Xinput48 probe_out[20] vssd1 vssd1 vccd1 vccd1 _5857_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4010_ _4065_/B _4029_/C vssd1 vssd1 vccd1 vccd1 _4041_/B sky130_fd_sc_hd__nand2_1
XFILLER_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5892_ _5892_/A vssd1 vssd1 vccd1 vccd1 _5892_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3725_ _5078_/Q input6/X _3728_/S vssd1 vssd1 vccd1 vccd1 _3725_/X sky130_fd_sc_hd__mux2_4
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3656_ _3656_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__or2_1
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3587_ _3605_/A1 _5035_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5035_/D sky130_fd_sc_hd__mux2_1
X_2607_ _3573_/A0 _5613_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5613_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2538_ _3574_/A0 _5705_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5705_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5326_ _5326_/CLK _5326_/D vssd1 vssd1 vccd1 vccd1 _5326_/Q sky130_fd_sc_hd__dfxtp_2
X_4770__355 _4786__371/A vssd1 vssd1 vccd1 vccd1 _5461_/CLK sky130_fd_sc_hd__inv_2
X_5257_ _5259_/CLK _5257_/D vssd1 vssd1 vccd1 vccd1 _5257_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2712 _2467_/A vssd1 vssd1 vccd1 vccd1 _3789_/A1 sky130_fd_sc_hd__buf_2
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2756 _4391_/X vssd1 vssd1 vccd1 vccd1 hold2756/X sky130_fd_sc_hd__buf_2
X_2469_ _5346_/Q vssd1 vssd1 vccd1 vccd1 _3125_/A sky130_fd_sc_hd__clkinv_4
X_4208_ _4217_/A _4208_/B vssd1 vssd1 vccd1 vccd1 _5550_/D sky130_fd_sc_hd__nor2_1
X_5188_ _5188_/CLK _5188_/D vssd1 vssd1 vccd1 vccd1 _5188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2778 _3954_/Y vssd1 vssd1 vccd1 vccd1 hold2778/X sky130_fd_sc_hd__buf_2
X_4811__396 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5502_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2789 hold2888/X vssd1 vssd1 vccd1 vccd1 hold2789/X sky130_fd_sc_hd__buf_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4139_ _5755_/Q _5539_/Q vssd1 vssd1 vccd1 vccd1 _4139_/X sky130_fd_sc_hd__or2_1
XFILLER_73_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4705__290 _5256_/CLK vssd1 vssd1 vccd1 vccd1 _5396_/CLK sky130_fd_sc_hd__inv_2
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3510_ _3591_/A1 _5152_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5152_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3441_ _5219_/Q _3596_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5219_/D sky130_fd_sc_hd__mux2_1
X_4754__339 _4786__371/A vssd1 vssd1 vccd1 vccd1 _5445_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3372_ _3564_/A1 _5307_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5307_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5111_/CLK _5111_/D vssd1 vssd1 vccd1 vccd1 _5111_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/CLK _5042_/D vssd1 vssd1 vccd1 vccd1 _5042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4456__41 _4456__41/A vssd1 vssd1 vccd1 vccd1 _5050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4648__233 _5248_/CLK vssd1 vssd1 vccd1 vccd1 _5334_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5875_ _5875_/A vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3708_ _4989_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3708_/X sky130_fd_sc_hd__or2_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3639_ _3639_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3639_/X sky130_fd_sc_hd__or2_1
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5309_ _5735_/CLK _5309_/D vssd1 vssd1 vccd1 vccd1 _5309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput205 input205/A vssd1 vssd1 vccd1 vccd1 _3624_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2542 hold2542/A vssd1 vssd1 vccd1 vccd1 hold2542/X sky130_fd_sc_hd__buf_2
XFILLER_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2553 hold512/X vssd1 vssd1 vccd1 vccd1 hold2553/X sky130_fd_sc_hd__buf_2
Xhold2564 hold2564/A vssd1 vssd1 vccd1 vccd1 hold2564/X sky130_fd_sc_hd__buf_2
XFILLER_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2575 hold2575/A vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__buf_2
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2586 hold2586/A vssd1 vssd1 vccd1 vccd1 hold383/A sky130_fd_sc_hd__buf_2
Xhold1830 hold2739/X vssd1 vssd1 vccd1 vccd1 hold2740/A sky130_fd_sc_hd__buf_2
Xhold1863 hold1863/A vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__buf_2
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1874 hold1874/A vssd1 vssd1 vccd1 vccd1 _4380_/B1 sky130_fd_sc_hd__buf_2
Xhold1885 hold1885/A vssd1 vssd1 vccd1 vccd1 _4394_/B1 sky130_fd_sc_hd__buf_2
Xhold1896 hold1896/A vssd1 vssd1 vccd1 vccd1 _4387_/B1 sky130_fd_sc_hd__buf_2
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4901__486/A
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_21_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4477__62/A
+ sky130_fd_sc_hd__clkbuf_16
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3990_ _5258_/Q _3653_/A _3997_/S vssd1 vssd1 vccd1 vccd1 _5258_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2941_ _5126_/Q _5158_/Q _5314_/Q _5359_/Q _2941_/S0 _3072_/S vssd1 vssd1 vccd1 vccd1
+ _2941_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5660_ _5660_/CLK _5660_/D vssd1 vssd1 vccd1 vccd1 _5660_/Q sky130_fd_sc_hd__dfxtp_1
X_2872_ _5367_/Q _2873_/B vssd1 vssd1 vccd1 vccd1 _2883_/B sky130_fd_sc_hd__and2_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5591_ _5591_/CLK _5591_/D vssd1 vssd1 vccd1 vccd1 _5591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold404 hold404/A vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__buf_2
Xhold426 _4313_/X vssd1 vssd1 vccd1 vccd1 _5676_/D sky130_fd_sc_hd__buf_2
Xhold415 hold415/A vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__buf_2
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3424_ _3597_/A1 _5234_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5234_/D sky130_fd_sc_hd__mux2_1
Xhold459 hold459/A vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__buf_2
Xhold437 hold437/A vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__buf_2
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3357_/A _3355_/B vssd1 vssd1 vccd1 vccd1 _3355_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3325_/A _3284_/X _3285_/X _3320_/C1 vssd1 vssd1 vccd1 vccd1 _3286_/X sky130_fd_sc_hd__o211a_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5025_/CLK _5025_/D vssd1 vssd1 vccd1 vccd1 _5025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1126 hold2052/X vssd1 vssd1 vccd1 vccd1 hold2053/A sky130_fd_sc_hd__buf_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4882__467 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5603_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5927_ _5927_/A vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _5858_/A vssd1 vssd1 vccd1 vccd1 _5858_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4776__361 _4937__522/A vssd1 vssd1 vccd1 vccd1 _5467_/CLK sky130_fd_sc_hd__inv_2
XFILLER_135_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold971 hold971/A vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__buf_2
Xhold960 hold960/A vssd1 vssd1 vccd1 vccd1 hold960/X sky130_fd_sc_hd__buf_2
XFILLER_1_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold982 hold982/A vssd1 vssd1 vccd1 vccd1 hold982/X sky130_fd_sc_hd__buf_2
XFILLER_89_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold993 hold993/A vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__buf_2
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2372 hold2372/A vssd1 vssd1 vccd1 vccd1 _5692_/D sky130_fd_sc_hd__buf_2
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2383 hold2383/A vssd1 vssd1 vccd1 vccd1 hold2383/X sky130_fd_sc_hd__buf_2
Xhold2394 _3671_/A vssd1 vssd1 vccd1 vccd1 hold2394/X sky130_fd_sc_hd__buf_2
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1660 hold2309/X vssd1 vssd1 vccd1 vccd1 hold2310/A sky130_fd_sc_hd__buf_2
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1693 hold2341/X vssd1 vssd1 vccd1 vccd1 hold2342/A sky130_fd_sc_hd__buf_2
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3140_ _3140_/A _3140_/B vssd1 vssd1 vccd1 vccd1 _3140_/X sky130_fd_sc_hd__or2_2
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3071_ _3074_/A1 _3069_/X _3070_/X vssd1 vssd1 vccd1 vccd1 _3071_/Y sky130_fd_sc_hd__o21ai_1
X_4426__11 _4469__54/A vssd1 vssd1 vccd1 vccd1 _4977_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4610__195 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5284_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3973_ _3638_/A _5243_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _5243_/D sky130_fd_sc_hd__mux2_1
X_5712_ _5712_/CLK _5712_/D vssd1 vssd1 vccd1 vccd1 _5712_/Q sky130_fd_sc_hd__dfxtp_1
X_2924_ _2945_/A _2924_/B vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__and2_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2855_ _5390_/Q _3391_/A0 _2860_/S vssd1 vssd1 vccd1 vccd1 _5390_/D sky130_fd_sc_hd__mux2_1
X_5643_ _5643_/CLK _5643_/D vssd1 vssd1 vccd1 vccd1 _5643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5574_ _5574_/CLK _5574_/D vssd1 vssd1 vccd1 vccd1 _5574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2786_ _5450_/Q _2850_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5450_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XCaravelHost_652 vssd1 vssd1 vccd1 vccd1 CaravelHost_652/HI caravel_irq[1] sky130_fd_sc_hd__conb_1
Xhold212 hold230/X vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__buf_2
XCaravelHost_674 vssd1 vssd1 vccd1 vccd1 CaravelHost_674/HI la_data_out[102] sky130_fd_sc_hd__conb_1
Xhold234 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__buf_2
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__buf_2
XCaravelHost_663 vssd1 vssd1 vccd1 vccd1 CaravelHost_663/HI core1Index[1] sky130_fd_sc_hd__conb_1
XFILLER_144_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold278 _3807_/X vssd1 vssd1 vccd1 vccd1 _5007_/D sky130_fd_sc_hd__buf_2
Xhold267 hold354/X vssd1 vssd1 vccd1 vccd1 hold355/A sky130_fd_sc_hd__buf_2
Xhold245 hold273/X vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__buf_2
Xhold256 hold272/X vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__buf_2
XCaravelHost_696 vssd1 vssd1 vccd1 vccd1 CaravelHost_696/HI la_data_out[124] sky130_fd_sc_hd__conb_1
XCaravelHost_685 vssd1 vssd1 vccd1 vccd1 CaravelHost_685/HI la_data_out[113] sky130_fd_sc_hd__conb_1
XFILLER_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3407_ _5273_/Q _3572_/A0 _3414_/S vssd1 vssd1 vccd1 vccd1 _5273_/D sky130_fd_sc_hd__mux2_1
X_4387_ _5742_/Q _4389_/C _4387_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4387_/X sky130_fd_sc_hd__o211a_1
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _5337_/Q _3125_/A _3156_/X _3337_/X vssd1 vssd1 vccd1 vccd1 _3338_/X sky130_fd_sc_hd__a211o_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3269_ _5475_/Q _3331_/A2 _3237_/B _5710_/Q vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__o22a_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ _5010_/CLK _5008_/D vssd1 vssd1 vccd1 vccd1 _5008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4553__138 _4418__3/A vssd1 vssd1 vccd1 vccd1 _5195_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2191 hold2803/X vssd1 vssd1 vccd1 vccd1 hold2804/A sky130_fd_sc_hd__buf_2
X_4510__95 _4510__95/A vssd1 vssd1 vccd1 vccd1 _5152_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1490 hold2260/X vssd1 vssd1 vccd1 vccd1 hold2261/A sky130_fd_sc_hd__buf_2
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2640_ _5603_/Q _3611_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5603_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput306 _5876_/X vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_12
X_2571_ _3576_/A0 _5642_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5642_/D sky130_fd_sc_hd__mux2_1
Xoutput317 _5886_/X vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_12
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4310_ _4248_/B _4318_/A2 _4322_/B _2443_/Y vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__o22a_1
X_5290_ _5733_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _5290_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput339 _5906_/X vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_12
Xoutput328 _5896_/X vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_12
X_4241_ _5343_/Q _3124_/Y _4164_/B _4240_/X hold741/X vssd1 vssd1 vccd1 vccd1 _4241_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ _5750_/Q _4130_/Y _4145_/A _4145_/C _4148_/B vssd1 vssd1 vccd1 vccd1 _4172_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_95_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3123_ _3123_/A _3123_/B _3123_/C _3122_/X vssd1 vssd1 vccd1 vccd1 _4093_/C sky130_fd_sc_hd__or4b_2
X_3054_ _3099_/B _3052_/X _3053_/X vssd1 vssd1 vccd1 vccd1 _3054_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3956_ _3930_/A split1/X _3778_/C _3897_/C vssd1 vssd1 vccd1 vccd1 _3956_/X sky130_fd_sc_hd__a31o_1
X_2907_ _5064_/Q _5040_/Q _5537_/Q _4981_/Q _2941_/S0 _3024_/S vssd1 vssd1 vccd1 vccd1
+ _2907_/X sky130_fd_sc_hd__mux4_1
X_3887_ _3887_/A _3887_/B vssd1 vssd1 vccd1 vccd1 _3887_/X sky130_fd_sc_hd__and2_2
X_5626_ _5626_/CLK _5626_/D vssd1 vssd1 vccd1 vccd1 _5626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2838_ _3584_/A0 _5405_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5405_/D sky130_fd_sc_hd__mux2_1
X_5557_ _5557_/CLK _5557_/D vssd1 vssd1 vccd1 vccd1 _5557_/Q sky130_fd_sc_hd__dfxtp_1
X_2769_ _2790_/A0 _5463_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5463_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5488_ _5488_/CLK _5488_/D vssd1 vssd1 vccd1 vccd1 _5488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout500 _3031_/B1 vssd1 vssd1 vccd1 vccd1 _3073_/B2 sky130_fd_sc_hd__buf_6
XFILLER_120_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout522 _3005_/S vssd1 vssd1 vccd1 vccd1 _3063_/S sky130_fd_sc_hd__buf_6
Xfanout511 _5372_/Q vssd1 vssd1 vccd1 vccd1 _3443_/B sky130_fd_sc_hd__buf_6
Xfanout533 _3126_/A vssd1 vssd1 vccd1 vccd1 _3184_/S1 sky130_fd_sc_hd__buf_4
XFILLER_113_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout555 _3797_/A3 vssd1 vssd1 vccd1 vccd1 _3810_/A3 sky130_fd_sc_hd__buf_6
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout566 _5698_/Q vssd1 vssd1 vccd1 vccd1 _3573_/A0 sky130_fd_sc_hd__buf_6
Xfanout544 fanout547/X vssd1 vssd1 vccd1 vccd1 _3318_/S sky130_fd_sc_hd__buf_4
X_4888__473 _4921__506/A vssd1 vssd1 vccd1 vccd1 _5609_/CLK sky130_fd_sc_hd__inv_2
Xfanout599 _2916_/A1 vssd1 vssd1 vccd1 vccd1 _3600_/A1 sky130_fd_sc_hd__clkbuf_8
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout588 _5692_/Q vssd1 vssd1 vccd1 vccd1 _3396_/A0 sky130_fd_sc_hd__buf_4
Xfanout577 _3567_/A1 vssd1 vssd1 vccd1 vccd1 _3576_/A0 sky130_fd_sc_hd__buf_4
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _5261_/Q hold358/X _3810_/A3 hold349/X _5010_/Q vssd1 vssd1 vccd1 vccd1 _3810_/X
+ sky130_fd_sc_hd__o32a_1
X_4681__266 _5383_/CLK vssd1 vssd1 vccd1 vccd1 _5370_/CLK sky130_fd_sc_hd__inv_2
X_3741_ _5000_/Q _3750_/B vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__or2_1
XANTENNA_18 _4389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 _3396_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3672_ _3672_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__and2_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2623_ _5370_/Q _5369_/Q vssd1 vssd1 vccd1 vccd1 _2777_/A sky130_fd_sc_hd__nand2_2
X_5411_ _5411_/CLK _5411_/D vssd1 vssd1 vccd1 vccd1 _5411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5342_ _5342_/CLK _5342_/D vssd1 vssd1 vccd1 vccd1 _5342_/Q sky130_fd_sc_hd__dfxtp_1
X_2554_ _5656_/Q _3395_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _5656_/D sky130_fd_sc_hd__mux2_1
X_4575__160 _4438__23/A vssd1 vssd1 vccd1 vccd1 _5225_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _5273_/CLK _5273_/D vssd1 vssd1 vccd1 vccd1 _5273_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2905 hold2905/A vssd1 vssd1 vccd1 vccd1 hold2905/X sky130_fd_sc_hd__buf_2
X_2485_ _2545_/A _3123_/C _3123_/B vssd1 vssd1 vccd1 vccd1 _2486_/B sky130_fd_sc_hd__a21oi_1
XFILLER_96_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4224_ _2454_/Y _4221_/C _4223_/X vssd1 vssd1 vccd1 vccd1 _5556_/D sky130_fd_sc_hd__a21oi_1
X_4155_ _5742_/Q _4155_/B vssd1 vssd1 vccd1 vccd1 _4170_/B sky130_fd_sc_hd__xor2_1
XFILLER_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3106_ _5360_/Q _3538_/A0 _3111_/S vssd1 vssd1 vccd1 vccd1 _5360_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4086_ _5687_/Q _4088_/B vssd1 vssd1 vccd1 vccd1 _4086_/X sky130_fd_sc_hd__and2_1
XFILLER_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3037_ _2867_/A _5187_/Q _2866_/B _5195_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3037_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4922__507 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5643_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4988_ _5022_/CLK _4988_/D vssd1 vssd1 vccd1 vccd1 _4988_/Q sky130_fd_sc_hd__dfxtp_1
X_3939_ _3939_/A0 _5096_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_wb_clk_i clkbuf_4_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4816__401 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5507_/CLK sky130_fd_sc_hd__inv_2
X_5609_ _5609_/CLK _5609_/D vssd1 vssd1 vccd1 vccd1 _5609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__clkbuf_2
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _3752_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput49 probe_out[21] vssd1 vssd1 vccd1 vccd1 _5858_/A sky130_fd_sc_hd__clkbuf_2
Xinput38 probe_out[11] vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__clkbuf_2
X_4559__144 _4423__8/A vssd1 vssd1 vccd1 vccd1 _5201_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _5891_/A vssd1 vssd1 vccd1 vccd1 _5891_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _3733_/A1 _3722_/X _3723_/X split2/A vssd1 vssd1 vccd1 vccd1 _3724_/X sky130_fd_sc_hd__o211a_1
XFILLER_146_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3655_ _3655_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3655_/X sky130_fd_sc_hd__or2_1
XFILLER_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2606_ _3159_/A _5614_/Q _2613_/S vssd1 vssd1 vccd1 vccd1 _5614_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3586_ _3604_/A1 _5036_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5036_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5325_ _5691_/CLK _5325_/D vssd1 vssd1 vccd1 vccd1 _5325_/Q sky130_fd_sc_hd__dfxtp_1
X_2537_ _3564_/A1 _5706_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5706_/D sky130_fd_sc_hd__mux2_1
X_5256_ _5256_/CLK _5256_/D vssd1 vssd1 vccd1 vccd1 _5256_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2468_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__inv_2
Xhold2713 _3787_/X vssd1 vssd1 vccd1 vccd1 hold2713/X sky130_fd_sc_hd__buf_2
Xhold2735 _4377_/X vssd1 vssd1 vccd1 vccd1 hold2735/X sky130_fd_sc_hd__buf_2
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4207_ _5550_/Q _4209_/B _4186_/X _4110_/B vssd1 vssd1 vccd1 vccd1 _4208_/B sky130_fd_sc_hd__o2bb2a_1
X_5187_ _5187_/CLK _5187_/D vssd1 vssd1 vccd1 vccd1 _5187_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2768 _4375_/X vssd1 vssd1 vccd1 vccd1 hold2768/X sky130_fd_sc_hd__buf_2
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4138_ _5755_/Q _5539_/Q vssd1 vssd1 vccd1 vccd1 _4138_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4069_ _4071_/B _4071_/C vssd1 vssd1 vccd1 vccd1 _4248_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4793__378 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5484_/CLK sky130_fd_sc_hd__inv_2
XFILLER_143_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3440_ _5220_/Q _3595_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5220_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3371_ _3572_/A0 _5308_/Q _3378_/S vssd1 vssd1 vccd1 vccd1 _5308_/D sky130_fd_sc_hd__mux2_1
X_5110_ _5256_/CLK _5110_/D vssd1 vssd1 vccd1 vccd1 _5110_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/CLK _5041_/D vssd1 vssd1 vccd1 vccd1 _5041_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4687__272 _5384_/CLK vssd1 vssd1 vccd1 vccd1 _5376_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4471__56 _5002_/CLK vssd1 vssd1 vccd1 vccd1 _5065_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5874_ _5874_/A vssd1 vssd1 vccd1 vccd1 _5874_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3707_ _5072_/Q input31/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__mux2_4
X_3638_ _3638_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__or2_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3569_ _5051_/Q _3569_/A1 _3570_/S vssd1 vssd1 vccd1 vccd1 _5051_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5308_ _5308_/CLK _5308_/D vssd1 vssd1 vccd1 vccd1 _5308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2510 hold2856/X vssd1 vssd1 vccd1 vccd1 hold2510/X sky130_fd_sc_hd__buf_2
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2543 hold2543/A vssd1 vssd1 vccd1 vccd1 _5321_/D sky130_fd_sc_hd__buf_2
X_5239_ _5239_/CLK _5239_/D vssd1 vssd1 vccd1 vccd1 _5239_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1820 hold2730/X vssd1 vssd1 vccd1 vccd1 hold2731/A sky130_fd_sc_hd__buf_2
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2565 hold2565/A vssd1 vssd1 vccd1 vccd1 hold548/A sky130_fd_sc_hd__buf_2
Xhold2554 hold2554/A vssd1 vssd1 vccd1 vccd1 hold2554/X sky130_fd_sc_hd__buf_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4928__513 _4455__40/A vssd1 vssd1 vccd1 vccd1 _5649_/CLK sky130_fd_sc_hd__inv_2
Xhold2576 hold203/X vssd1 vssd1 vccd1 vccd1 hold2576/X sky130_fd_sc_hd__buf_2
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2587 hold383/X vssd1 vssd1 vccd1 vccd1 hold2587/X sky130_fd_sc_hd__buf_2
Xhold1831 hold1831/A vssd1 vssd1 vccd1 vccd1 _3825_/A2 sky130_fd_sc_hd__buf_2
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1875 _4380_/X vssd1 vssd1 vccd1 vccd1 hold1875/X sky130_fd_sc_hd__buf_2
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1886 _4394_/X vssd1 vssd1 vccd1 vccd1 hold1886/X sky130_fd_sc_hd__buf_2
Xhold1864 _3830_/X vssd1 vssd1 vccd1 vccd1 hold1864/X sky130_fd_sc_hd__buf_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1897 _4387_/X vssd1 vssd1 vccd1 vccd1 hold1897/X sky130_fd_sc_hd__buf_2
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _5261_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2940_ _5062_/Q _5038_/Q _5535_/Q _4979_/Q _2867_/B _3063_/S vssd1 vssd1 vccd1 vccd1
+ _2940_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4721__306 _5244_/CLK vssd1 vssd1 vccd1 vccd1 _5412_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2871_ _5145_/Q _5153_/Q _5217_/Q _5137_/Q _3036_/S _2944_/S0 vssd1 vssd1 vccd1 vccd1
+ _2871_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5590_ _5590_/CLK _5590_/D vssd1 vssd1 vccd1 vccd1 _5590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 _3970_/B vssd1 vssd1 vccd1 vccd1 _5363_/D sky130_fd_sc_hd__buf_2
Xhold416 hold416/A vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__buf_2
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3423_ _3596_/A1 _5235_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5235_/D sky130_fd_sc_hd__mux2_1
Xhold449 hold449/A vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__buf_2
X_4615__200 _4909__494/A vssd1 vssd1 vccd1 vccd1 _5289_/CLK sky130_fd_sc_hd__inv_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _5329_/Q _3353_/A _3353_/Y _4093_/B vssd1 vssd1 vccd1 vccd1 _5329_/D sky130_fd_sc_hd__o211a_1
XFILLER_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3285_ _5648_/Q _3331_/A2 _3326_/B2 _5640_/Q vssd1 vssd1 vccd1 vccd1 _3285_/X sky130_fd_sc_hd__o22a_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5024_ _5024_/CLK _5024_/D vssd1 vssd1 vccd1 vccd1 _5024_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5926_ _5926_/A vssd1 vssd1 vccd1 vccd1 _5926_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5857_ _5857_/A vssd1 vssd1 vccd1 vccd1 _5857_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold972 hold972/A vssd1 vssd1 vccd1 vccd1 hold972/X sky130_fd_sc_hd__buf_2
Xhold961 hold961/A vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__buf_2
XFILLER_135_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold983 hold983/A vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__buf_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold994 hold994/A vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__buf_2
XFILLER_135_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2340 hold2340/A vssd1 vssd1 vccd1 vccd1 hold2340/X sky130_fd_sc_hd__buf_2
XFILLER_103_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1650 hold206/X vssd1 vssd1 vccd1 vccd1 hold1650/X sky130_fd_sc_hd__buf_2
Xhold2384 hold2384/A vssd1 vssd1 vccd1 vccd1 hold2384/X sky130_fd_sc_hd__buf_2
Xhold2395 hold2395/A vssd1 vssd1 vccd1 vccd1 hold987/A sky130_fd_sc_hd__buf_2
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1683 hold2820/X vssd1 vssd1 vccd1 vccd1 hold2821/A sky130_fd_sc_hd__buf_2
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1694 hold2343/X vssd1 vssd1 vccd1 vccd1 hold2344/A sky130_fd_sc_hd__buf_2
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3070_ _5433_/Q _2460_/Y _3073_/B2 _5425_/Q _3097_/B vssd1 vssd1 vccd1 vccd1 _3070_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4441__26 _5001_/CLK vssd1 vssd1 vccd1 vccd1 _5035_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3972_ _3637_/A _5242_/Q _3979_/S vssd1 vssd1 vccd1 vccd1 _5242_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5711_ _5711_/CLK _5711_/D vssd1 vssd1 vccd1 vccd1 _5711_/Q sky130_fd_sc_hd__dfxtp_1
X_2923_ _5031_/Q _5175_/Q _5239_/Q _5223_/Q _2944_/S0 _3040_/S vssd1 vssd1 vccd1 vccd1
+ _2924_/B sky130_fd_sc_hd__mux4_2
XFILLER_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2854_ _5391_/Q _3390_/A0 _2860_/S vssd1 vssd1 vccd1 vccd1 _5391_/D sky130_fd_sc_hd__mux2_1
X_4799__384 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5490_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5642_ _5642_/CLK _5642_/D vssd1 vssd1 vccd1 vccd1 _5642_/Q sky130_fd_sc_hd__dfxtp_1
X_5573_ _5573_/CLK _5573_/D vssd1 vssd1 vccd1 vccd1 _5573_/Q sky130_fd_sc_hd__dfxtp_1
X_2785_ _5451_/Q _2849_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5451_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__buf_2
XCaravelHost_653 vssd1 vssd1 vccd1 vccd1 CaravelHost_653/HI caravel_irq[2] sky130_fd_sc_hd__conb_1
XFILLER_144_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold213 _3992_/X vssd1 vssd1 vccd1 vccd1 _5260_/D sky130_fd_sc_hd__buf_2
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__buf_2
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__buf_2
XCaravelHost_664 vssd1 vssd1 vccd1 vccd1 CaravelHost_664/HI core1Index[2] sky130_fd_sc_hd__conb_1
XFILLER_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold246 _3806_/X vssd1 vssd1 vccd1 vccd1 _5006_/D sky130_fd_sc_hd__buf_2
Xhold268 _3810_/X vssd1 vssd1 vccd1 vccd1 _5010_/D sky130_fd_sc_hd__buf_2
Xhold257 hold274/X vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__buf_2
XCaravelHost_697 vssd1 vssd1 vccd1 vccd1 CaravelHost_697/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XCaravelHost_686 vssd1 vssd1 vccd1 vccd1 CaravelHost_686/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XCaravelHost_675 vssd1 vssd1 vccd1 vccd1 CaravelHost_675/HI la_data_out[103] sky130_fd_sc_hd__conb_1
XFILLER_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4386_ _3642_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4386_/X sky130_fd_sc_hd__a21bo_1
X_3406_ _3406_/A _3571_/A vssd1 vssd1 vccd1 vccd1 _3414_/S sky130_fd_sc_hd__nor2_8
XFILLER_140_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _3334_/X _3336_/X _3357_/A vssd1 vssd1 vccd1 vccd1 _3337_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _5443_/Q _5459_/Q _3299_/S vssd1 vssd1 vccd1 vccd1 _3268_/X sky130_fd_sc_hd__mux2_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5007_/CLK _5007_/D vssd1 vssd1 vccd1 vccd1 _5007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3199_ _3574_/A0 _3159_/B _3198_/X _3277_/C1 vssd1 vssd1 vccd1 vccd1 _5342_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5909_ _5909_/A vssd1 vssd1 vccd1 vccd1 _5909_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4592__177 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5266_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2192 hold2805/X vssd1 vssd1 vccd1 vccd1 hold2806/A sky130_fd_sc_hd__buf_2
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1480 hold2253/X vssd1 vssd1 vccd1 vccd1 hold2254/A sky130_fd_sc_hd__buf_2
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1491 hold2262/X vssd1 vssd1 vccd1 vccd1 hold2263/A sky130_fd_sc_hd__buf_2
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4833__418 _4456__41/A vssd1 vssd1 vccd1 vccd1 _5524_/CLK sky130_fd_sc_hd__inv_2
Xoutput307 _5840_/X vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_12
X_2570_ _3575_/A0 _5643_/Q _2574_/S vssd1 vssd1 vccd1 vccd1 _5643_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput329 _5842_/X vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_12
Xoutput318 _5841_/X vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_12
XFILLER_141_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4240_ _5564_/Q _4242_/B vssd1 vssd1 vccd1 vccd1 _4240_/X sky130_fd_sc_hd__or2_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4171_ _4171_/A _4171_/B _4171_/C vssd1 vssd1 vccd1 vccd1 _4171_/X sky130_fd_sc_hd__and3_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3122_ _3122_/A _3122_/B _3122_/C vssd1 vssd1 vccd1 vccd1 _3122_/X sky130_fd_sc_hd__and3_1
X_3053_ _2460_/A _5130_/Q _2866_/B _5138_/Q _3064_/C1 vssd1 vssd1 vccd1 vccd1 _3053_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4727__312 _4941__526/A vssd1 vssd1 vccd1 vccd1 _5418_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ _3955_/A _3959_/C vssd1 vssd1 vccd1 vccd1 _3955_/Y sky130_fd_sc_hd__nor2_1
X_2906_ _5589_/Q _5573_/Q _5455_/Q _5605_/Q _3024_/S _2941_/S0 vssd1 vssd1 vccd1 vccd1
+ _2906_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3886_ _4401_/A _5208_/Q _3897_/C _3855_/X vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__a31o_1
X_5625_ _5625_/CLK _5625_/D vssd1 vssd1 vccd1 vccd1 _5625_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_118_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4956__541/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2837_ _3538_/A0 _5406_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5406_/D sky130_fd_sc_hd__mux2_1
X_5556_ _5557_/CLK _5556_/D vssd1 vssd1 vccd1 vccd1 _5556_/Q sky130_fd_sc_hd__dfxtp_2
X_2768_ _3389_/A0 _5464_/Q _2775_/S vssd1 vssd1 vccd1 vccd1 _5464_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2699_ _5524_/Q _3402_/A1 _2702_/S vssd1 vssd1 vccd1 vccd1 _5524_/D sky130_fd_sc_hd__mux2_1
X_5487_ _5487_/CLK _5487_/D vssd1 vssd1 vccd1 vccd1 _5487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout501 _2865_/X vssd1 vssd1 vccd1 vccd1 _3031_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout523 _3005_/S vssd1 vssd1 vccd1 vccd1 _3036_/S sky130_fd_sc_hd__clkbuf_16
Xfanout512 _5371_/Q vssd1 vssd1 vccd1 vccd1 _3453_/C sky130_fd_sc_hd__buf_12
Xfanout556 _3797_/A3 vssd1 vssd1 vccd1 vccd1 _3814_/A3 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4369_ _4369_/A _4399_/C _4369_/C _4369_/D vssd1 vssd1 vccd1 vccd1 _4401_/B sky130_fd_sc_hd__nor4_2
Xfanout545 fanout547/X vssd1 vssd1 vccd1 vccd1 _3324_/S sky130_fd_sc_hd__buf_8
Xfanout534 _3126_/A vssd1 vssd1 vccd1 vccd1 _3130_/B sky130_fd_sc_hd__buf_8
XFILLER_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout567 _5698_/Q vssd1 vssd1 vccd1 vccd1 _3564_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout589 _3387_/A1 vssd1 vssd1 vccd1 vccd1 _3579_/A0 sky130_fd_sc_hd__buf_4
Xfanout578 _3402_/A1 vssd1 vssd1 vccd1 vccd1 _3567_/A1 sky130_fd_sc_hd__buf_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4520__105 _4432__17/A vssd1 vssd1 vccd1 vccd1 _5162_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 _3657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3740_ _5083_/Q input11/X _3763_/B vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3671_ _3671_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3671_/X sky130_fd_sc_hd__and2_1
X_2622_ _5373_/Q _5368_/Q vssd1 vssd1 vccd1 vccd1 _2862_/B sky130_fd_sc_hd__xnor2_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5410_ _5410_/CLK _5410_/D vssd1 vssd1 vccd1 vccd1 _5410_/Q sky130_fd_sc_hd__dfxtp_1
X_5341_ _5341_/CLK _5341_/D vssd1 vssd1 vccd1 vccd1 _5341_/Q sky130_fd_sc_hd__dfxtp_1
X_2553_ _5657_/Q _3394_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _5657_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5272_ _5272_/CLK _5272_/D vssd1 vssd1 vccd1 vccd1 _5272_/Q sky130_fd_sc_hd__dfxtp_1
X_2484_ _2545_/A _3123_/C _2483_/X vssd1 vssd1 vccd1 vccd1 _2487_/C sky130_fd_sc_hd__o21ai_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4223_ _4220_/B _4222_/X _4217_/A vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__a21o_1
Xhold2906 hold2906/A vssd1 vssd1 vccd1 vccd1 hold2906/X sky130_fd_sc_hd__buf_2
X_4154_ _5552_/Q _4210_/A vssd1 vssd1 vccd1 vccd1 _4155_/B sky130_fd_sc_hd__xnor2_2
X_3105_ _5361_/Q _3600_/A1 _3111_/S vssd1 vssd1 vccd1 vccd1 _5361_/D sky130_fd_sc_hd__mux2_1
X_4085_ _5686_/Q _4088_/B vssd1 vssd1 vccd1 vccd1 _4085_/X sky130_fd_sc_hd__and2_1
XFILLER_83_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3036_ _4968_/Q _5179_/Q _3036_/S vssd1 vssd1 vccd1 vccd1 _3036_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4961__546 _4961__546/A vssd1 vssd1 vccd1 vccd1 _5719_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4987_ _5019_/CLK _4987_/D vssd1 vssd1 vccd1 vccd1 _4987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3938_ _3938_/A0 _5095_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3938_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3869_ _4399_/B _3866_/X _3868_/X _4361_/A vssd1 vssd1 vccd1 vccd1 _3869_/X sky130_fd_sc_hd__a31o_1
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855__440 _4892__477/A vssd1 vssd1 vccd1 vccd1 _5576_/CLK sky130_fd_sc_hd__inv_2
X_5608_ _5608_/CLK _5608_/D vssd1 vssd1 vccd1 vccd1 _5608_/Q sky130_fd_sc_hd__dfxtp_1
X_5539_ _5566_/CLK _5539_/D vssd1 vssd1 vccd1 vccd1 _5539_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4451__36/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i _4676__261/A vssd1 vssd1 vccd1 vccd1 _4435__20/A sky130_fd_sc_hd__clkbuf_16
XFILLER_87_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4477__62 _4477__62/A vssd1 vssd1 vccd1 vccd1 _5119_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__clkbuf_2
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
Xinput39 probe_out[12] vssd1 vssd1 vccd1 vccd1 _5849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4598__183 _4964__549/A vssd1 vssd1 vccd1 vccd1 _5272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5890_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5890_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4839__424 _5001_/CLK vssd1 vssd1 vccd1 vccd1 _5532_/CLK sky130_fd_sc_hd__inv_2
X_3723_ _4994_/Q _3729_/B vssd1 vssd1 vccd1 vccd1 _3723_/X sky130_fd_sc_hd__or2_1
X_3654_ _3654_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__or2_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2605_ _3562_/A _2664_/B vssd1 vssd1 vccd1 vccd1 _2613_/S sky130_fd_sc_hd__or2_4
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3585_ _3603_/A1 _5037_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5037_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5324_ _5691_/CLK _5324_/D vssd1 vssd1 vccd1 vccd1 _5324_/Q sky130_fd_sc_hd__dfxtp_1
X_2536_ _3572_/A0 _5707_/Q _2543_/S vssd1 vssd1 vccd1 vccd1 _5707_/D sky130_fd_sc_hd__mux2_1
X_5255_ _5256_/CLK _5255_/D vssd1 vssd1 vccd1 vccd1 _5255_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2467_ _2467_/A vssd1 vssd1 vccd1 vccd1 _2467_/Y sky130_fd_sc_hd__inv_4
Xhold2714 hold2714/A vssd1 vssd1 vccd1 vccd1 hold2714/X sky130_fd_sc_hd__buf_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2736 hold2736/A vssd1 vssd1 vccd1 vccd1 hold2736/X sky130_fd_sc_hd__buf_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4206_ _4217_/A _4206_/B vssd1 vssd1 vccd1 vccd1 _5549_/D sky130_fd_sc_hd__nor2_1
X_5186_ _5186_/CLK _5186_/D vssd1 vssd1 vccd1 vccd1 _5186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _5754_/Q _4137_/B vssd1 vssd1 vccd1 vccd1 _4137_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ _4021_/B _4021_/C _4029_/C _5675_/Q vssd1 vssd1 vccd1 vccd1 _4071_/C sky130_fd_sc_hd__a31o_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3019_ _2867_/A _5131_/Q _3041_/A2 _5139_/Q _2947_/S vssd1 vssd1 vccd1 vccd1 _3019_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4632__217 _5084_/CLK vssd1 vssd1 vccd1 vccd1 _5310_/CLK sky130_fd_sc_hd__inv_2
XFILLER_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4526__111 _4510__95/A vssd1 vssd1 vccd1 vccd1 _5168_/CLK sky130_fd_sc_hd__inv_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3370_ _3370_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3378_/S sky130_fd_sc_hd__or2_4
XFILLER_112_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/CLK _5040_/D vssd1 vssd1 vccd1 vccd1 _5040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5873_ _5873_/A vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3706_ _3718_/A1 _3704_/X _3705_/X split4/X vssd1 vssd1 vccd1 vccd1 _3706_/X sky130_fd_sc_hd__o211a_1
XFILLER_147_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3637_ _3637_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3637_/X sky130_fd_sc_hd__or2_1
X_3568_ _5052_/Q _3568_/A1 _3570_/S vssd1 vssd1 vccd1 vccd1 _5052_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5307_ _5307_/CLK _5307_/D vssd1 vssd1 vccd1 vccd1 _5307_/Q sky130_fd_sc_hd__dfxtp_1
X_2519_ _3566_/A1 _5720_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5720_/D sky130_fd_sc_hd__mux2_1
X_3499_ _3607_/A _3535_/B vssd1 vssd1 vccd1 vccd1 _3507_/S sky130_fd_sc_hd__nor2_8
XFILLER_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2500 hold2500/A vssd1 vssd1 vccd1 vccd1 hold799/A sky130_fd_sc_hd__buf_2
XFILLER_88_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2511 hold2511/A vssd1 vssd1 vccd1 vccd1 hold2511/X sky130_fd_sc_hd__buf_2
Xhold1810 hold2542/X vssd1 vssd1 vccd1 vccd1 hold2543/A sky130_fd_sc_hd__buf_2
X_5238_ _5238_/CLK _5238_/D vssd1 vssd1 vccd1 vccd1 _5238_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2555 hold2555/A vssd1 vssd1 vccd1 vccd1 hold2555/X sky130_fd_sc_hd__buf_2
XFILLER_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5169_ _5169_/CLK _5169_/D vssd1 vssd1 vccd1 vccd1 _5169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1843 hold2735/X vssd1 vssd1 vccd1 vccd1 hold2736/A sky130_fd_sc_hd__buf_2
Xhold2577 hold2577/A vssd1 vssd1 vccd1 vccd1 hold2577/X sky130_fd_sc_hd__buf_2
Xhold1821 hold1821/A vssd1 vssd1 vccd1 vccd1 hold727/A sky130_fd_sc_hd__buf_2
Xhold2588 hold2588/A vssd1 vssd1 vccd1 vccd1 hold2588/X sky130_fd_sc_hd__buf_2
Xhold1854 hold2583/X vssd1 vssd1 vccd1 vccd1 hold2584/A sky130_fd_sc_hd__buf_2
Xhold2566 hold548/X vssd1 vssd1 vccd1 vccd1 hold2566/X sky130_fd_sc_hd__buf_2
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1832 _3825_/X vssd1 vssd1 vccd1 vccd1 hold1832/X sky130_fd_sc_hd__buf_2
X_4447__32 _5002_/CLK vssd1 vssd1 vccd1 vccd1 _5041_/CLK sky130_fd_sc_hd__inv_2
Xhold1876 hold1876/A vssd1 vssd1 vccd1 vccd1 hold585/A sky130_fd_sc_hd__buf_2
Xhold1887 hold1887/A vssd1 vssd1 vccd1 vccd1 hold868/A sky130_fd_sc_hd__buf_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1865 hold1865/A vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__buf_2
XFILLER_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1898 hold1898/A vssd1 vssd1 vccd1 vccd1 hold842/A sky130_fd_sc_hd__buf_2
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4423__8/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__buf_2
XFILLER_75_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4760__345 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5451_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _2873_/B _2870_/B vssd1 vssd1 vccd1 vccd1 _2870_/X sky130_fd_sc_hd__or2_1
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4801__386 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5492_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3422_ _3595_/A1 _5236_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5236_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3353_/A _3353_/B vssd1 vssd1 vccd1 vccd1 _3353_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1106 hold2340/X vssd1 vssd1 vccd1 vccd1 hold2341/A sky130_fd_sc_hd__buf_2
X_3284_ _5043_/Q _5632_/Q _3284_/S vssd1 vssd1 vccd1 vccd1 _3284_/X sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5023_ _5024_/CLK _5023_/D vssd1 vssd1 vccd1 vccd1 _5023_/Q sky130_fd_sc_hd__dfxtp_2
Xhold1139 hold2402/X vssd1 vssd1 vccd1 vccd1 hold2403/A sky130_fd_sc_hd__buf_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5925_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5856_ _5856_/A vssd1 vssd1 vccd1 vccd1 _5856_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2999_ _5395_/Q _5403_/Q _3069_/S vssd1 vssd1 vccd1 vccd1 _2999_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold973 hold973/A vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__buf_2
XFILLER_1_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold962 hold962/A vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__buf_2
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold995 hold995/A vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__buf_2
Xhold984 hold984/A vssd1 vssd1 vccd1 vccd1 hold984/X sky130_fd_sc_hd__buf_2
XFILLER_1_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2330 hold992/X vssd1 vssd1 vccd1 vccd1 hold2330/X sky130_fd_sc_hd__buf_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2352 _4352_/X vssd1 vssd1 vccd1 vccd1 hold2352/X sky130_fd_sc_hd__buf_2
Xhold2341 hold2341/A vssd1 vssd1 vccd1 vccd1 hold2341/X sky130_fd_sc_hd__buf_2
Xhold1651 hold1651/A vssd1 vssd1 vccd1 vccd1 _5754_/D sky130_fd_sc_hd__buf_2
Xhold2385 hold2385/A vssd1 vssd1 vccd1 vccd1 _5750_/D sky130_fd_sc_hd__buf_2
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1640 hold2193/X vssd1 vssd1 vccd1 vccd1 hold2194/A sky130_fd_sc_hd__buf_2
Xhold1684 hold2216/X vssd1 vssd1 vccd1 vccd1 hold2217/A sky130_fd_sc_hd__buf_2
XFILLER_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1695 hold2345/X vssd1 vssd1 vccd1 vccd1 hold2346/A sky130_fd_sc_hd__buf_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4744__329 _4744__329/A vssd1 vssd1 vccd1 vccd1 _5435_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4638__223 _5007_/CLK vssd1 vssd1 vccd1 vccd1 _5316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3971_ _3971_/A _3989_/B vssd1 vssd1 vccd1 vccd1 _3971_/Y sky130_fd_sc_hd__nand2_8
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2922_ _5199_/Q _5183_/Q _4972_/Q _5191_/Q _3036_/S _2943_/S1 vssd1 vssd1 vccd1 vccd1
+ _2922_/X sky130_fd_sc_hd__mux4_2
X_5710_ _5710_/CLK _5710_/D vssd1 vssd1 vccd1 vccd1 _5710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5641_ _5641_/CLK _5641_/D vssd1 vssd1 vccd1 vccd1 _5641_/Q sky130_fd_sc_hd__dfxtp_1
X_2853_ _5392_/Q _2853_/A1 _2860_/S vssd1 vssd1 vccd1 vccd1 _5392_/D sky130_fd_sc_hd__mux2_1
X_5572_ _5572_/CLK _5572_/D vssd1 vssd1 vccd1 vccd1 _5572_/Q sky130_fd_sc_hd__dfxtp_1
X_2784_ _5452_/Q _2848_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5452_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XCaravelHost_654 vssd1 vssd1 vccd1 vccd1 CaravelHost_654/HI caravel_irq[3] sky130_fd_sc_hd__conb_1
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__buf_2
Xhold214 hold235/X vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__buf_2
Xhold225 _3628_/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__buf_2
XCaravelHost_665 vssd1 vssd1 vccd1 vccd1 CaravelHost_665/HI core1Index[3] sky130_fd_sc_hd__conb_1
XFILLER_132_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold258 hold276/X vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__buf_2
XCaravelHost_698 vssd1 vssd1 vccd1 vccd1 CaravelHost_698/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XCaravelHost_687 vssd1 vssd1 vccd1 vccd1 CaravelHost_687/HI la_data_out[115] sky130_fd_sc_hd__conb_1
XCaravelHost_676 vssd1 vssd1 vccd1 vccd1 CaravelHost_676/HI la_data_out[104] sky130_fd_sc_hd__conb_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__buf_2
XFILLER_132_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4385_ _5741_/Q _4389_/C _4385_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__o211a_1
X_3405_ _5274_/Q _3579_/A0 _3405_/S vssd1 vssd1 vccd1 vccd1 _5274_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _3336_/A1 _3317_/X _3320_/X _3335_/X _3136_/X vssd1 vssd1 vccd1 vccd1 _3336_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_140_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5006_/CLK _5006_/D vssd1 vssd1 vccd1 vccd1 _5006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _5419_/Q _2482_/B _3237_/B _5411_/Q _3282_/C1 vssd1 vssd1 vccd1 vccd1 _3267_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198_ _5342_/Q _3125_/A _3353_/A _3197_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3198_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5908_ _5908_/A vssd1 vssd1 vccd1 vccd1 _5908_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5839_ _5839_/A vssd1 vssd1 vccd1 vccd1 _5839_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2182 hold2796/X vssd1 vssd1 vccd1 vccd1 hold2797/A sky130_fd_sc_hd__buf_2
Xhold2171 hold2885/X vssd1 vssd1 vccd1 vccd1 hold2886/A sky130_fd_sc_hd__buf_2
XFILLER_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1470 hold13/X vssd1 vssd1 vccd1 vccd1 hold958/A sky130_fd_sc_hd__buf_2
Xhold2193 hold2807/X vssd1 vssd1 vccd1 vccd1 hold2193/X sky130_fd_sc_hd__buf_2
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1492 hold2264/X vssd1 vssd1 vccd1 vccd1 hold2265/A sky130_fd_sc_hd__buf_2
Xhold1481 hold2255/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__buf_2
XFILLER_72_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4872__457 _4892__477/A vssd1 vssd1 vccd1 vccd1 _5593_/CLK sky130_fd_sc_hd__inv_2
Xoutput308 _5877_/X vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_12
XFILLER_113_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput319 _5887_/X vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_12
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4170_/A _4170_/B _4170_/C _4170_/D vssd1 vssd1 vccd1 vccd1 _4177_/C sky130_fd_sc_hd__and4_1
X_4913__498 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5634_/CLK sky130_fd_sc_hd__inv_2
X_3121_ _3597_/A1 _5347_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5347_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3052_ _5210_/Q _5146_/Q _3063_/S vssd1 vssd1 vccd1 vccd1 _3052_/X sky130_fd_sc_hd__mux2_1
X_4501__86 _4509__94/A vssd1 vssd1 vccd1 vccd1 _5143_/CLK sky130_fd_sc_hd__inv_2
X_4766__351 _4786__371/A vssd1 vssd1 vccd1 vccd1 _5457_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3954_ _3827_/C split1/X _3920_/B vssd1 vssd1 vccd1 vccd1 _3954_/Y sky130_fd_sc_hd__a21oi_1
X_4807__392 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5498_/CLK sky130_fd_sc_hd__inv_2
X_2905_ _3043_/A _2900_/X _2904_/X _3094_/B vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__o211a_2
X_3885_ _5071_/Q _3959_/A _3885_/B1 vssd1 vssd1 vccd1 vccd1 _3885_/X sky130_fd_sc_hd__a21o_1
X_2836_ _3501_/A1 _5407_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5407_/D sky130_fd_sc_hd__mux2_1
X_5624_ _5624_/CLK _5624_/D vssd1 vssd1 vccd1 vccd1 _5624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5555_ _5557_/CLK _5555_/D vssd1 vssd1 vccd1 vccd1 _5555_/Q sky130_fd_sc_hd__dfxtp_2
X_2767_ _2788_/A _3397_/A vssd1 vssd1 vccd1 vccd1 _2775_/S sky130_fd_sc_hd__or2_4
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2698_ _5525_/Q _3566_/A1 _2702_/S vssd1 vssd1 vccd1 vccd1 _5525_/D sky130_fd_sc_hd__mux2_1
X_5486_ _5486_/CLK _5486_/D vssd1 vssd1 vccd1 vccd1 _5486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout513 _2460_/A vssd1 vssd1 vccd1 vccd1 _2867_/A sky130_fd_sc_hd__buf_8
Xfanout524 _5364_/Q vssd1 vssd1 vccd1 vccd1 _3005_/S sky130_fd_sc_hd__buf_8
XFILLER_59_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout502 split2/A vssd1 vssd1 vccd1 vccd1 split4/A sky130_fd_sc_hd__buf_8
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout557 _3779_/Y vssd1 vssd1 vccd1 vccd1 _3797_/A3 sky130_fd_sc_hd__buf_8
X_4368_ _4368_/A _5728_/Q vssd1 vssd1 vccd1 vccd1 _5734_/D sky130_fd_sc_hd__and2_1
Xfanout546 fanout547/X vssd1 vssd1 vccd1 vccd1 _3290_/S sky130_fd_sc_hd__buf_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout535 _3126_/A vssd1 vssd1 vccd1 vccd1 _3201_/S1 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4299_ _4298_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5669_/D sky130_fd_sc_hd__and2b_1
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _5647_/Q _2464_/Y _3326_/B2 _5639_/Q vssd1 vssd1 vccd1 vccd1 _3319_/X sky130_fd_sc_hd__o22a_1
Xfanout579 _5695_/Q vssd1 vssd1 vccd1 vccd1 _3402_/A1 sky130_fd_sc_hd__buf_6
Xfanout568 _3409_/A1 vssd1 vssd1 vccd1 vccd1 _3391_/A0 sky130_fd_sc_hd__clkbuf_8
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4600__185 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5274_/CLK sky130_fd_sc_hd__inv_2
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3670_ _3670_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3670_/X sky130_fd_sc_hd__and2_1
XFILLER_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2621_ _5370_/Q _2620_/Y _2862_/A vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5340_ _5340_/CLK _5340_/D vssd1 vssd1 vccd1 vccd1 _5340_/Q sky130_fd_sc_hd__dfxtp_1
X_2552_ _5658_/Q _3393_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _5658_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5271_ _5271_/CLK _5271_/D vssd1 vssd1 vccd1 vccd1 _5271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4222_ _4226_/B _4222_/B vssd1 vssd1 vccd1 vccd1 _4222_/X sky130_fd_sc_hd__or2_1
X_2483_ _5334_/Q _2463_/Y _2486_/A _3122_/C vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__a31o_1
Xhold2907 hold2907/A vssd1 vssd1 vccd1 vccd1 hold2907/X sky130_fd_sc_hd__buf_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4153_ _5741_/Q _4153_/B _4153_/C vssd1 vssd1 vccd1 vccd1 _4153_/X sky130_fd_sc_hd__and3_1
X_3104_ _5362_/Q _3599_/A1 _3111_/S vssd1 vssd1 vccd1 vccd1 _5362_/D sky130_fd_sc_hd__mux2_1
X_4084_ _5685_/Q _4088_/B vssd1 vssd1 vccd1 vccd1 _4084_/X sky130_fd_sc_hd__and2_1
XFILLER_56_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3035_ _2460_/A _5356_/Q _5123_/Q _3073_/B2 _3073_/C1 vssd1 vssd1 vccd1 vccd1 _3035_/X
+ sky130_fd_sc_hd__o221a_1
X_4417__2 _4418__3/A vssd1 vssd1 vccd1 vccd1 _4968_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4986_ _5019_/CLK _4986_/D vssd1 vssd1 vccd1 vccd1 _4986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4543__128 _4423__8/A vssd1 vssd1 vccd1 vccd1 _5185_/CLK sky130_fd_sc_hd__inv_2
X_3937_ _3937_/A0 _5094_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3937_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3868_ _5731_/Q _3857_/Y _3867_/X _3887_/B _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3868_/X
+ sky130_fd_sc_hd__a221o_1
X_3799_ hold277/X _5250_/Q _3810_/A3 hold349/X _4999_/Q vssd1 vssd1 vccd1 vccd1 _4999_/D
+ sky130_fd_sc_hd__o32a_1
X_5607_ _5607_/CLK _5607_/D vssd1 vssd1 vccd1 vccd1 _5607_/Q sky130_fd_sc_hd__dfxtp_1
X_2819_ _3391_/A0 _5422_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5422_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5538_ _5538_/CLK _5538_/D vssd1 vssd1 vccd1 vccd1 _5538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5469_ _5469_/CLK _5469_/D vssd1 vssd1 vccd1 vccd1 _5469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_55_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _5256_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4492__77 _4508__93/A vssd1 vssd1 vccd1 vccd1 _5134_/CLK sky130_fd_sc_hd__inv_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4878__463 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5599_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3722_ _5077_/Q input5/X _3728_/S vssd1 vssd1 vccd1 vccd1 _3722_/X sky130_fd_sc_hd__mux2_4
X_3653_ _3653_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3653_/X sky130_fd_sc_hd__or2_1
X_2604_ _3339_/A1 _5615_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5615_/D sky130_fd_sc_hd__mux2_1
X_3584_ _3584_/A0 _5038_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5038_/D sky130_fd_sc_hd__mux2_1
X_5323_ _5691_/CLK _5323_/D vssd1 vssd1 vccd1 vccd1 _5323_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_142_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2535_ _3406_/A _3370_/A vssd1 vssd1 vccd1 vccd1 _2543_/S sky130_fd_sc_hd__or2_4
X_5254_ _5256_/CLK _5254_/D vssd1 vssd1 vccd1 vccd1 _5254_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2466_ _3711_/B vssd1 vssd1 vccd1 vccd1 _2466_/Y sky130_fd_sc_hd__inv_2
X_5185_ _5185_/CLK _5185_/D vssd1 vssd1 vccd1 vccd1 _5185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4205_ _5549_/Q _4209_/B _4186_/X _4112_/Y vssd1 vssd1 vccd1 vccd1 _4206_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2748 _4393_/X vssd1 vssd1 vccd1 vccd1 hold2748/X sky130_fd_sc_hd__buf_2
X_4136_ _5540_/Q _5539_/Q vssd1 vssd1 vccd1 vccd1 _4137_/B sky130_fd_sc_hd__xor2_4
X_4067_ _4275_/B _4271_/C _4275_/C _4271_/D vssd1 vssd1 vccd1 vccd1 _4073_/C sky130_fd_sc_hd__and4_1
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3018_ _5211_/Q _5147_/Q _3063_/S vssd1 vssd1 vccd1 vccd1 _3018_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4969_ _4969_/CLK _4969_/D vssd1 vssd1 vccd1 vccd1 _4969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4459__44/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4671__256 _4514__99/A vssd1 vssd1 vccd1 vccd1 _5359_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4712__297 _4744__329/A vssd1 vssd1 vccd1 vccd1 _5403_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4565__150 _4509__94/A vssd1 vssd1 vccd1 vccd1 _5215_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606__191 _4463__48/A vssd1 vssd1 vccd1 vccd1 _5280_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5872_ _5872_/A vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4905__490/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3705_ _4988_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3705_/X sky130_fd_sc_hd__or2_1
XFILLER_134_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3636_ _4357_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3636_/X sky130_fd_sc_hd__or2_1
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3567_ _5053_/Q _3567_/A1 _3570_/S vssd1 vssd1 vccd1 vccd1 _5053_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2518_ _3574_/A0 _5721_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5721_/D sky130_fd_sc_hd__mux2_1
X_5306_ _5306_/CLK _5306_/D vssd1 vssd1 vccd1 vccd1 _5306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3498_ _3597_/A1 _5162_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5162_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5237_ _5237_/CLK _5237_/D vssd1 vssd1 vccd1 vccd1 _5237_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2501 hold799/X vssd1 vssd1 vccd1 vccd1 hold2501/X sky130_fd_sc_hd__buf_2
Xhold2512 hold2512/A vssd1 vssd1 vccd1 vccd1 hold2512/X sky130_fd_sc_hd__buf_2
XFILLER_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2523 hold2868/X vssd1 vssd1 vccd1 vccd1 hold2523/X sky130_fd_sc_hd__buf_2
Xhold1800 hold2514/X vssd1 vssd1 vccd1 vccd1 hold2515/A sky130_fd_sc_hd__buf_2
X_2449_ _5669_/Q vssd1 vssd1 vccd1 vccd1 _2449_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2556 hold2556/A vssd1 vssd1 vccd1 vccd1 _5755_/D sky130_fd_sc_hd__buf_2
X_5168_ _5168_/CLK _5168_/D vssd1 vssd1 vccd1 vccd1 _5168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2578 hold2578/A vssd1 vssd1 vccd1 vccd1 hold2578/X sky130_fd_sc_hd__buf_2
Xhold1844 hold1844/A vssd1 vssd1 vccd1 vccd1 hold786/A sky130_fd_sc_hd__buf_2
Xhold1822 hold727/X vssd1 vssd1 vccd1 vccd1 hold1822/X sky130_fd_sc_hd__buf_2
XFILLER_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1833 hold1833/A vssd1 vssd1 vccd1 vccd1 hold192/A sky130_fd_sc_hd__buf_2
Xhold2567 hold2567/A vssd1 vssd1 vccd1 vccd1 hold2567/X sky130_fd_sc_hd__buf_2
Xhold1877 hold585/X vssd1 vssd1 vccd1 vccd1 hold1877/X sky130_fd_sc_hd__buf_2
X_5099_ _5383_/CLK _5099_/D vssd1 vssd1 vccd1 vccd1 _5099_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1855 hold2585/X vssd1 vssd1 vccd1 vccd1 hold2586/A sky130_fd_sc_hd__buf_2
X_4119_ _5547_/Q _4132_/B _4119_/C vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__nand3_2
Xhold1866 hold193/X vssd1 vssd1 vccd1 vccd1 hold1866/X sky130_fd_sc_hd__buf_2
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4549__134 _4421__6/A vssd1 vssd1 vccd1 vccd1 _5191_/CLK sky130_fd_sc_hd__inv_2
Xhold1899 hold842/X vssd1 vssd1 vccd1 vccd1 hold1899/X sky130_fd_sc_hd__buf_2
Xhold1888 hold868/X vssd1 vssd1 vccd1 vccd1 hold1888/X sky130_fd_sc_hd__buf_2
X_4462__47 _4463__48/A vssd1 vssd1 vccd1 vccd1 _5056_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5684_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__buf_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3421_ _3594_/A1 _5237_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5237_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _5330_/Q _3357_/A _3169_/Y _4093_/B vssd1 vssd1 vccd1 vccd1 _5330_/D sky130_fd_sc_hd__o211a_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3283_ _3301_/A1 _3281_/X _3282_/X vssd1 vssd1 vccd1 vccd1 _3283_/X sky130_fd_sc_hd__o21a_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1107 hold2344/X vssd1 vssd1 vccd1 vccd1 hold2345/A sky130_fd_sc_hd__buf_2
X_5022_ _5022_/CLK hold81/X vssd1 vssd1 vccd1 vccd1 _5022_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _5924_/A vssd1 vssd1 vccd1 vccd1 _5924_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5855_ _5855_/A vssd1 vssd1 vccd1 vccd1 _5855_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5025_/CLK sky130_fd_sc_hd__clkbuf_8
X_2998_ _3034_/A _2996_/X _2997_/X vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3619_ _4389_/B _3617_/B _3618_/X _4966_/Q vssd1 vssd1 vccd1 vccd1 _3619_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold963 hold963/A vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__buf_2
X_4507__92 _4507__92/A vssd1 vssd1 vccd1 vccd1 _5149_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold996 hold996/A vssd1 vssd1 vccd1 vccd1 hold996/X sky130_fd_sc_hd__buf_2
Xhold985 hold985/A vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__buf_2
Xhold974 hold974/A vssd1 vssd1 vccd1 vccd1 hold974/X sky130_fd_sc_hd__buf_2
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2320 hold723/X vssd1 vssd1 vccd1 vccd1 hold2320/X sky130_fd_sc_hd__buf_2
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2331 hold2331/A vssd1 vssd1 vccd1 vccd1 input166/A sky130_fd_sc_hd__buf_2
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2353 hold2353/A vssd1 vssd1 vccd1 vccd1 hold2353/X sky130_fd_sc_hd__buf_2
Xhold2342 hold2342/A vssd1 vssd1 vccd1 vccd1 hold748/A sky130_fd_sc_hd__buf_2
Xhold1630 hold2206/X vssd1 vssd1 vccd1 vccd1 hold2207/A sky130_fd_sc_hd__buf_2
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2386 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 hold2386/X sky130_fd_sc_hd__buf_2
Xhold1641 hold2195/X vssd1 vssd1 vccd1 vccd1 hold2196/A sky130_fd_sc_hd__buf_2
Xhold1685 hold2218/X vssd1 vssd1 vccd1 vccd1 hold2219/A sky130_fd_sc_hd__buf_2
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4783__368 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5474_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4677__262 _4425__10/A vssd1 vssd1 vccd1 vccd1 _5366_/CLK sky130_fd_sc_hd__inv_2
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _5382_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _5209_/D sky130_fd_sc_hd__and2_1
XFILLER_51_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2921_ _5063_/Q _5039_/Q _5536_/Q _4980_/Q _2941_/S0 _3024_/S vssd1 vssd1 vccd1 vccd1
+ _2921_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5640_ _5640_/CLK _5640_/D vssd1 vssd1 vccd1 vccd1 _5640_/Q sky130_fd_sc_hd__dfxtp_1
X_4918__503 _4457__42/A vssd1 vssd1 vccd1 vccd1 _5639_/CLK sky130_fd_sc_hd__inv_2
X_2852_ _2852_/A _3397_/A vssd1 vssd1 vccd1 vccd1 _2860_/S sky130_fd_sc_hd__nor2_8
X_5571_ _5571_/CLK _5571_/D vssd1 vssd1 vccd1 vccd1 _5571_/Q sky130_fd_sc_hd__dfxtp_1
X_2783_ _5453_/Q _3602_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5453_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__buf_2
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_655 vssd1 vssd1 vccd1 vccd1 CaravelHost_655/HI core0Index[0] sky130_fd_sc_hd__conb_1
Xhold215 hold223/X vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__buf_2
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold675/A sky130_fd_sc_hd__buf_2
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold259 _3802_/X vssd1 vssd1 vccd1 vccd1 _5002_/D sky130_fd_sc_hd__buf_2
Xhold248 hold271/X vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__buf_2
XCaravelHost_688 vssd1 vssd1 vccd1 vccd1 CaravelHost_688/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XCaravelHost_677 vssd1 vssd1 vccd1 vccd1 CaravelHost_677/HI la_data_out[105] sky130_fd_sc_hd__conb_1
X_3404_ _5275_/Q _3569_/A1 _3405_/S vssd1 vssd1 vccd1 vccd1 _5275_/D sky130_fd_sc_hd__mux2_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__buf_2
XCaravelHost_666 vssd1 vssd1 vccd1 vccd1 CaravelHost_666/HI core1Index[4] sky130_fd_sc_hd__conb_1
XFILLER_113_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_699 vssd1 vssd1 vccd1 vccd1 CaravelHost_699/HI la_data_out[127] sky130_fd_sc_hd__conb_1
X_4384_ _3643_/A _4389_/B _4398_/A2 vssd1 vssd1 vccd1 vccd1 _4384_/X sky130_fd_sc_hd__a21bo_1
XFILLER_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3335_ _3325_/X _3326_/X _3353_/B _3323_/X vssd1 vssd1 vccd1 vccd1 _3335_/X sky130_fd_sc_hd__a211o_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3328_/A _3266_/B vssd1 vssd1 vccd1 vccd1 _3266_/X sky130_fd_sc_hd__or2_1
X_5005_ _5005_/CLK _5005_/D vssd1 vssd1 vccd1 vccd1 _5005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ _3136_/X _3191_/X _3195_/X _3196_/X vssd1 vssd1 vccd1 vccd1 _3197_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5907_ _5907_/A vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__clkbuf_4
X_4432__17 _4432__17/A vssd1 vssd1 vccd1 vccd1 _5026_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5838_ _5838_/A vssd1 vssd1 vccd1 vccd1 _5838_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold760 hold760/A vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__buf_2
Xhold782 hold782/A vssd1 vssd1 vccd1 vccd1 hold782/X sky130_fd_sc_hd__buf_2
Xhold793 hold793/A vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__buf_2
XFILLER_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2172 hold2789/X vssd1 vssd1 vccd1 vccd1 hold2790/A sky130_fd_sc_hd__buf_2
Xhold2183 hold2798/X vssd1 vssd1 vccd1 vccd1 hold2799/A sky130_fd_sc_hd__buf_2
Xhold2194 hold2194/A vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__buf_2
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1493 hold969/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__buf_2
Xhold1482 hold19/X vssd1 vssd1 vccd1 vccd1 hold964/A sky130_fd_sc_hd__buf_2
Xhold1471 hold958/X vssd1 vssd1 vccd1 vccd1 _3934_/A0 sky130_fd_sc_hd__buf_2
XFILLER_33_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput309 _5878_/X vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_12
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4498__83 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5140_/CLK sky130_fd_sc_hd__inv_2
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3120_ _3596_/A1 _5348_/Q _3121_/S vssd1 vssd1 vccd1 vccd1 _5348_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _3099_/B _3049_/X _3050_/X vssd1 vssd1 vccd1 vccd1 _3051_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3953_ _5257_/Q _5110_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _5110_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2904_ _2947_/S _2901_/X _2903_/X vssd1 vssd1 vccd1 vccd1 _2904_/X sky130_fd_sc_hd__a21o_1
X_3884_ _4399_/B _3881_/X _3883_/X _4361_/A vssd1 vssd1 vccd1 vccd1 _3884_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2835_ _3536_/A0 _5408_/Q _2842_/S vssd1 vssd1 vccd1 vccd1 _5408_/D sky130_fd_sc_hd__mux2_1
X_5623_ _5623_/CLK _5623_/D vssd1 vssd1 vccd1 vccd1 _5623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5554_ _5566_/CLK _5554_/D vssd1 vssd1 vccd1 vccd1 _5554_/Q sky130_fd_sc_hd__dfxtp_1
X_2766_ _3396_/A0 _5465_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5465_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2697_ _5526_/Q _3409_/A1 _2702_/S vssd1 vssd1 vccd1 vccd1 _5526_/D sky130_fd_sc_hd__mux2_1
X_5485_ _5485_/CLK _5485_/D vssd1 vssd1 vccd1 vccd1 _5485_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout514 _5366_/Q vssd1 vssd1 vccd1 vccd1 _2460_/A sky130_fd_sc_hd__buf_8
X_4367_ _4368_/A _5727_/Q vssd1 vssd1 vccd1 vccd1 _5733_/D sky130_fd_sc_hd__and2_1
XFILLER_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout503 _3777_/A3 vssd1 vssd1 vccd1 vccd1 split2/A sky130_fd_sc_hd__buf_12
Xfanout525 _3002_/S vssd1 vssd1 vccd1 vccd1 _3072_/S sky130_fd_sc_hd__buf_6
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout536 _3126_/A vssd1 vssd1 vccd1 vccd1 _3127_/A sky130_fd_sc_hd__buf_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout547 _5326_/Q vssd1 vssd1 vccd1 vccd1 fanout547/X sky130_fd_sc_hd__buf_6
X_3318_ _5042_/Q _5631_/Q _3318_/S vssd1 vssd1 vccd1 vccd1 _3318_/X sky130_fd_sc_hd__mux2_1
X_4298_ _4262_/B _4308_/A2 _4308_/B1 _2449_/Y vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__o22a_1
Xfanout558 _3897_/C vssd1 vssd1 vccd1 vccd1 _3882_/A3 sky130_fd_sc_hd__buf_4
XFILLER_59_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout569 _3574_/A0 vssd1 vssd1 vccd1 vccd1 _2743_/A0 sky130_fd_sc_hd__buf_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3249_ _3301_/A1 _3247_/X _3248_/X vssd1 vssd1 vccd1 vccd1 _3249_/X sky130_fd_sc_hd__o21a_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold590 hold590/A vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__buf_2
XFILLER_110_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4789__374 _5697_/CLK vssd1 vssd1 vccd1 vccd1 _5480_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1290 hold2541/X vssd1 vssd1 vccd1 vccd1 hold2542/A sky130_fd_sc_hd__buf_2
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2620_ _2861_/A vssd1 vssd1 vccd1 vccd1 _2620_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2551_ _5659_/Q _5696_/Q _2555_/S vssd1 vssd1 vccd1 vccd1 _5659_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5270_ _5270_/CLK _5270_/D vssd1 vssd1 vccd1 vccd1 _5270_/Q sky130_fd_sc_hd__dfxtp_1
X_2482_ _3346_/A _2482_/B vssd1 vssd1 vccd1 vccd1 _3123_/C sky130_fd_sc_hd__xor2_2
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4221_ _4244_/S _4221_/B _4221_/C vssd1 vssd1 vccd1 vccd1 _5555_/D sky130_fd_sc_hd__and3_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2908 hold2908/A vssd1 vssd1 vccd1 vccd1 hold2908/X sky130_fd_sc_hd__buf_2
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4152_ _4153_/B _4153_/C _5741_/Q vssd1 vssd1 vccd1 vccd1 _4152_/Y sky130_fd_sc_hd__a21oi_2
X_3103_ _3598_/A _3535_/B vssd1 vssd1 vccd1 vccd1 _3111_/S sky130_fd_sc_hd__nor2_8
X_4083_ _5684_/Q _4088_/B vssd1 vssd1 vccd1 vccd1 _4083_/X sky130_fd_sc_hd__and2_1
XFILLER_83_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3034_ _3034_/A _3034_/B vssd1 vssd1 vccd1 vccd1 _3034_/X sky130_fd_sc_hd__or2_1
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4985_ _5024_/CLK _4985_/D vssd1 vssd1 vccd1 vccd1 _4985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4582__167 _4510__95/A vssd1 vssd1 vccd1 vccd1 _5232_/CLK sky130_fd_sc_hd__inv_2
X_3936_ _3936_/A0 _5093_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3867_ _3998_/A1 _5204_/Q _3882_/A3 _3855_/X vssd1 vssd1 vccd1 vccd1 _3867_/X sky130_fd_sc_hd__a31o_1
X_5606_ _5606_/CLK _5606_/D vssd1 vssd1 vccd1 vccd1 _5606_/Q sky130_fd_sc_hd__dfxtp_1
X_3798_ hold277/X _5249_/Q _3810_/A3 hold349/X _4998_/Q vssd1 vssd1 vccd1 vccd1 _4998_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2818_ _3390_/A0 _5423_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5423_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5537_ _5537_/CLK _5537_/D vssd1 vssd1 vccd1 vccd1 _5537_/Q sky130_fd_sc_hd__dfxtp_1
X_2749_ _2788_/A _3370_/A vssd1 vssd1 vccd1 vccd1 _2757_/S sky130_fd_sc_hd__or2_4
XFILLER_105_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5468_ _5468_/CLK _5468_/D vssd1 vssd1 vccd1 vccd1 _5468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5399_ _5399_/CLK _5399_/D vssd1 vssd1 vccd1 vccd1 _5399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_95_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4897__482/A
+ sky130_fd_sc_hd__clkbuf_16
X_4823__408 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5514_/CLK sky130_fd_sc_hd__inv_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4433__18/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4717__302 _5010_/CLK vssd1 vssd1 vccd1 vccd1 _5408_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4468__53 _4468__53/A vssd1 vssd1 vccd1 vccd1 _5062_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3721_ _3733_/A1 _3719_/X _3720_/X split2/A vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__o211a_1
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3652_ _3652_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3652_/X sky130_fd_sc_hd__or2_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3583_ _3601_/A1 _5039_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5039_/D sky130_fd_sc_hd__mux2_1
X_2603_ _3569_/A1 _5616_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5616_/D sky130_fd_sc_hd__mux2_1
X_5322_ _5691_/CLK _5322_/D vssd1 vssd1 vccd1 vccd1 _5322_/Q sky130_fd_sc_hd__dfxtp_2
X_2534_ _5332_/Q _5331_/Q _3350_/B split3/A vssd1 vssd1 vccd1 vccd1 _3370_/A sky130_fd_sc_hd__or4b_4
XFILLER_114_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5253_ _5256_/CLK _5253_/D vssd1 vssd1 vccd1 vccd1 _5253_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2465_ _3920_/B vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__inv_4
X_5184_ _5184_/CLK _5184_/D vssd1 vssd1 vccd1 vccd1 _5184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4204_ _4204_/A _4204_/B vssd1 vssd1 vccd1 vccd1 _5548_/D sky130_fd_sc_hd__nor2_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _5752_/Q _4135_/B vssd1 vssd1 vccd1 vccd1 _4171_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _5751_/Q _4262_/B vssd1 vssd1 vccd1 vccd1 _4271_/D sky130_fd_sc_hd__xor2_2
X_3017_ _3595_/A1 _2895_/Y _3016_/X _3080_/B1 vssd1 vssd1 vccd1 vccd1 _5377_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _4968_/CLK _4968_/D vssd1 vssd1 vccd1 vccd1 _4968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3919_ _5083_/Q _3926_/A2 _3923_/B1 _3918_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5083_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951__536 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5709_/CLK sky130_fd_sc_hd__inv_2
XFILLER_124_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4845__430 _5002_/CLK vssd1 vssd1 vccd1 vccd1 _5538_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5871_ _5871_/A vssd1 vssd1 vccd1 vccd1 _5871_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3704_ _5071_/Q input30/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3704_/X sky130_fd_sc_hd__mux2_4
XFILLER_147_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3635_ _4356_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3635_/X sky130_fd_sc_hd__or2_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3566_ _5054_/Q _3566_/A1 _3570_/S vssd1 vssd1 vccd1 vccd1 _5054_/D sky130_fd_sc_hd__mux2_1
X_4694__279 _5244_/CLK vssd1 vssd1 vccd1 vccd1 _5385_/CLK sky130_fd_sc_hd__inv_2
XFILLER_130_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3497_ _3596_/A1 _5163_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5163_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2517_ _3564_/A1 _5722_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5722_/D sky130_fd_sc_hd__mux2_1
X_5305_ _5305_/CLK _5305_/D vssd1 vssd1 vccd1 vccd1 _5305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5236_ _5236_/CLK _5236_/D vssd1 vssd1 vccd1 vccd1 _5236_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2502 hold2502/A vssd1 vssd1 vccd1 vccd1 hold2502/X sky130_fd_sc_hd__buf_2
Xhold2513 hold2513/A vssd1 vssd1 vccd1 vccd1 hold816/A sky130_fd_sc_hd__buf_2
X_2448_ _5670_/Q vssd1 vssd1 vccd1 vccd1 _2448_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2524 hold2524/A vssd1 vssd1 vccd1 vccd1 hold2524/X sky130_fd_sc_hd__buf_2
Xhold1801 hold2516/X vssd1 vssd1 vccd1 vccd1 hold2517/A sky130_fd_sc_hd__buf_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5167_ _5167_/CLK _5167_/D vssd1 vssd1 vccd1 vccd1 _5167_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1845 hold786/X vssd1 vssd1 vccd1 vccd1 hold1845/X sky130_fd_sc_hd__buf_2
Xhold2579 hold2579/A vssd1 vssd1 vccd1 vccd1 _5724_/D sky130_fd_sc_hd__buf_2
Xhold1823 hold1823/A vssd1 vssd1 vccd1 vccd1 _4372_/B1 sky130_fd_sc_hd__buf_2
XFILLER_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2568 hold2568/A vssd1 vssd1 vccd1 vccd1 hold2568/X sky130_fd_sc_hd__buf_2
Xhold1834 hold192/X vssd1 vssd1 vccd1 vccd1 hold1834/X sky130_fd_sc_hd__buf_2
Xhold1878 hold1878/A vssd1 vssd1 vccd1 vccd1 _5739_/D sky130_fd_sc_hd__buf_2
X_5098_ _5384_/CLK _5098_/D vssd1 vssd1 vccd1 vccd1 _5098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1856 hold2587/X vssd1 vssd1 vccd1 vccd1 hold2588/A sky130_fd_sc_hd__buf_2
X_4118_ _4169_/A _4118_/B _4118_/C _4169_/B vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__and4_1
Xhold1867 hold1867/A vssd1 vssd1 vccd1 vccd1 _5024_/D sky130_fd_sc_hd__buf_2
X_4588__173 _5111_/CLK vssd1 vssd1 vccd1 vccd1 _5238_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4049_ _4254_/B _4254_/C _5750_/Q vssd1 vssd1 vccd1 vccd1 _4049_/Y sky130_fd_sc_hd__a21oi_1
Xhold1889 hold1889/A vssd1 vssd1 vccd1 vccd1 _5745_/D sky130_fd_sc_hd__buf_2
XFILLER_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__buf_2
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4829__414 _4909__494/A vssd1 vssd1 vccd1 vccd1 _5520_/CLK sky130_fd_sc_hd__inv_2
X_4438__23 _4438__23/A vssd1 vssd1 vccd1 vccd1 _5032_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold408 _3962_/Y vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__buf_2
XFILLER_143_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3420_ _3593_/A1 _5238_/Q _3424_/S vssd1 vssd1 vccd1 vccd1 _5238_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3351_ _2489_/Y split3/X _3351_/C vssd1 vssd1 vccd1 vccd1 _5331_/D sky130_fd_sc_hd__and3b_1
XFILLER_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3282_ _5506_/Q _2482_/B _3298_/B1 _5498_/Q _3282_/C1 vssd1 vssd1 vccd1 vccd1 _3282_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1119 hold2778/X vssd1 vssd1 vccd1 vccd1 hold1119/X sky130_fd_sc_hd__buf_2
X_5021_ _5022_/CLK _5021_/D vssd1 vssd1 vccd1 vccd1 _5021_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5923_ _5923_/A vssd1 vssd1 vccd1 vccd1 _5923_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5854_ _5854_/A vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4622__207 _4964__549/A vssd1 vssd1 vccd1 vccd1 _5299_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2997_ _5601_/Q _2460_/A _3073_/B2 _5585_/Q _3073_/C1 vssd1 vssd1 vccd1 vccd1 _2997_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3618_ _5258_/Q _5259_/Q _5260_/Q _5261_/Q vssd1 vssd1 vccd1 vccd1 _3618_/X sky130_fd_sc_hd__and4_4
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold953 hold953/A vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__buf_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold964 hold964/A vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__buf_2
XFILLER_131_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3549_ _5117_/Q _3594_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5117_/D sky130_fd_sc_hd__mux2_1
X_4516__101 _4485__70/A vssd1 vssd1 vccd1 vccd1 _5158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold975 hold975/A vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__buf_2
Xhold986 hold986/A vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__buf_2
Xhold997 hold997/A vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__buf_2
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2310 hold2310/A vssd1 vssd1 vccd1 vccd1 _5697_/D sky130_fd_sc_hd__buf_2
Xhold2321 hold2321/A vssd1 vssd1 vccd1 vccd1 hold2321/X sky130_fd_sc_hd__buf_2
X_5219_ _5219_/CLK _5219_/D vssd1 vssd1 vccd1 vccd1 _5219_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2354 hold2354/A vssd1 vssd1 vccd1 vccd1 hold2354/X sky130_fd_sc_hd__buf_2
Xhold2343 hold748/X vssd1 vssd1 vccd1 vccd1 hold2343/X sky130_fd_sc_hd__buf_2
Xhold2332 _3670_/A vssd1 vssd1 vccd1 vccd1 hold2332/X sky130_fd_sc_hd__buf_2
Xhold1631 hold2208/X vssd1 vssd1 vccd1 vccd1 hold2209/A sky130_fd_sc_hd__buf_2
Xhold2387 hold2387/A vssd1 vssd1 vccd1 vccd1 hold985/A sky130_fd_sc_hd__buf_2
Xhold1642 hold2197/X vssd1 vssd1 vccd1 vccd1 hold2198/A sky130_fd_sc_hd__buf_2
Xhold2365 _4350_/X vssd1 vssd1 vccd1 vccd1 hold2365/X sky130_fd_sc_hd__buf_2
Xhold1686 hold2220/X vssd1 vssd1 vccd1 vccd1 hold2221/A sky130_fd_sc_hd__buf_2
Xhold1675 hold2352/X vssd1 vssd1 vccd1 vccd1 hold2353/A sky130_fd_sc_hd__buf_2
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2920_ _5588_/Q _5572_/Q _5454_/Q _5604_/Q _3024_/S _2941_/S0 vssd1 vssd1 vccd1 vccd1
+ _2920_/X sky130_fd_sc_hd__mux4_2
X_2851_ _5393_/Q _3543_/A0 _2851_/S vssd1 vssd1 vccd1 vccd1 _5393_/D sky130_fd_sc_hd__mux2_1
X_4957__542 _5697_/CLK vssd1 vssd1 vccd1 vccd1 _5715_/CLK sky130_fd_sc_hd__inv_2
X_2782_ _5454_/Q _3601_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5454_/D sky130_fd_sc_hd__mux2_1
X_5570_ _5570_/CLK _5570_/D vssd1 vssd1 vccd1 vccd1 _5570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__buf_2
XCaravelHost_656 vssd1 vssd1 vccd1 vccd1 CaravelHost_656/HI core0Index[1] sky130_fd_sc_hd__conb_1
Xhold216 hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__buf_2
Xhold249 hold275/X vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__buf_2
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__buf_2
XCaravelHost_689 vssd1 vssd1 vccd1 vccd1 CaravelHost_689/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XCaravelHost_678 vssd1 vssd1 vccd1 vccd1 CaravelHost_678/HI la_data_out[106] sky130_fd_sc_hd__conb_1
X_3403_ _5276_/Q _3577_/A0 _3405_/S vssd1 vssd1 vccd1 vccd1 _5276_/D sky130_fd_sc_hd__mux2_1
XCaravelHost_667 vssd1 vssd1 vccd1 vccd1 CaravelHost_667/HI core1Index[5] sky130_fd_sc_hd__conb_1
XFILLER_113_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4383_ _5740_/Q _4389_/C _4383_/B1 _3778_/A vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__o211a_1
XFILLER_112_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3334_/A1 _3311_/X _3314_/X _3333_/X _3169_/B vssd1 vssd1 vccd1 vccd1 _3334_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _5657_/Q _5387_/Q _3327_/S vssd1 vssd1 vccd1 vccd1 _3266_/B sky130_fd_sc_hd__mux2_1
X_5004_ _5004_/CLK _5004_/D vssd1 vssd1 vccd1 vccd1 _5004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3334_/A1 _3183_/X _3185_/X _3187_/X _3169_/B vssd1 vssd1 vccd1 vccd1 _3196_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5906_ _5906_/A vssd1 vssd1 vccd1 vccd1 _5906_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5837_ _5837_/A vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5699_ _5751_/CLK _5699_/D vssd1 vssd1 vccd1 vccd1 _5699_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_49_wb_clk_i clkbuf_4_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5004_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750__335 _4786__371/A vssd1 vssd1 vccd1 vccd1 _5441_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2173 hold2791/X vssd1 vssd1 vccd1 vccd1 hold2792/A sky130_fd_sc_hd__buf_2
XFILLER_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2184 hold2800/X vssd1 vssd1 vccd1 vccd1 hold2801/A sky130_fd_sc_hd__buf_2
Xhold1450 hold453/X vssd1 vssd1 vccd1 vccd1 _4403_/B1 sky130_fd_sc_hd__buf_2
Xhold2195 hold186/X vssd1 vssd1 vccd1 vccd1 hold2195/X sky130_fd_sc_hd__buf_2
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1472 _3934_/X vssd1 vssd1 vccd1 vccd1 hold959/A sky130_fd_sc_hd__buf_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1494 hold25/X vssd1 vssd1 vccd1 vccd1 hold970/A sky130_fd_sc_hd__buf_2
Xhold1483 hold964/X vssd1 vssd1 vccd1 vccd1 _3935_/A0 sky130_fd_sc_hd__buf_2
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _5226_/Q _2866_/A _2866_/B _5114_/Q _3097_/B vssd1 vssd1 vccd1 vccd1 _3050_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _5256_/Q _5109_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _5109_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2903_ _2945_/A _2902_/X _2919_/B vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__a21o_1
X_3883_ _5734_/Q _3857_/Y _3882_/X _3887_/B _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3883_/X
+ sky130_fd_sc_hd__a221o_1
X_2834_ _3508_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2842_/S sky130_fd_sc_hd__or2_4
X_5622_ _5622_/CLK _5622_/D vssd1 vssd1 vccd1 vccd1 _5622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5553_ _5553_/CLK _5553_/D vssd1 vssd1 vccd1 vccd1 _5553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2765_ _3395_/A0 _5466_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5466_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4734__319 _5005_/CLK vssd1 vssd1 vccd1 vccd1 _5425_/CLK sky130_fd_sc_hd__inv_2
X_2696_ _5527_/Q _3573_/A0 _2702_/S vssd1 vssd1 vccd1 vccd1 _5527_/D sky130_fd_sc_hd__mux2_1
X_5484_ _5484_/CLK _5484_/D vssd1 vssd1 vccd1 vccd1 _5484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout515 _2867_/B vssd1 vssd1 vccd1 vccd1 _2944_/S0 sky130_fd_sc_hd__clkbuf_16
Xfanout504 _3777_/A3 vssd1 vssd1 vccd1 vccd1 _3766_/C1 sky130_fd_sc_hd__buf_8
X_4366_ _4368_/A _5726_/Q vssd1 vssd1 vccd1 vccd1 _5732_/D sky130_fd_sc_hd__and2_1
Xfanout526 _3002_/S vssd1 vssd1 vccd1 vccd1 _3024_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout548 _4282_/Y vssd1 vssd1 vccd1 vccd1 _4308_/B1 sky130_fd_sc_hd__buf_4
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3325_/A _3315_/X _3316_/X vssd1 vssd1 vccd1 vccd1 _3317_/X sky130_fd_sc_hd__o21a_1
Xfanout537 _5327_/Q vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__buf_6
XFILLER_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4297_ _4296_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5668_/D sky130_fd_sc_hd__and2b_1
Xfanout559 _2501_/X vssd1 vssd1 vccd1 vccd1 _3897_/C sky130_fd_sc_hd__buf_6
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _5507_/Q _2482_/B _3298_/B1 _5499_/Q _3282_/C1 vssd1 vssd1 vccd1 vccd1 _3248_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3179_ _5343_/Q _3125_/A _3353_/A _3178_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3179_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4628__213 _4460__45/A vssd1 vssd1 vccd1 vccd1 _5305_/CLK sky130_fd_sc_hd__inv_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold580 hold580/A vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__buf_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2550_ _5660_/Q _3391_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _5660_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2481_ _5334_/Q _2463_/Y _3122_/C _2486_/A vssd1 vssd1 vccd1 vccd1 _2487_/B sky130_fd_sc_hd__o211a_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4220_ _5555_/Q _4220_/B vssd1 vssd1 vccd1 vccd1 _4221_/C sky130_fd_sc_hd__nand2_1
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4151_ _4153_/B _4153_/C vssd1 vssd1 vccd1 vccd1 _4151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3102_ _3066_/S _3099_/A _3101_/Y vssd1 vssd1 vccd1 vccd1 _5364_/D sky130_fd_sc_hd__a21oi_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4082_ _4082_/A _4325_/A vssd1 vssd1 vccd1 vccd1 _5309_/D sky130_fd_sc_hd__and2_1
X_3033_ _5155_/Q _5311_/Q _3072_/S vssd1 vssd1 vccd1 vccd1 _3034_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4984_ _5016_/CLK _4984_/D vssd1 vssd1 vccd1 vccd1 _4984_/Q sky130_fd_sc_hd__dfxtp_1
X_3935_ _3935_/A0 _5092_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3935_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5605_ _5605_/CLK _5605_/D vssd1 vssd1 vccd1 vccd1 _5605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3866_ _5753_/Q _3998_/A1 _3882_/A3 _3887_/A vssd1 vssd1 vccd1 vccd1 _3866_/X sky130_fd_sc_hd__a31o_1
X_2817_ _3389_/A0 _5424_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _5424_/D sky130_fd_sc_hd__mux2_1
X_3797_ _4360_/A _5248_/Q _3797_/A3 hold364/X _4997_/Q vssd1 vssd1 vccd1 vccd1 _3797_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5536_ _5536_/CLK _5536_/D vssd1 vssd1 vccd1 vccd1 _5536_/Q sky130_fd_sc_hd__dfxtp_1
X_2748_ _3339_/A1 _5481_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5481_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5467_/CLK _5467_/D vssd1 vssd1 vccd1 vccd1 _5467_/Q sky130_fd_sc_hd__dfxtp_1
X_2679_ _2848_/A1 _5570_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5570_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5398_ _5398_/CLK _5398_/D vssd1 vssd1 vccd1 vccd1 _5398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4349_ _4281_/X _4324_/X _4348_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5691_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4862__447 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5583_/CLK sky130_fd_sc_hd__inv_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903__488 _4937__522/A vssd1 vssd1 vccd1 vccd1 _5624_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5007_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4756__341 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5447_/CLK sky130_fd_sc_hd__inv_2
XFILLER_136_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4483__68 _5006_/CLK vssd1 vssd1 vccd1 vccd1 _5125_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _4993_/Q _3729_/B vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__or2_1
XFILLER_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ _3651_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3651_/X sky130_fd_sc_hd__or2_1
X_3582_ _3600_/A1 _5040_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5040_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2602_ _3577_/A0 _5617_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5617_/D sky130_fd_sc_hd__mux2_1
X_5321_ _5691_/CLK _5321_/D vssd1 vssd1 vccd1 vccd1 _5321_/Q sky130_fd_sc_hd__dfxtp_4
X_2533_ _3396_/A0 _5708_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5708_/D sky130_fd_sc_hd__mux2_1
X_5252_ _5252_/CLK _5252_/D vssd1 vssd1 vccd1 vccd1 _5252_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2464_ _2464_/A vssd1 vssd1 vccd1 vccd1 _2464_/Y sky130_fd_sc_hd__inv_2
X_5183_ _5183_/CLK _5183_/D vssd1 vssd1 vccd1 vccd1 _5183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2706 _4093_/X vssd1 vssd1 vccd1 vccd1 hold2706/X sky130_fd_sc_hd__buf_2
X_4203_ _5548_/Q _4187_/B1 _4186_/X _4157_/B vssd1 vssd1 vccd1 vccd1 _4204_/B sky130_fd_sc_hd__o2bb2a_1
Xhold2717 hold2720/X vssd1 vssd1 vccd1 vccd1 _2467_/A sky130_fd_sc_hd__buf_2
XFILLER_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2739 hold191/X vssd1 vssd1 vccd1 vccd1 hold2739/X sky130_fd_sc_hd__buf_2
X_4134_ _5542_/Q _4142_/B vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__xor2_2
XFILLER_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4065_ _5669_/Q _4065_/B vssd1 vssd1 vccd1 vccd1 _4262_/B sky130_fd_sc_hd__xnor2_4
X_3016_ _2863_/A _5377_/Q _3094_/A _3015_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _3016_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_71_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _4967_/CLK _4967_/D vssd1 vssd1 vccd1 vccd1 _4967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3918_ _5738_/Q _3920_/B _5292_/Q vssd1 vssd1 vccd1 vccd1 _3918_/X sky130_fd_sc_hd__and3_1
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3849_ _5090_/Q _3959_/B vssd1 vssd1 vccd1 vccd1 _3850_/D sky130_fd_sc_hd__nand2_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _5519_/CLK _5519_/D vssd1 vssd1 vccd1 vccd1 _5519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_111_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4941__526/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4533__118 _5111_/CLK vssd1 vssd1 vccd1 vccd1 _5175_/CLK sky130_fd_sc_hd__inv_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5870_ _5870_/A vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3703_ _3718_/A1 _3701_/X _3702_/X split4/X vssd1 vssd1 vccd1 vccd1 _3703_/X sky130_fd_sc_hd__o211a_1
XFILLER_147_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3634_ _4355_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3634_/X sky130_fd_sc_hd__or2_1
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3565_ _5055_/Q _3574_/A0 _3570_/S vssd1 vssd1 vccd1 vccd1 _5055_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3496_ _3595_/A1 _5164_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5164_/D sky130_fd_sc_hd__mux2_1
X_2516_ _3572_/A0 _5723_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _5723_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5304_ _5304_/CLK _5304_/D vssd1 vssd1 vccd1 vccd1 _5304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5235_ _5235_/CLK _5235_/D vssd1 vssd1 vccd1 vccd1 _5235_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2503 hold2503/A vssd1 vssd1 vccd1 vccd1 hold2503/X sky130_fd_sc_hd__buf_2
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2447_ _5671_/Q vssd1 vssd1 vccd1 vccd1 _4034_/A sky130_fd_sc_hd__inv_2
XFILLER_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2525 hold2525/A vssd1 vssd1 vccd1 vccd1 hold2525/X sky130_fd_sc_hd__buf_2
Xhold2536 hold2862/X vssd1 vssd1 vccd1 vccd1 hold2536/X sky130_fd_sc_hd__buf_2
Xhold2514 hold816/X vssd1 vssd1 vccd1 vccd1 hold2514/X sky130_fd_sc_hd__buf_2
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5166_ _5166_/CLK _5166_/D vssd1 vssd1 vccd1 vccd1 _5166_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1813 hold2572/X vssd1 vssd1 vccd1 vccd1 hold2573/A sky130_fd_sc_hd__buf_2
Xhold1824 _4372_/X vssd1 vssd1 vccd1 vccd1 hold1824/X sky130_fd_sc_hd__buf_2
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2569 hold2569/A vssd1 vssd1 vccd1 vccd1 _5753_/D sky130_fd_sc_hd__buf_2
Xhold1835 hold1835/A vssd1 vssd1 vccd1 vccd1 _3830_/B sky130_fd_sc_hd__buf_2
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1846 hold1846/A vssd1 vssd1 vccd1 vccd1 _4378_/B1 sky130_fd_sc_hd__buf_2
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5097_ _5384_/CLK _5097_/D vssd1 vssd1 vccd1 vccd1 _5097_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1857 hold1857/A vssd1 vssd1 vccd1 vccd1 _5727_/D sky130_fd_sc_hd__buf_2
X_4117_ _4210_/A _4210_/B _5743_/Q vssd1 vssd1 vccd1 vccd1 _4169_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4048_ _4254_/B _4254_/C vssd1 vssd1 vccd1 vccd1 _4048_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput290 _5861_/X vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_12
X_4868__453 _5252_/CLK vssd1 vssd1 vccd1 vccd1 _5589_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__buf_2
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4453__38 _4453__38/A vssd1 vssd1 vccd1 vccd1 _5047_/CLK sky130_fd_sc_hd__inv_2
X_4909__494 _4909__494/A vssd1 vssd1 vccd1 vccd1 _5630_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3350_ _3350_/A _3350_/B vssd1 vssd1 vccd1 vccd1 _3351_/C sky130_fd_sc_hd__nand2_1
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5020_ _5022_/CLK _5020_/D vssd1 vssd1 vccd1 vccd1 _5020_/Q sky130_fd_sc_hd__dfxtp_1
X_3281_ _5482_/Q _5490_/Q _3281_/S vssd1 vssd1 vccd1 vccd1 _3281_/X sky130_fd_sc_hd__mux2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5922_ _5922_/A vssd1 vssd1 vccd1 vccd1 _5922_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4661__246 _4439__24/A vssd1 vssd1 vccd1 vccd1 _5349_/CLK sky130_fd_sc_hd__inv_2
X_5853_ _5853_/A vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _5451_/Q _5569_/Q _3024_/S vssd1 vssd1 vccd1 vccd1 _2996_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4702__287 _5002_/CLK vssd1 vssd1 vccd1 vccd1 _5393_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3617_ _4389_/B _3617_/B vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__nand2_1
X_3548_ _5118_/Q _3593_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5118_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold954 hold954/A vssd1 vssd1 vccd1 vccd1 hold954/X sky130_fd_sc_hd__buf_2
XFILLER_142_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4555__140 _4419__4/A vssd1 vssd1 vccd1 vccd1 _5197_/CLK sky130_fd_sc_hd__inv_2
Xhold965 hold965/A vssd1 vssd1 vccd1 vccd1 hold965/X sky130_fd_sc_hd__buf_2
Xhold998 hold998/A vssd1 vssd1 vccd1 vccd1 hold998/X sky130_fd_sc_hd__buf_2
Xhold987 hold987/A vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__buf_2
Xhold976 hold976/A vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__buf_2
X_3479_ _3614_/A1 _5179_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5179_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2322 hold2322/A vssd1 vssd1 vccd1 vccd1 hold2322/X sky130_fd_sc_hd__buf_2
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5218_ _5218_/CLK _5218_/D vssd1 vssd1 vccd1 vccd1 _5218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2355 hold2355/A vssd1 vssd1 vccd1 vccd1 hold766/A sky130_fd_sc_hd__buf_2
Xhold2344 hold2344/A vssd1 vssd1 vccd1 vccd1 hold2344/X sky130_fd_sc_hd__buf_2
Xhold1610 hold2452/X vssd1 vssd1 vccd1 vccd1 hold2453/A sky130_fd_sc_hd__buf_2
Xhold2333 hold2333/A vssd1 vssd1 vccd1 vccd1 hold993/A sky130_fd_sc_hd__buf_2
X_5149_ _5149_/CLK _5149_/D vssd1 vssd1 vccd1 vccd1 _5149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1621 hold2797/X vssd1 vssd1 vccd1 vccd1 hold2798/A sky130_fd_sc_hd__buf_2
Xhold1643 hold1643/A vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__buf_2
Xhold2388 hold985/X vssd1 vssd1 vccd1 vccd1 hold2388/X sky130_fd_sc_hd__buf_2
Xhold2366 hold2366/A vssd1 vssd1 vccd1 vccd1 hold2366/X sky130_fd_sc_hd__buf_2
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1676 hold2354/X vssd1 vssd1 vccd1 vccd1 hold2355/A sky130_fd_sc_hd__buf_2
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2850_ _5394_/Q _2850_/A1 _2851_/S vssd1 vssd1 vccd1 vccd1 _5394_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2781_ _5455_/Q _3600_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5455_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 hold227/X vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__buf_2
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__buf_2
X_4539__124 _4419__4/A vssd1 vssd1 vccd1 vccd1 _5181_/CLK sky130_fd_sc_hd__inv_2
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__buf_2
XCaravelHost_679 vssd1 vssd1 vccd1 vccd1 CaravelHost_679/HI la_data_out[107] sky130_fd_sc_hd__conb_1
XCaravelHost_668 vssd1 vssd1 vccd1 vccd1 CaravelHost_668/HI core1Index[6] sky130_fd_sc_hd__conb_1
X_3402_ _5277_/Q _3402_/A1 _3405_/S vssd1 vssd1 vccd1 vccd1 _5277_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_657 vssd1 vssd1 vccd1 vccd1 CaravelHost_657/HI core0Index[2] sky130_fd_sc_hd__conb_1
XFILLER_131_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4382_ _3644_/A _4389_/B _4398_/A2 vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__a21bo_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3328_/X _3329_/X _3332_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3333_/X sky130_fd_sc_hd__a211o_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3264_ _2464_/A _5303_/Q _5052_/Q _3128_/B _3326_/C1 vssd1 vssd1 vccd1 vccd1 _3264_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5004_/CLK _5003_/D vssd1 vssd1 vccd1 vccd1 _5003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3326_/C1 _3192_/X _3194_/X vssd1 vssd1 vccd1 vccd1 _3195_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5905_ _5905_/A vssd1 vssd1 vccd1 vccd1 _5905_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2979_ _2460_/A _5358_/Q _5125_/Q _3073_/B2 _3073_/C1 vssd1 vssd1 vccd1 vccd1 _2979_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5698_ _5751_/CLK _5698_/D vssd1 vssd1 vccd1 vccd1 _5698_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold740 hold740/A vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__buf_2
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2130 hold2130/A vssd1 vssd1 vccd1 vccd1 hold494/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_89_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4453__38/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2163 _3080_/B1 vssd1 vssd1 vccd1 vccd1 hold2163/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5730_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2152 _3859_/X vssd1 vssd1 vccd1 vccd1 hold2152/X sky130_fd_sc_hd__buf_2
XFILLER_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1451 _3961_/Y vssd1 vssd1 vccd1 vccd1 hold416/A sky130_fd_sc_hd__buf_2
Xhold2185 hold2185/A vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__buf_2
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2174 hold2793/X vssd1 vssd1 vccd1 vccd1 hold2794/A sky130_fd_sc_hd__buf_2
Xhold2196 hold2196/A vssd1 vssd1 vccd1 vccd1 hold2196/X sky130_fd_sc_hd__buf_2
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1495 hold970/X vssd1 vssd1 vccd1 vccd1 _3936_/A0 sky130_fd_sc_hd__buf_2
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1462 hold2887/X vssd1 vssd1 vccd1 vccd1 hold2888/A sky130_fd_sc_hd__buf_2
Xhold1473 hold959/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__buf_2
Xhold1484 _3935_/X vssd1 vssd1 vccd1 vccd1 hold965/A sky130_fd_sc_hd__buf_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xsplit1 split1/A vssd1 vssd1 vccd1 vccd1 split1/X sky130_fd_sc_hd__buf_4
XFILLER_0_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3951_ _5255_/Q _5108_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _5108_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2902_ _5032_/Q _5176_/Q _5240_/Q _5224_/Q _2944_/S0 _3040_/S vssd1 vssd1 vccd1 vccd1
+ _2902_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3882_ _4401_/A _5207_/Q _3882_/A3 _3855_/X vssd1 vssd1 vccd1 vccd1 _3882_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5621_ _5621_/CLK _5621_/D vssd1 vssd1 vccd1 vccd1 _5621_/Q sky130_fd_sc_hd__dfxtp_1
X_2833_ _5692_/Q _5409_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5409_/D sky130_fd_sc_hd__mux2_1
X_5552_ _5553_/CLK _5552_/D vssd1 vssd1 vccd1 vccd1 _5552_/Q sky130_fd_sc_hd__dfxtp_2
X_2764_ _5694_/Q _5467_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5467_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2695_ _5528_/Q _3572_/A0 _2702_/S vssd1 vssd1 vccd1 vccd1 _5528_/D sky130_fd_sc_hd__mux2_1
X_5483_ _5483_/CLK _5483_/D vssd1 vssd1 vccd1 vccd1 _5483_/Q sky130_fd_sc_hd__dfxtp_1
X_4773__358 _5697_/CLK vssd1 vssd1 vccd1 vccd1 _5464_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout505 _3777_/A3 vssd1 vssd1 vccd1 vccd1 _3774_/C1 sky130_fd_sc_hd__buf_6
X_4365_ _4365_/A _5725_/Q vssd1 vssd1 vccd1 vccd1 _5731_/D sky130_fd_sc_hd__and2_1
Xfanout516 _2867_/B vssd1 vssd1 vccd1 vccd1 _2943_/S1 sky130_fd_sc_hd__buf_4
Xfanout527 _3002_/S vssd1 vssd1 vccd1 vccd1 _3069_/S sky130_fd_sc_hd__buf_6
XFILLER_101_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _5615_/Q _2464_/A _3128_/B _5607_/Q _3316_/C1 vssd1 vssd1 vccd1 vccd1 _3316_/X
+ sky130_fd_sc_hd__o221a_1
X_4814__399 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5505_/CLK sky130_fd_sc_hd__inv_2
Xfanout538 _3299_/S vssd1 vssd1 vccd1 vccd1 _3330_/S sky130_fd_sc_hd__buf_6
X_4489__74 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5131_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4296_ _4261_/B _4308_/A2 _4308_/B1 _2450_/Y vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__o22a_1
Xfanout549 _4282_/Y vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _5483_/Q _5491_/Q _3281_/S vssd1 vssd1 vccd1 vccd1 _3247_/X sky130_fd_sc_hd__mux2_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3178_ _3136_/X _3164_/X _3168_/X _3177_/X vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__a31o_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4667__252 _5084_/CLK vssd1 vssd1 vccd1 vccd1 _5355_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4708__293 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5399_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold570 hold822/X vssd1 vssd1 vccd1 vccd1 hold823/A sky130_fd_sc_hd__buf_2
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2480_ _5334_/Q _5329_/Q vssd1 vssd1 vccd1 vccd1 _3123_/B sky130_fd_sc_hd__xor2_1
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ _5552_/Q _4210_/A _5553_/Q vssd1 vssd1 vccd1 vccd1 _4153_/C sky130_fd_sc_hd__a21o_1
X_3101_ _3066_/S _3099_/A _2778_/A vssd1 vssd1 vccd1 vccd1 _3101_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4081_ _4081_/A _4081_/B _4279_/B vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__and3_2
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3032_ _3074_/A1 _3030_/X _3031_/X _3097_/B vssd1 vssd1 vccd1 vccd1 _3032_/X sky130_fd_sc_hd__o211a_1
Xinput190 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__buf_6
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _5016_/CLK _4983_/D vssd1 vssd1 vccd1 vccd1 _4983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3934_ _3934_/A0 _5091_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3865_ _5067_/Q _3959_/A _3865_/B1 vssd1 vssd1 vccd1 vccd1 _3865_/X sky130_fd_sc_hd__a21o_1
X_5604_ _5604_/CLK _5604_/D vssd1 vssd1 vccd1 vccd1 _5604_/Q sky130_fd_sc_hd__dfxtp_1
X_2816_ _3370_/A _2852_/A vssd1 vssd1 vccd1 vccd1 _2824_/S sky130_fd_sc_hd__or2_4
XFILLER_118_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3796_ hold137/X _5247_/Q _3796_/A3 _3796_/B1 _4996_/Q vssd1 vssd1 vccd1 vccd1 _3796_/X
+ sky130_fd_sc_hd__o32a_1
X_5535_ _5535_/CLK _5535_/D vssd1 vssd1 vccd1 vccd1 _5535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2747_ _3308_/A1 _5482_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5482_/D sky130_fd_sc_hd__mux2_1
X_2678_ _3602_/A1 _5571_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5571_/D sky130_fd_sc_hd__mux2_1
X_5466_ _5466_/CLK _5466_/D vssd1 vssd1 vccd1 vccd1 _5466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5397_ _5397_/CLK _5397_/D vssd1 vssd1 vccd1 vccd1 _5397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4348_ _5691_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4348_/X sky130_fd_sc_hd__or2_1
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4279_ _4324_/A _4279_/B vssd1 vssd1 vccd1 vccd1 _4279_/X sky130_fd_sc_hd__or2_1
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4795__380 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5486_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4507__92/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _3650_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__or2_1
XFILLER_127_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3581_ _3599_/A1 _5041_/Q _3588_/S vssd1 vssd1 vccd1 vccd1 _5041_/D sky130_fd_sc_hd__mux2_1
X_2601_ _3567_/A1 _5618_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5618_/D sky130_fd_sc_hd__mux2_1
X_5320_ _5684_/CLK _5320_/D vssd1 vssd1 vccd1 vccd1 _5320_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2532_ _5693_/Q _5709_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5709_/D sky130_fd_sc_hd__mux2_1
X_5251_ _5252_/CLK _5251_/D vssd1 vssd1 vccd1 vccd1 _5251_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4202_ _4204_/A _4202_/B vssd1 vssd1 vccd1 vccd1 _5547_/D sky130_fd_sc_hd__nor2_1
X_2463_ _5329_/Q vssd1 vssd1 vccd1 vccd1 _2463_/Y sky130_fd_sc_hd__inv_2
X_5182_ _5182_/CLK _5182_/D vssd1 vssd1 vccd1 vccd1 _5182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2707 hold2707/A vssd1 vssd1 vccd1 vccd1 hold2707/X sky130_fd_sc_hd__buf_2
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4133_ _5751_/Q _4133_/B vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__xor2_1
X_4459__44 _4459__44/A vssd1 vssd1 vccd1 vccd1 _5053_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4064_ _5752_/Q _4261_/B vssd1 vssd1 vccd1 vccd1 _4275_/C sky130_fd_sc_hd__xor2_2
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3015_ _3094_/B _3011_/X _3012_/X _3014_/X vssd1 vssd1 vccd1 vccd1 _3015_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ _5684_/CLK _4966_/D vssd1 vssd1 vccd1 vccd1 _4966_/Q sky130_fd_sc_hd__dfxtp_2
X_3917_ _5082_/Q _3926_/A2 _3923_/B1 _3916_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5082_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3848_ _5090_/Q _3850_/C _2501_/X vssd1 vssd1 vccd1 vccd1 _4369_/D sky130_fd_sc_hd__o21a_1
X_4779__364 _5019_/CLK vssd1 vssd1 vccd1 vccd1 _5470_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3779_ _5023_/Q _5024_/Q vssd1 vssd1 vccd1 vccd1 _3779_/Y sky130_fd_sc_hd__nand2b_1
X_5518_ _5518_/CLK _5518_/D vssd1 vssd1 vccd1 vccd1 _5518_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5449_ _5449_/CLK _5449_/D vssd1 vssd1 vccd1 vccd1 _5449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4572__157 _5111_/CLK vssd1 vssd1 vccd1 vccd1 _5222_/CLK sky130_fd_sc_hd__inv_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4613__198 _5019_/CLK vssd1 vssd1 vccd1 vccd1 _5287_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3702_ _4987_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3702_/X sky130_fd_sc_hd__or2_1
X_3633_ _4354_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__or2_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3564_ _5056_/Q _3564_/A1 _3570_/S vssd1 vssd1 vccd1 vccd1 _5056_/D sky130_fd_sc_hd__mux2_1
X_3495_ _3594_/A1 _5165_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5165_/D sky130_fd_sc_hd__mux2_1
X_5303_ _5303_/CLK _5303_/D vssd1 vssd1 vccd1 vccd1 _5303_/Q sky130_fd_sc_hd__dfxtp_1
X_2515_ _3406_/A _3562_/A vssd1 vssd1 vccd1 vccd1 _2523_/S sky130_fd_sc_hd__or2_4
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2504 hold2504/A vssd1 vssd1 vccd1 vccd1 _5320_/D sky130_fd_sc_hd__buf_2
X_5234_ _5234_/CLK _5234_/D vssd1 vssd1 vccd1 vccd1 _5234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2446_ _5672_/Q vssd1 vssd1 vccd1 vccd1 _2446_/Y sky130_fd_sc_hd__inv_2
X_5165_ _5165_/CLK _5165_/D vssd1 vssd1 vccd1 vccd1 _5165_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2537 hold2537/A vssd1 vssd1 vccd1 vccd1 hold2537/X sky130_fd_sc_hd__buf_2
Xhold2526 hold2526/A vssd1 vssd1 vccd1 vccd1 hold833/A sky130_fd_sc_hd__buf_2
Xhold2515 hold2515/A vssd1 vssd1 vccd1 vccd1 hold2515/X sky130_fd_sc_hd__buf_2
Xhold1814 hold2574/X vssd1 vssd1 vccd1 vccd1 hold2575/A sky130_fd_sc_hd__buf_2
Xhold1825 hold1825/A vssd1 vssd1 vccd1 vccd1 hold728/A sky130_fd_sc_hd__buf_2
Xhold1836 _3828_/X vssd1 vssd1 vccd1 vccd1 hold1836/X sky130_fd_sc_hd__buf_2
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4116_ _5743_/Q _4210_/A _4210_/B vssd1 vssd1 vccd1 vccd1 _4118_/C sky130_fd_sc_hd__or3_1
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1847 _4378_/X vssd1 vssd1 vccd1 vccd1 hold1847/X sky130_fd_sc_hd__buf_2
X_5096_ _5542_/CLK _5096_/D vssd1 vssd1 vccd1 vccd1 _5096_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1858 wbs_we_i vssd1 vssd1 vccd1 vccd1 hold1858/X sky130_fd_sc_hd__buf_2
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4047_ _5669_/Q _4065_/B _5670_/Q vssd1 vssd1 vccd1 vccd1 _4254_/C sky130_fd_sc_hd__a21o_2
XFILLER_72_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput280 _5852_/X vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_12
XFILLER_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput291 _5862_/X vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_12
XFILLER_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3280_ _3328_/A _3278_/X _3279_/X vssd1 vssd1 vccd1 vccd1 _3280_/X sky130_fd_sc_hd__o21a_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4429__14 _4424__9/A vssd1 vssd1 vccd1 vccd1 _4980_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _5921_/A vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5852_ _5852_/A vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2995_ _5060_/Q _3031_/B1 _3029_/B1 _2994_/X vssd1 vssd1 vccd1 vccd1 _2995_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3616_ _5264_/Q _5265_/Q _5262_/Q _5263_/Q vssd1 vssd1 vccd1 vccd1 _3617_/B sky130_fd_sc_hd__and4bb_4
X_3547_ _5119_/Q _3592_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5119_/D sky130_fd_sc_hd__mux2_1
Xhold955 hold955/A vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__buf_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold988 hold988/A vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__buf_2
Xhold977 hold977/A vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__buf_2
Xhold966 hold966/A vssd1 vssd1 vccd1 vccd1 hold966/X sky130_fd_sc_hd__buf_2
X_3478_ _3613_/A1 _5180_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5180_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold999 hold999/A vssd1 vssd1 vccd1 vccd1 hold999/X sky130_fd_sc_hd__buf_2
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5217_ _5217_/CLK _5217_/D vssd1 vssd1 vccd1 vccd1 _5217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2345 hold2345/A vssd1 vssd1 vccd1 vccd1 hold2345/X sky130_fd_sc_hd__buf_2
Xhold1600 hold2465/X vssd1 vssd1 vccd1 vccd1 hold1600/X sky130_fd_sc_hd__buf_2
Xhold2323 hold2323/A vssd1 vssd1 vccd1 vccd1 _5695_/D sky130_fd_sc_hd__buf_2
X_5148_ _5148_/CLK _5148_/D vssd1 vssd1 vccd1 vccd1 _5148_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1644 hold2590/X vssd1 vssd1 vccd1 vccd1 hold2591/A sky130_fd_sc_hd__buf_2
Xhold2378 _4406_/X vssd1 vssd1 vccd1 vccd1 hold2378/X sky130_fd_sc_hd__buf_2
Xhold1622 hold2801/X vssd1 vssd1 vccd1 vccd1 hold2185/A sky130_fd_sc_hd__buf_2
Xhold2356 hold766/X vssd1 vssd1 vccd1 vccd1 hold2356/X sky130_fd_sc_hd__buf_2
Xhold1611 hold2454/X vssd1 vssd1 vccd1 vccd1 hold2455/A sky130_fd_sc_hd__buf_2
Xhold2389 hold2389/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__buf_2
Xhold2367 hold2367/A vssd1 vssd1 vccd1 vccd1 hold2367/X sky130_fd_sc_hd__buf_2
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5742_/CLK _5079_/D vssd1 vssd1 vccd1 vccd1 _5079_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1677 hold2356/X vssd1 vssd1 vccd1 vccd1 hold2357/A sky130_fd_sc_hd__buf_2
XFILLER_45_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1666 hold2316/X vssd1 vssd1 vccd1 vccd1 hold2317/A sky130_fd_sc_hd__buf_2
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4941__526 _4941__526/A vssd1 vssd1 vccd1 vccd1 _5662_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4835__420 _5683_/CLK vssd1 vssd1 vccd1 vccd1 _5526_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4513__98 _5684_/CLK vssd1 vssd1 vccd1 vccd1 _5155_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2890 hold2906/X vssd1 vssd1 vccd1 vccd1 hold2907/A sky130_fd_sc_hd__buf_2
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4684__269 _4425__10/A vssd1 vssd1 vccd1 vccd1 _5373_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2780_ _5456_/Q _3599_/A1 _2787_/S vssd1 vssd1 vccd1 vccd1 _5456_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4578__163 _4510__95/A vssd1 vssd1 vccd1 vccd1 _5228_/CLK sky130_fd_sc_hd__inv_2
Xhold218 hold229/X vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__buf_2
Xhold229 _3989_/X vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__buf_2
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4381_ _5291_/Q _4381_/B vssd1 vssd1 vccd1 vccd1 _4381_/X sky130_fd_sc_hd__and2_1
X_3401_ _5278_/Q _3575_/A0 _3405_/S vssd1 vssd1 vccd1 vccd1 _5278_/D sky130_fd_sc_hd__mux2_1
XCaravelHost_669 vssd1 vssd1 vccd1 vccd1 CaravelHost_669/HI core1Index[7] sky130_fd_sc_hd__conb_1
XCaravelHost_658 vssd1 vssd1 vccd1 vccd1 CaravelHost_658/HI core0Index[3] sky130_fd_sc_hd__conb_1
X_3332_ _3328_/A _3330_/X _3331_/X _3171_/A vssd1 vssd1 vccd1 vccd1 _3332_/X sky130_fd_sc_hd__o211a_1
XFILLER_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3263_ _3357_/B _3263_/B vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__or2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/CLK _5002_/D vssd1 vssd1 vccd1 vccd1 _5002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3194_ _3320_/C1 _3193_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3194_/X sky130_fd_sc_hd__a21o_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5904_ _5904_/A vssd1 vssd1 vccd1 vccd1 _5904_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2978_ _3034_/A _2978_/B vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__or2_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5697_ _5697_/CLK _5697_/D vssd1 vssd1 vccd1 vccd1 _5697_/Q sky130_fd_sc_hd__dfxtp_1
X_4819__404 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_147_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap460 _4401_/B vssd1 vssd1 vccd1 vccd1 _4381_/B sky130_fd_sc_hd__buf_2
Xhold741 hold741/A vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__buf_2
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold774 hold774/A vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__buf_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2120 _3870_/X vssd1 vssd1 vccd1 vccd1 hold2120/X sky130_fd_sc_hd__buf_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2164 hold2164/A vssd1 vssd1 vccd1 vccd1 hold953/A sky130_fd_sc_hd__buf_2
Xhold2153 hold2153/A vssd1 vssd1 vccd1 vccd1 hold560/A sky130_fd_sc_hd__buf_2
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1452 hold416/X vssd1 vssd1 vccd1 vccd1 _5113_/D sky130_fd_sc_hd__buf_2
Xhold2186 hold61/X vssd1 vssd1 vccd1 vccd1 hold2186/X sky130_fd_sc_hd__buf_2
XFILLER_18_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2197 hold2197/A vssd1 vssd1 vccd1 vccd1 hold2197/X sky130_fd_sc_hd__buf_2
Xhold1474 hold14/X vssd1 vssd1 vccd1 vccd1 hold960/A sky130_fd_sc_hd__buf_2
Xhold1485 hold965/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__buf_2
Xhold1463 hold2792/X vssd1 vssd1 vccd1 vccd1 hold2793/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_58_wb_clk_i _5025_/CLK vssd1 vssd1 vccd1 vccd1 _5006_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1496 _3936_/X vssd1 vssd1 vccd1 vccd1 hold971/A sky130_fd_sc_hd__buf_2
XFILLER_26_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xsplit2 split2/A vssd1 vssd1 vccd1 vccd1 split2/X sky130_fd_sc_hd__buf_4
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__buf_2
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3950_ _5254_/Q _5107_/Q _3953_/S vssd1 vssd1 vccd1 vccd1 _3950_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2901_ _5200_/Q _5184_/Q _4973_/Q _5192_/Q _3036_/S _2943_/S1 vssd1 vssd1 vccd1 vccd1
+ _2901_/X sky130_fd_sc_hd__mux4_2
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3881_ _5750_/Q _3998_/A1 _3882_/A3 _3887_/A vssd1 vssd1 vccd1 vccd1 _3881_/X sky130_fd_sc_hd__a31o_1
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5620_ _5620_/CLK _5620_/D vssd1 vssd1 vccd1 vccd1 _5620_/Q sky130_fd_sc_hd__dfxtp_1
X_2832_ _5693_/Q _5410_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5410_/D sky130_fd_sc_hd__mux2_1
X_5551_ _5551_/CLK _5551_/D vssd1 vssd1 vccd1 vccd1 _5551_/Q sky130_fd_sc_hd__dfxtp_2
X_2763_ _3393_/A0 _5468_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5468_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5482_ _5482_/CLK _5482_/D vssd1 vssd1 vccd1 vccd1 _5482_/Q sky130_fd_sc_hd__dfxtp_1
X_2694_ _3571_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _2702_/S sky130_fd_sc_hd__nor2_8
XFILLER_145_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4364_ _4365_/A _5724_/Q vssd1 vssd1 vccd1 vccd1 _5730_/D sky130_fd_sc_hd__and2_1
Xfanout506 _2497_/Y vssd1 vssd1 vccd1 vccd1 _3777_/A3 sky130_fd_sc_hd__buf_12
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout528 _5364_/Q vssd1 vssd1 vccd1 vccd1 _3002_/S sky130_fd_sc_hd__buf_6
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout517 _5365_/Q vssd1 vssd1 vccd1 vccd1 _2867_/B sky130_fd_sc_hd__buf_12
X_4295_ _4294_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5667_/D sky130_fd_sc_hd__and2b_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3315_ _5575_/Q _5591_/Q _3318_/S vssd1 vssd1 vccd1 vccd1 _3315_/X sky130_fd_sc_hd__mux2_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout539 _3327_/S vssd1 vssd1 vccd1 vccd1 _3299_/S sky130_fd_sc_hd__buf_6
XFILLER_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3246_ _3567_/A1 _3159_/B _3245_/X _3277_/C1 vssd1 vssd1 vccd1 vccd1 _5340_/D sky130_fd_sc_hd__o211a_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3177_ _3171_/X _3173_/X _3176_/X _3334_/A1 _3169_/B vssd1 vssd1 vccd1 vccd1 _3177_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5749_ _5751_/CLK _5749_/D vssd1 vssd1 vccd1 vccd1 _5749_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_105_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5566_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_135_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold560 hold560/A vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__buf_2
Xhold571 hold826/X vssd1 vssd1 vccd1 vccd1 hold690/A sky130_fd_sc_hd__buf_2
XFILLER_104_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4947__532 _4965__550/A vssd1 vssd1 vccd1 vccd1 _5705_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1293 hold2573/X vssd1 vssd1 vccd1 vccd1 hold2574/A sky130_fd_sc_hd__buf_2
Xhold1282 hold2511/X vssd1 vssd1 vccd1 vccd1 hold2512/A sky130_fd_sc_hd__buf_2
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3100_ _2867_/B _3099_/A _3099_/Y _2778_/A vssd1 vssd1 vccd1 vccd1 _5365_/D sky130_fd_sc_hd__o211a_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4080_ _4080_/A _4080_/B vssd1 vssd1 vccd1 vccd1 _4279_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3031_ _5434_/Q _2460_/Y _3031_/B1 _5426_/Q vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__o22a_1
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput180 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput191 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__buf_4
X_4982_ _4982_/CLK _4982_/D vssd1 vssd1 vccd1 vccd1 _4982_/Q sky130_fd_sc_hd__dfxtp_1
X_4740__325 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5431_/CLK sky130_fd_sc_hd__inv_2
X_3933_ _3933_/A0 _5090_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3933_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5734_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3864_ _4399_/B _3861_/X _3863_/X _4361_/A vssd1 vssd1 vccd1 vccd1 _3864_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5603_ _5603_/CLK _5603_/D vssd1 vssd1 vccd1 vccd1 _5603_/Q sky130_fd_sc_hd__dfxtp_1
X_2815_ _3543_/A0 _5425_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5425_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3795_ hold137/X _5246_/Q _3796_/A3 _3795_/B1 _4995_/Q vssd1 vssd1 vccd1 vccd1 _3795_/X
+ sky130_fd_sc_hd__o32a_1
X_5534_ _5534_/CLK _5534_/D vssd1 vssd1 vccd1 vccd1 _5534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2746_ _3277_/A1 _5483_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5483_/D sky130_fd_sc_hd__mux2_1
X_2677_ _3601_/A1 _5572_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5572_/D sky130_fd_sc_hd__mux2_1
X_5465_ _5465_/CLK _5465_/D vssd1 vssd1 vccd1 vccd1 _5465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4416_ _5755_/Q _4401_/Y _4415_/X vssd1 vssd1 vccd1 vccd1 _4416_/X sky130_fd_sc_hd__a21o_1
X_5396_ _5396_/CLK _5396_/D vssd1 vssd1 vccd1 vccd1 _5396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4347_ _5691_/Q _4324_/X _4346_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _5690_/D sky130_fd_sc_hd__o211a_1
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4278_ _4081_/A _4324_/A _4269_/A _4269_/B vssd1 vssd1 vccd1 vccd1 _4278_/X sky130_fd_sc_hd__o22a_2
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3229_ _3357_/B _3227_/X _3228_/X vssd1 vssd1 vccd1 vccd1 _3242_/B sky130_fd_sc_hd__o21a_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5557_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4724__309 _5244_/CLK vssd1 vssd1 vccd1 vccd1 _5415_/CLK sky130_fd_sc_hd__inv_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3580_ _3598_/B _3607_/A vssd1 vssd1 vccd1 vccd1 _3588_/S sky130_fd_sc_hd__or2_4
XFILLER_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2600_ _3575_/A0 _5619_/Q _2604_/S vssd1 vssd1 vccd1 vccd1 _5619_/D sky130_fd_sc_hd__mux2_1
X_4618__203 _4960__545/A vssd1 vssd1 vccd1 vccd1 _5295_/CLK sky130_fd_sc_hd__inv_2
X_2531_ _3394_/A0 _5710_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5710_/D sky130_fd_sc_hd__mux2_1
X_5250_ _5252_/CLK _5250_/D vssd1 vssd1 vccd1 vccd1 _5250_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4201_ _5547_/Q _4187_/B1 _4210_/C _4121_/Y vssd1 vssd1 vccd1 vccd1 _4202_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2462_ _5331_/Q vssd1 vssd1 vccd1 vccd1 _3350_/A sky130_fd_sc_hd__inv_2
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5181_ _5181_/CLK _5181_/D vssd1 vssd1 vccd1 vccd1 _5181_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2708 hold2708/A vssd1 vssd1 vccd1 vccd1 hold2708/X sky130_fd_sc_hd__buf_2
XFILLER_110_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4132_ _5543_/Q _4132_/B vssd1 vssd1 vccd1 vccd1 _4133_/B sky130_fd_sc_hd__xnor2_2
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4063_ _4063_/A _4063_/B vssd1 vssd1 vccd1 vccd1 _4261_/B sky130_fd_sc_hd__nand2_2
XFILLER_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3014_ _3045_/A1 _2995_/X _2998_/X _3013_/X _2883_/X vssd1 vssd1 vccd1 vccd1 _3014_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4474__59 _4510__95/A vssd1 vssd1 vccd1 vccd1 _5116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3916_ _5739_/Q _3924_/B _5292_/Q vssd1 vssd1 vccd1 vccd1 _3916_/X sky130_fd_sc_hd__and3_1
XFILLER_51_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3847_ _5755_/Q _3998_/A1 _3882_/A3 _3887_/A vssd1 vssd1 vccd1 vccd1 _3847_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _3778_/A _3778_/B _3778_/C vssd1 vssd1 vccd1 vccd1 _3778_/X sky130_fd_sc_hd__and3_1
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5517_ _5517_/CLK _5517_/D vssd1 vssd1 vccd1 vccd1 _5517_/Q sky130_fd_sc_hd__dfxtp_1
X_2729_ _3308_/A1 _5498_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5498_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5448_ _5448_/CLK _5448_/D vssd1 vssd1 vccd1 vccd1 _5448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5379_ _5379_/CLK _5379_/D vssd1 vssd1 vccd1 vccd1 _5379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5022_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3701_ _5070_/Q input29/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3701_/X sky130_fd_sc_hd__mux2_4
XFILLER_147_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3632_ _4353_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3632_/X sky130_fd_sc_hd__or2_1
XFILLER_128_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4852__437 _5252_/CLK vssd1 vssd1 vccd1 vccd1 _5573_/CLK sky130_fd_sc_hd__inv_2
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3563_ _5057_/Q _3572_/A0 _3570_/S vssd1 vssd1 vccd1 vccd1 _5057_/D sky130_fd_sc_hd__mux2_1
X_5302_ _5302_/CLK _5302_/D vssd1 vssd1 vccd1 vccd1 _5302_/Q sky130_fd_sc_hd__dfxtp_1
X_3494_ _3593_/A1 _5166_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5166_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2514_ _5332_/Q _3350_/A _3350_/B split3/A vssd1 vssd1 vccd1 vccd1 _3562_/A sky130_fd_sc_hd__or4b_4
X_5233_ _5233_/CLK _5233_/D vssd1 vssd1 vccd1 vccd1 _5233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2445_ _5673_/Q vssd1 vssd1 vccd1 vccd1 _2445_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5164_ _5164_/CLK _5164_/D vssd1 vssd1 vccd1 vccd1 _5164_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2538 hold2538/A vssd1 vssd1 vccd1 vccd1 hold2538/X sky130_fd_sc_hd__buf_2
Xhold2527 hold833/X vssd1 vssd1 vccd1 vccd1 hold2527/X sky130_fd_sc_hd__buf_2
Xhold2516 hold2516/A vssd1 vssd1 vccd1 vccd1 hold2516/X sky130_fd_sc_hd__buf_2
Xhold1826 hold728/X vssd1 vssd1 vccd1 vccd1 hold1826/X sky130_fd_sc_hd__buf_2
Xhold1815 hold2576/X vssd1 vssd1 vccd1 vccd1 hold2577/A sky130_fd_sc_hd__buf_2
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2549 hold2875/X vssd1 vssd1 vccd1 vccd1 hold2549/X sky130_fd_sc_hd__buf_2
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4115_ _4108_/B _4119_/C _4104_/D _5551_/Q vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__a31oi_4
Xhold1848 hold1848/A vssd1 vssd1 vccd1 vccd1 hold787/A sky130_fd_sc_hd__buf_2
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1837 hold1837/A vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__buf_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5095_ _5542_/CLK _5095_/D vssd1 vssd1 vccd1 vccd1 _5095_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1859 hold1859/A vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__buf_2
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4046_ _5749_/Q _4046_/B _4046_/C vssd1 vssd1 vccd1 vccd1 _4271_/B sky130_fd_sc_hd__nand3b_1
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4746__331 _4746__331/A vssd1 vssd1 vccd1 vccd1 _5437_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput270 _3627_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput281 _5853_/X vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_12
Xoutput292 _5863_/X vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_12
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4444__29 _4468__53/A vssd1 vssd1 vccd1 vccd1 _5038_/CLK sky130_fd_sc_hd__inv_2
X_5920_ _5920_/A vssd1 vssd1 vccd1 vccd1 _5920_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5851_ _5851_/A vssd1 vssd1 vccd1 vccd1 _5851_/X sky130_fd_sc_hd__clkbuf_4
X_2994_ _4977_/Q _2870_/B _2993_/X _3034_/A vssd1 vssd1 vccd1 vccd1 _2994_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3615_ _4967_/Q _3615_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4967_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3546_ _5120_/Q _3591_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5120_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold989 hold989/A vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__buf_2
Xhold978 hold978/A vssd1 vssd1 vccd1 vccd1 hold978/X sky130_fd_sc_hd__buf_2
Xhold967 hold967/A vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__buf_2
Xhold956 hold956/A vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__buf_2
X_3477_ _3612_/A1 _5181_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5181_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5216_ _5216_/CLK _5216_/D vssd1 vssd1 vccd1 vccd1 _5216_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2346 hold2346/A vssd1 vssd1 vccd1 vccd1 _5696_/D sky130_fd_sc_hd__buf_2
Xhold2324 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 hold2324/X sky130_fd_sc_hd__buf_2
Xhold1601 hold1601/A vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__buf_2
XFILLER_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5147_ _5147_/CLK _5147_/D vssd1 vssd1 vccd1 vccd1 _5147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1623 hold2186/X vssd1 vssd1 vccd1 vccd1 hold2187/A sky130_fd_sc_hd__buf_2
Xhold2357 hold2357/A vssd1 vssd1 vccd1 vccd1 hold2357/X sky130_fd_sc_hd__buf_2
Xhold2379 hold2379/A vssd1 vssd1 vccd1 vccd1 hold2379/X sky130_fd_sc_hd__buf_2
Xhold1612 hold2456/X vssd1 vssd1 vccd1 vccd1 hold1612/X sky130_fd_sc_hd__buf_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2368 hold2368/A vssd1 vssd1 vccd1 vccd1 hold754/A sky130_fd_sc_hd__buf_2
X_5078_ _5383_/CLK _5078_/D vssd1 vssd1 vccd1 vccd1 _5078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1645 hold2592/X vssd1 vssd1 vccd1 vccd1 hold2593/A sky130_fd_sc_hd__buf_2
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1678 hold2358/X vssd1 vssd1 vccd1 vccd1 hold2359/A sky130_fd_sc_hd__buf_2
Xhold1667 hold2318/X vssd1 vssd1 vccd1 vccd1 hold2319/A sky130_fd_sc_hd__buf_2
X_4029_ _5673_/Q _4065_/B _4029_/C vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__and3_2
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4523__108 _4435__20/A vssd1 vssd1 vccd1 vccd1 _5165_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold219 hold231/X vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__buf_2
X_4380_ _5739_/Q _4370_/X _4380_/B1 hold875/X vssd1 vssd1 vccd1 vccd1 _4380_/X sky130_fd_sc_hd__o211a_1
X_3400_ _5279_/Q _3574_/A0 _3405_/S vssd1 vssd1 vccd1 vccd1 _5279_/D sky130_fd_sc_hd__mux2_1
XCaravelHost_659 vssd1 vssd1 vccd1 vccd1 CaravelHost_659/HI core0Index[4] sky130_fd_sc_hd__conb_1
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3331_ _5473_/Q _3331_/A2 _3237_/B _5708_/Q vssd1 vssd1 vccd1 vccd1 _3331_/X sky130_fd_sc_hd__o22a_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3262_ _5523_/Q _5276_/Q _3324_/S vssd1 vssd1 vccd1 vccd1 _3263_/B sky130_fd_sc_hd__mux2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/CLK _5001_/D vssd1 vssd1 vccd1 vccd1 _5001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3193_ _5721_/Q _5298_/Q _5271_/Q _5705_/Q _3290_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3193_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4964__549 _4964__549/A vssd1 vssd1 vccd1 vccd1 _5722_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5903_ _5903_/A vssd1 vssd1 vccd1 vccd1 _5903_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2977_ _5157_/Q _5313_/Q _3002_/S vssd1 vssd1 vccd1 vccd1 _2978_/B sky130_fd_sc_hd__mux2_1
X_4858__443 _4898__483/A vssd1 vssd1 vccd1 vccd1 _5579_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5696_ _5734_/CLK _5696_/D vssd1 vssd1 vccd1 vccd1 _5696_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold742 hold742/A vssd1 vssd1 vccd1 vccd1 _4244_/S sky130_fd_sc_hd__buf_2
X_3529_ _5135_/Q _3610_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5135_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold786 hold786/A vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__buf_2
XFILLER_103_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2121 hold2121/A vssd1 vssd1 vccd1 vccd1 hold489/A sky130_fd_sc_hd__buf_2
Xhold2110 hold2110/A vssd1 vssd1 vccd1 vccd1 hold474/A sky130_fd_sc_hd__buf_2
XFILLER_130_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2154 hold560/X vssd1 vssd1 vccd1 vccd1 hold2154/X sky130_fd_sc_hd__buf_2
Xhold2143 _3884_/X vssd1 vssd1 vccd1 vccd1 hold2143/X sky130_fd_sc_hd__buf_2
XFILLER_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2165 hold953/X vssd1 vssd1 vccd1 vccd1 hold2165/X sky130_fd_sc_hd__buf_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2187 hold2187/A vssd1 vssd1 vccd1 vccd1 hold2187/X sky130_fd_sc_hd__buf_2
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1475 hold960/X vssd1 vssd1 vccd1 vccd1 _5091_/D sky130_fd_sc_hd__buf_2
Xhold1486 hold20/X vssd1 vssd1 vccd1 vccd1 hold966/A sky130_fd_sc_hd__buf_2
Xhold1464 hold2234/X vssd1 vssd1 vccd1 vccd1 hold2235/A sky130_fd_sc_hd__buf_2
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2198 hold2198/A vssd1 vssd1 vccd1 vccd1 _4997_/D sky130_fd_sc_hd__buf_2
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1497 hold971/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__buf_2
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_98_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4821__406/A
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_27_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4508__93/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4651__236 _4658__243/A vssd1 vssd1 vccd1 vccd1 _5337_/CLK sky130_fd_sc_hd__inv_2
XFILLER_122_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xsplit3 split3/A vssd1 vssd1 vccd1 vccd1 split3/X sky130_fd_sc_hd__buf_2
XFILLER_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__buf_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__buf_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4545__130 _4418__3/A vssd1 vssd1 vccd1 vccd1 _5187_/CLK sky130_fd_sc_hd__inv_2
X_2900_ _2898_/X _2899_/X _2947_/S vssd1 vssd1 vccd1 vccd1 _2900_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3880_ _5070_/Q _3959_/A hold526/X vssd1 vssd1 vccd1 vccd1 _3880_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2831_ _3394_/A0 _5411_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5411_/D sky130_fd_sc_hd__mux2_1
X_4422__7 _4422__7/A vssd1 vssd1 vccd1 vccd1 _4973_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _5551_/CLK _5550_/D vssd1 vssd1 vccd1 vccd1 _5550_/Q sky130_fd_sc_hd__dfxtp_1
X_2762_ _3392_/A0 _5469_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5469_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5481_ _5481_/CLK _5481_/D vssd1 vssd1 vccd1 vccd1 _5481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2693_ _5335_/Q _5334_/Q _3346_/A vssd1 vssd1 vccd1 vccd1 _3562_/B sky130_fd_sc_hd__nand3_4
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4363_ _4368_/A _5363_/Q vssd1 vssd1 vccd1 vccd1 _5729_/D sky130_fd_sc_hd__and2_1
Xfanout518 _5365_/Q vssd1 vssd1 vccd1 vccd1 _2941_/S0 sky130_fd_sc_hd__clkbuf_16
XFILLER_112_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4294_ _4058_/Y _4308_/A2 _4308_/B1 _2451_/Y vssd1 vssd1 vccd1 vccd1 _4294_/X sky130_fd_sc_hd__o22a_1
Xfanout507 _4369_/A vssd1 vssd1 vccd1 vccd1 _4399_/B sky130_fd_sc_hd__buf_4
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _3357_/B _3312_/X _3313_/X vssd1 vssd1 vccd1 vccd1 _3314_/X sky130_fd_sc_hd__o21a_1
Xfanout529 _5333_/Q vssd1 vssd1 vccd1 vccd1 _3346_/A sky130_fd_sc_hd__buf_6
XFILLER_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3245_ _5340_/Q _3125_/A _3156_/X _3244_/X vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__a211o_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3176_ _3174_/X _3175_/X _3240_/S vssd1 vssd1 vccd1 vccd1 _3176_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5748_ _5752_/CLK _5748_/D vssd1 vssd1 vccd1 vccd1 _5748_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ _5738_/CLK _5679_/D vssd1 vssd1 vccd1 vccd1 _5679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold561 hold561/A vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__buf_2
Xhold572 hold739/X vssd1 vssd1 vccd1 vccd1 hold740/A sky130_fd_sc_hd__buf_2
XFILLER_2_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold594 hold759/X vssd1 vssd1 vccd1 vccd1 hold760/A sky130_fd_sc_hd__buf_2
XFILLER_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1261 hold2485/X vssd1 vssd1 vccd1 vccd1 hold2486/A sky130_fd_sc_hd__buf_2
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1283 hold2515/X vssd1 vssd1 vccd1 vccd1 hold2516/A sky130_fd_sc_hd__buf_2
Xhold1294 hold2577/X vssd1 vssd1 vccd1 vccd1 hold2578/A sky130_fd_sc_hd__buf_2
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4529__114 _4435__20/A vssd1 vssd1 vccd1 vccd1 _5171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3030_ _5394_/Q _5402_/Q _3069_/S vssd1 vssd1 vccd1 vccd1 _3030_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput170 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__clkbuf_8
Xinput181 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__buf_4
Xinput192 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _3660_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_64_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _4981_/CLK _4981_/D vssd1 vssd1 vccd1 vccd1 _4981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _3932_/A0 _5089_/Q _3999_/S vssd1 vssd1 vccd1 vccd1 _3932_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3863_ _5730_/Q _3857_/Y _3862_/X _3887_/B _3925_/B1 vssd1 vssd1 vccd1 vccd1 _3863_/X
+ sky130_fd_sc_hd__a221o_1
X_2814_ _2850_/A1 _5426_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5426_/D sky130_fd_sc_hd__mux2_1
X_5602_ _5602_/CLK _5602_/D vssd1 vssd1 vccd1 vccd1 _5602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5533_ _5533_/CLK _5533_/D vssd1 vssd1 vccd1 vccd1 _5533_/Q sky130_fd_sc_hd__dfxtp_1
X_3794_ hold137/X _5245_/Q _3796_/A3 _3795_/B1 _4994_/Q vssd1 vssd1 vccd1 vccd1 _3794_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2745_ _3567_/A1 _5484_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5484_/D sky130_fd_sc_hd__mux2_1
X_2676_ _3600_/A1 _5573_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5573_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _5464_/CLK _5464_/D vssd1 vssd1 vccd1 vccd1 _5464_/Q sky130_fd_sc_hd__dfxtp_1
X_5395_ _5395_/CLK _5395_/D vssd1 vssd1 vccd1 vccd1 _5395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4415_ _4350_/A split5/A _4415_/A3 hold453/X vssd1 vssd1 vccd1 vccd1 _4415_/X sky130_fd_sc_hd__a31o_1
X_4346_ _5690_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4346_/X sky130_fd_sc_hd__or2_1
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4277_ _4277_/A _4277_/B _4277_/C _4276_/X vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__or4b_2
X_3228_ _2464_/A _5304_/Q _5053_/Q _3128_/B _3326_/C1 vssd1 vssd1 vccd1 vccd1 _3228_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3159_ _3159_/A _3159_/B vssd1 vssd1 vccd1 vccd1 _3159_/X sky130_fd_sc_hd__or2_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold391 hold398/X vssd1 vssd1 vccd1 vccd1 hold399/A sky130_fd_sc_hd__buf_2
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4763__348 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5454_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4804__389 _4821__406/A vssd1 vssd1 vccd1 vccd1 _5495_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4657__242 _4459__44/A vssd1 vssd1 vccd1 vccd1 _5343_/CLK sky130_fd_sc_hd__inv_2
X_2530_ _3393_/A0 _5711_/Q _2533_/S vssd1 vssd1 vccd1 vccd1 _5711_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2461_ _5334_/Q vssd1 vssd1 vccd1 vccd1 _3344_/A sky130_fd_sc_hd__inv_2
XFILLER_130_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _4204_/A _4200_/B vssd1 vssd1 vccd1 vccd1 _5546_/D sky130_fd_sc_hd__nor2_1
X_5180_ _5180_/CLK _5180_/D vssd1 vssd1 vccd1 vccd1 _5180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2709 hold2709/A vssd1 vssd1 vccd1 vccd1 hold929/A sky130_fd_sc_hd__buf_2
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4131_ _4122_/X _4123_/Y _4130_/Y _5750_/Q _4171_/A vssd1 vssd1 vccd1 vccd1 _4149_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4062_ _5667_/Q _5666_/Q _5665_/Q _5668_/Q vssd1 vssd1 vccd1 vccd1 _4063_/B sky130_fd_sc_hd__a31o_1
XFILLER_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3013_ _3003_/X _3004_/X _3075_/B1 _3001_/X vssd1 vssd1 vccd1 vccd1 _3013_/X sky130_fd_sc_hd__a211o_1
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3915_ _5081_/Q _3926_/A2 _3923_/B1 _3914_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5081_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3846_ _4399_/C _3888_/C vssd1 vssd1 vccd1 vccd1 _3887_/A sky130_fd_sc_hd__or2_4
X_3777_ _3824_/A1 _5113_/Q _3777_/A3 _3776_/X vssd1 vssd1 vccd1 vccd1 _3777_/X sky130_fd_sc_hd__a31o_4
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2728_ _3277_/A1 _5499_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5499_/D sky130_fd_sc_hd__mux2_1
X_5516_ _5516_/CLK _5516_/D vssd1 vssd1 vccd1 vccd1 _5516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5447_ _5447_/CLK _5447_/D vssd1 vssd1 vccd1 vccd1 _5447_/Q sky130_fd_sc_hd__dfxtp_1
X_2659_ _3602_/A1 _5587_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5587_/D sky130_fd_sc_hd__mux2_1
X_5378_ _5378_/CLK _5378_/D vssd1 vssd1 vccd1 vccd1 _5378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4329_ _4081_/B _4080_/B _4328_/X _4325_/B _4325_/A vssd1 vssd1 vccd1 vccd1 _4329_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3718_/A1 _3698_/X _3699_/X split4/X vssd1 vssd1 vccd1 vccd1 _3700_/X sky130_fd_sc_hd__o211a_1
XFILLER_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3631_ _4352_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3631_/X sky130_fd_sc_hd__or2_1
XFILLER_128_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3562_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3570_/S sky130_fd_sc_hd__nor2_8
XFILLER_127_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2513_ _2499_/X _2511_/Y _3782_/A vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__a21oi_4
X_5301_ _5301_/CLK _5301_/D vssd1 vssd1 vccd1 vccd1 _5301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4891__476 _4892__477/A vssd1 vssd1 vccd1 vccd1 _5612_/CLK sky130_fd_sc_hd__inv_2
X_3493_ _3592_/A1 _5167_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5167_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5232_ _5232_/CLK _5232_/D vssd1 vssd1 vccd1 vccd1 _5232_/Q sky130_fd_sc_hd__dfxtp_1
X_2444_ _5674_/Q vssd1 vssd1 vccd1 vccd1 _2444_/Y sky130_fd_sc_hd__inv_2
X_5163_ _5163_/CLK _5163_/D vssd1 vssd1 vccd1 vccd1 _5163_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2528 hold2528/A vssd1 vssd1 vccd1 vccd1 hold2528/X sky130_fd_sc_hd__buf_2
Xhold2517 hold2517/A vssd1 vssd1 vccd1 vccd1 _5323_/D sky130_fd_sc_hd__buf_2
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2539 hold2539/A vssd1 vssd1 vccd1 vccd1 hold848/A sky130_fd_sc_hd__buf_2
Xhold1816 hold2578/X vssd1 vssd1 vccd1 vccd1 hold2579/A sky130_fd_sc_hd__buf_2
Xhold1827 hold1827/A vssd1 vssd1 vccd1 vccd1 _5735_/D sky130_fd_sc_hd__buf_2
X_4114_ _5745_/Q _4114_/B _4114_/C vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__nand3b_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1849 hold787/X vssd1 vssd1 vccd1 vccd1 hold1849/X sky130_fd_sc_hd__buf_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1838 hold151/X vssd1 vssd1 vccd1 vccd1 hold1838/X sky130_fd_sc_hd__buf_2
X_5094_ _5542_/CLK _5094_/D vssd1 vssd1 vccd1 vccd1 _5094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4045_ _4046_/B _4046_/C _5749_/Q vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__a21bo_1
X_4785__370 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5476_/CLK sky130_fd_sc_hd__inv_2
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3829_ _3829_/A _3829_/B _3829_/C vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__and3_1
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput271 _3628_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__clkbuf_2
Xoutput260 _3660_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput282 _5854_/X vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_12
Xoutput293 _5864_/X vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_12
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4769__354 _4786__371/A vssd1 vssd1 vccd1 vccd1 _5460_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5850_ _5850_/A vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2993_ _5036_/Q _5533_/Q _3072_/S vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3614_ _4968_/Q _3614_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4968_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3545_ _5121_/Q _3608_/A1 _3552_/S vssd1 vssd1 vccd1 vccd1 _5121_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3476_ _3611_/A1 _5182_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5182_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold957 hold957/A vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__buf_2
Xhold968 hold968/A vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__buf_2
Xhold979 hold979/A vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__buf_2
XFILLER_143_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5215_ _5215_/CLK _5215_/D vssd1 vssd1 vccd1 vccd1 _5215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2303 _4355_/X vssd1 vssd1 vccd1 vccd1 hold2303/X sky130_fd_sc_hd__buf_2
XFILLER_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2325 hold2325/A vssd1 vssd1 vccd1 vccd1 hold991/A sky130_fd_sc_hd__buf_2
X_5146_ _5146_/CLK _5146_/D vssd1 vssd1 vccd1 vccd1 _5146_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1602 hold43/X vssd1 vssd1 vccd1 vccd1 hold1602/X sky130_fd_sc_hd__buf_2
XFILLER_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1624 hold2188/X vssd1 vssd1 vccd1 vccd1 hold2189/A sky130_fd_sc_hd__buf_2
Xhold2358 hold2358/A vssd1 vssd1 vccd1 vccd1 hold2358/X sky130_fd_sc_hd__buf_2
Xhold2369 hold754/X vssd1 vssd1 vccd1 vccd1 hold2369/X sky130_fd_sc_hd__buf_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1613 hold1613/A vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__buf_2
X_5077_ _5383_/CLK _5077_/D vssd1 vssd1 vccd1 vccd1 _5077_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1646 hold2594/X vssd1 vssd1 vccd1 vccd1 hold2595/A sky130_fd_sc_hd__buf_2
Xhold1657 hold2303/X vssd1 vssd1 vccd1 vccd1 hold2304/A sky130_fd_sc_hd__buf_2
Xhold1668 hold2320/X vssd1 vssd1 vccd1 vccd1 hold2321/A sky130_fd_sc_hd__buf_2
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4028_ _5743_/Q _4266_/B vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__xor2_2
XFILLER_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4562__147 _4506__91/A vssd1 vssd1 vccd1 vccd1 _5212_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4603__188 _4456__41/A vssd1 vssd1 vccd1 vccd1 _5277_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold209 hold401/X vssd1 vssd1 vccd1 vccd1 hold402/A sky130_fd_sc_hd__buf_2
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3330_ _5441_/Q _5457_/Q _3330_/S vssd1 vssd1 vccd1 vccd1 _3330_/X sky130_fd_sc_hd__mux2_2
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5739_/CLK _5000_/D vssd1 vssd1 vccd1 vccd1 _5000_/Q sky130_fd_sc_hd__dfxtp_1
X_3261_ _3357_/B _3259_/X _3260_/X _3323_/C1 vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__o211a_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4504__89 _4504__89/A vssd1 vssd1 vccd1 vccd1 _5146_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3192_ _5055_/Q _5279_/Q _5526_/Q _5306_/Q _3312_/S _3127_/A vssd1 vssd1 vccd1 vccd1
+ _3192_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5902_ _5902_/A vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2976_ _3034_/A _2974_/X _2975_/X _3097_/B vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__o211a_1
X_4897__482 _4897__482/A vssd1 vssd1 vccd1 vccd1 _5618_/CLK sky130_fd_sc_hd__inv_2
X_5695_ _5697_/CLK _5695_/D vssd1 vssd1 vccd1 vccd1 _5695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold710 hold710/A vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__buf_2
Xhold732 _3832_/X vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__buf_2
Xhold754 hold754/A vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__buf_2
X_3528_ _5136_/Q _3609_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5136_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold787 hold787/A vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__buf_2
X_3459_ _3612_/A1 _5197_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5197_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2111 hold474/X vssd1 vssd1 vccd1 vccd1 hold2111/X sky130_fd_sc_hd__buf_2
XFILLER_130_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2144 hold2144/A vssd1 vssd1 vccd1 vccd1 hold541/A sky130_fd_sc_hd__buf_2
X_5129_ _5129_/CLK _5129_/D vssd1 vssd1 vccd1 vccd1 _5129_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2166 hold2166/A vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__buf_2
Xhold2155 hold2155/A vssd1 vssd1 vccd1 vccd1 _3860_/B1 sky130_fd_sc_hd__buf_2
Xhold2188 hold2188/A vssd1 vssd1 vccd1 vccd1 hold2188/X sky130_fd_sc_hd__buf_2
Xhold1443 hold2109/X vssd1 vssd1 vccd1 vccd1 hold2110/A sky130_fd_sc_hd__buf_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1476 hold2245/X vssd1 vssd1 vccd1 vccd1 hold2246/A sky130_fd_sc_hd__buf_2
Xhold1465 hold2236/X vssd1 vssd1 vccd1 vccd1 hold2237/A sky130_fd_sc_hd__buf_2
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1498 hold26/X vssd1 vssd1 vccd1 vccd1 hold972/A sky130_fd_sc_hd__buf_2
Xhold1487 hold966/X vssd1 vssd1 vccd1 vccd1 _5092_/D sky130_fd_sc_hd__buf_2
XFILLER_26_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_67_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5691_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4690__275 _5384_/CLK vssd1 vssd1 vccd1 vccd1 _5379_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xsplit4 split4/A vssd1 vssd1 vccd1 vccd1 split4/X sky130_fd_sc_hd__buf_2
XFILLER_0_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__buf_2
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__buf_2
XFILLER_36_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold70 hold99/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__buf_2
XFILLER_91_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2830_ _3393_/A0 _5412_/Q _2833_/S vssd1 vssd1 vccd1 vccd1 _5412_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2761_ _3391_/A0 _5470_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5470_/D sky130_fd_sc_hd__mux2_1
X_2692_ _3597_/A1 _5531_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5531_/D sky130_fd_sc_hd__mux2_1
X_5480_ _5480_/CLK _5480_/D vssd1 vssd1 vccd1 vccd1 _5480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _2892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931__516 _4454__39/A vssd1 vssd1 vccd1 vccd1 _5652_/CLK sky130_fd_sc_hd__inv_2
X_4362_ _5336_/Q _4368_/A vssd1 vssd1 vccd1 vccd1 _5728_/D sky130_fd_sc_hd__and2_1
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout519 _5365_/Q vssd1 vssd1 vccd1 vccd1 _2942_/S1 sky130_fd_sc_hd__buf_4
X_4293_ _4292_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5666_/D sky130_fd_sc_hd__and2b_1
Xfanout508 _2490_/X vssd1 vssd1 vccd1 vccd1 _3926_/A2 sky130_fd_sc_hd__buf_6
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _5505_/Q _2464_/A _3128_/B _5497_/Q _3316_/C1 vssd1 vssd1 vccd1 vccd1 _3313_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3241_/X _3243_/X _3357_/A vssd1 vssd1 vccd1 vccd1 _3244_/X sky130_fd_sc_hd__o21a_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3175_ _5503_/Q _5495_/Q _5487_/Q _5511_/Q _3327_/S _3219_/S0 vssd1 vssd1 vccd1 vccd1
+ _3175_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4825__410 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5516_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2959_ _5165_/Q _5350_/Q _3005_/S vssd1 vssd1 vccd1 vccd1 _2959_/X sky130_fd_sc_hd__mux2_1
X_5747_ _5747_/CLK _5747_/D vssd1 vssd1 vccd1 vccd1 _5747_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5678_ _5738_/CLK _5678_/D vssd1 vssd1 vccd1 vccd1 _5678_/Q sky130_fd_sc_hd__dfxtp_4
X_4674__259 _4485__70/A vssd1 vssd1 vccd1 vccd1 _5362_/CLK sky130_fd_sc_hd__inv_2
Xhold551 hold576/X vssd1 vssd1 vccd1 vccd1 hold577/A sky130_fd_sc_hd__buf_2
XFILLER_2_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold584 hold584/A vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__buf_2
Xhold595 hold740/X vssd1 vssd1 vccd1 vccd1 hold741/A sky130_fd_sc_hd__buf_2
Xhold573 _4241_/X vssd1 vssd1 vccd1 vccd1 _5564_/D sky130_fd_sc_hd__buf_2
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1240 hold1950/X vssd1 vssd1 vccd1 vccd1 hold1951/A sky130_fd_sc_hd__buf_2
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_114_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5246_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1262 hold2489/X vssd1 vssd1 vccd1 vccd1 hold2490/A sky130_fd_sc_hd__buf_2
X_4568__153 _4432__17/A vssd1 vssd1 vccd1 vccd1 _5218_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4609__194 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5283_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2471__1 _4419__4/A vssd1 vssd1 vccd1 vccd1 _4967_/CLK sky130_fd_sc_hd__inv_2
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput160 input160/A vssd1 vssd1 vccd1 vccd1 _3664_/A sky130_fd_sc_hd__buf_4
Xinput171 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__buf_4
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput193 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__buf_6
Xinput182 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__buf_4
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _4980_/CLK _4980_/D vssd1 vssd1 vccd1 vccd1 _4980_/Q sky130_fd_sc_hd__dfxtp_1
X_3931_ _3931_/A _3931_/B _3931_/C split1/A vssd1 vssd1 vccd1 vccd1 _3931_/X sky130_fd_sc_hd__or4b_2
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3862_ _3998_/A1 _5203_/Q _3882_/A3 _3855_/X vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__a31o_1
X_2813_ _2849_/A1 _5427_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5427_/D sky130_fd_sc_hd__mux2_1
X_5601_ _5601_/CLK _5601_/D vssd1 vssd1 vccd1 vccd1 _5601_/Q sky130_fd_sc_hd__dfxtp_1
X_5532_ _5532_/CLK _5532_/D vssd1 vssd1 vccd1 vccd1 _5532_/Q sky130_fd_sc_hd__dfxtp_1
X_3793_ hold137/X _5244_/Q _3796_/A3 _3796_/B1 _4993_/Q vssd1 vssd1 vccd1 vccd1 _3793_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2744_ _3218_/A1 _5485_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5485_/D sky130_fd_sc_hd__mux2_1
X_2675_ _3599_/A1 _5574_/Q _2682_/S vssd1 vssd1 vccd1 vccd1 _5574_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5463_ _5463_/CLK _5463_/D vssd1 vssd1 vccd1 vccd1 _5463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5394_ _5394_/CLK _5394_/D vssd1 vssd1 vccd1 vccd1 _5394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4414_ _5754_/Q _4401_/Y _4414_/B1 vssd1 vssd1 vccd1 vccd1 _4414_/X sky130_fd_sc_hd__a21o_1
X_4345_ _5690_/Q _4324_/X _4344_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _5689_/D sky130_fd_sc_hd__o211a_1
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4276_ _4070_/Y _4071_/X _4275_/X _4031_/X vssd1 vssd1 vccd1 vccd1 _4276_/X sky130_fd_sc_hd__o211a_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3227_ _5524_/Q _5277_/Q _3324_/S vssd1 vssd1 vccd1 vccd1 _3227_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3158_ _5344_/Q _3125_/A _3353_/A _3155_/X vssd1 vssd1 vccd1 vccd1 _3158_/X sky130_fd_sc_hd__a22o_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3089_ _3089_/A _3089_/B vssd1 vssd1 vccd1 vccd1 _5371_/D sky130_fd_sc_hd__nor2_1
XFILLER_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold392 hold400/X vssd1 vssd1 vccd1 vccd1 hold401/A sky130_fd_sc_hd__buf_2
XFILLER_78_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1092 hold2317/X vssd1 vssd1 vccd1 vccd1 hold2318/A sky130_fd_sc_hd__buf_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_wb_clk_i _5743_/CLK vssd1 vssd1 vccd1 vccd1 _5747_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4696__281 _5543_/CLK vssd1 vssd1 vccd1 vccd1 _5387_/CLK sky130_fd_sc_hd__inv_2
X_2460_ _2460_/A vssd1 vssd1 vccd1 vccd1 _2460_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _4130_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _4130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4061_ _4059_/X _4060_/Y _4055_/X _4056_/X vssd1 vssd1 vccd1 vccd1 _4271_/C sky130_fd_sc_hd__o211a_1
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3012_ _3043_/A _3012_/B _3012_/C vssd1 vssd1 vccd1 vccd1 _3012_/X sky130_fd_sc_hd__or3_1
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3914_ _5740_/Q _3924_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3914_/X sky130_fd_sc_hd__and3_1
XFILLER_60_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3845_ _4399_/C _3888_/C vssd1 vssd1 vccd1 vccd1 _3845_/Y sky130_fd_sc_hd__nor2_1
X_4937__522 _4937__522/A vssd1 vssd1 vccd1 vccd1 _5658_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3776_ input35/X input2/X _3638_/B _3775_/X split1/A vssd1 vssd1 vccd1 vccd1 _3776_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_145_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2727_ _3567_/A1 _5500_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5500_/D sky130_fd_sc_hd__mux2_1
X_5515_ _5515_/CLK _5515_/D vssd1 vssd1 vccd1 vccd1 _5515_/Q sky130_fd_sc_hd__dfxtp_1
X_5446_ _5446_/CLK _5446_/D vssd1 vssd1 vccd1 vccd1 _5446_/Q sky130_fd_sc_hd__dfxtp_1
X_2658_ _3601_/A1 _5588_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5588_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5377_ _5377_/CLK _5377_/D vssd1 vssd1 vccd1 vccd1 _5377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2589_ _3391_/A0 _5628_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5628_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4328_ _5682_/Q _5681_/Q vssd1 vssd1 vccd1 vccd1 _4328_/X sky130_fd_sc_hd__or2_1
X_4259_ _5752_/Q _4259_/B _4259_/C vssd1 vssd1 vccd1 vccd1 _4260_/D sky130_fd_sc_hd__and3b_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730__315 _4731__316/A vssd1 vssd1 vccd1 vccd1 _5421_/CLK sky130_fd_sc_hd__inv_2
XFILLER_144_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3630_ _4351_/B _3638_/B vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__or2_1
XFILLER_128_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3561_ _5058_/Q _3606_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5058_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2512_ _3930_/C _2512_/B _2512_/C _2512_/D vssd1 vssd1 vccd1 vccd1 _4369_/C sky130_fd_sc_hd__or4_1
X_5300_ _5300_/CLK _5300_/D vssd1 vssd1 vccd1 vccd1 _5300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3492_ _3591_/A1 _5168_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5168_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5231_ _5231_/CLK _5231_/D vssd1 vssd1 vccd1 vccd1 _5231_/Q sky130_fd_sc_hd__dfxtp_1
X_2443_ _5675_/Q vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5162_ _5162_/CLK _5162_/D vssd1 vssd1 vccd1 vccd1 _5162_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2529 hold2529/A vssd1 vssd1 vccd1 vccd1 hold2529/X sky130_fd_sc_hd__buf_2
X_4113_ _4114_/B _4114_/C _5745_/Q vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__a21bo_1
X_5093_ _5542_/CLK _5093_/D vssd1 vssd1 vccd1 vccd1 _5093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1839 hold1839/A vssd1 vssd1 vccd1 vccd1 _5023_/D sky130_fd_sc_hd__buf_2
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _4046_/B _4046_/C vssd1 vssd1 vccd1 vccd1 _4253_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3828_ _3830_/B _3828_/B _3829_/C vssd1 vssd1 vccd1 vccd1 _3828_/X sky130_fd_sc_hd__and3_1
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3759_ _3759_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3759_/X sky130_fd_sc_hd__and2_1
XFILLER_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput250 _3651_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput261 _3632_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5429_ _5429_/CLK _5429_/D vssd1 vssd1 vccd1 vccd1 _5429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput272 _3623_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__clkbuf_2
XFILLER_58_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput294 _5865_/X vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_12
Xoutput283 _5855_/X vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_12
XFILLER_102_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2992_ _5116_/Q _3041_/A2 _2945_/A _2991_/X vssd1 vssd1 vccd1 vccd1 _3012_/C sky130_fd_sc_hd__o211a_1
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3613_ _4969_/Q _3613_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4969_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold903 hold903/A vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__buf_2
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3544_ _3589_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3552_/S sky130_fd_sc_hd__nor2_8
X_3475_ _3610_/A1 _5183_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5183_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold969 hold969/A vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__buf_2
Xhold958 hold958/A vssd1 vssd1 vccd1 vccd1 hold958/X sky130_fd_sc_hd__buf_2
XFILLER_142_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _5214_/CLK _5214_/D vssd1 vssd1 vccd1 vccd1 _5214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2304 hold2304/A vssd1 vssd1 vccd1 vccd1 hold2304/X sky130_fd_sc_hd__buf_2
Xhold2326 hold991/X vssd1 vssd1 vccd1 vccd1 hold2326/X sky130_fd_sc_hd__buf_2
X_5145_ _5145_/CLK _5145_/D vssd1 vssd1 vccd1 vccd1 _5145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1603 hold1603/A vssd1 vssd1 vccd1 vccd1 _3944_/A0 sky130_fd_sc_hd__buf_2
Xhold1614 hold49/X vssd1 vssd1 vccd1 vccd1 hold1614/X sky130_fd_sc_hd__buf_2
Xhold2359 hold2359/A vssd1 vssd1 vccd1 vccd1 _5694_/D sky130_fd_sc_hd__buf_2
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5076_ _5725_/CLK _5076_/D vssd1 vssd1 vccd1 vccd1 _5076_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1647 hold2596/X vssd1 vssd1 vccd1 vccd1 _4414_/B1 sky130_fd_sc_hd__buf_2
Xhold1658 hold2305/X vssd1 vssd1 vccd1 vccd1 hold2306/A sky130_fd_sc_hd__buf_2
XFILLER_38_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1669 hold2322/X vssd1 vssd1 vccd1 vccd1 hold2323/A sky130_fd_sc_hd__buf_2
X_4027_ _4027_/A _4027_/B vssd1 vssd1 vccd1 vccd1 _4266_/B sky130_fd_sc_hd__xnor2_4
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2893 hold2904/X vssd1 vssd1 vccd1 vccd1 hold2905/A sky130_fd_sc_hd__buf_2
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842__427 _4468__53/A vssd1 vssd1 vccd1 vccd1 _5535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4736__321 _4744__329/A vssd1 vssd1 vccd1 vccd1 _5427_/CLK sky130_fd_sc_hd__inv_2
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3260_ _5702_/Q _3331_/A2 _3326_/B2 _5718_/Q vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__o22a_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3316_/C1 _3188_/X _3190_/X vssd1 vssd1 vccd1 vccd1 _3191_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5901_ _5901_/A vssd1 vssd1 vccd1 vccd1 _5901_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ _5436_/Q _2460_/Y _3031_/B1 _5428_/Q vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5694_ _5734_/CLK _5694_/D vssd1 vssd1 vccd1 vccd1 _5694_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold711 hold711/A vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__buf_2
Xhold700 hold732/X vssd1 vssd1 vccd1 vccd1 hold733/A sky130_fd_sc_hd__buf_2
X_3527_ _5137_/Q _3590_/A1 _3534_/S vssd1 vssd1 vccd1 vccd1 _5137_/D sky130_fd_sc_hd__mux2_1
Xhold733 hold733/A vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__buf_2
XFILLER_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold766 hold766/A vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__buf_2
X_3458_ _3611_/A1 _5198_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5198_/D sky130_fd_sc_hd__mux2_1
Xhold799 hold799/A vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__buf_2
Xhold2112 hold2112/A vssd1 vssd1 vccd1 vccd1 _4984_/D sky130_fd_sc_hd__buf_2
XFILLER_39_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2134 _3874_/X vssd1 vssd1 vccd1 vccd1 hold2134/X sky130_fd_sc_hd__buf_2
Xhold2145 hold541/X vssd1 vssd1 vccd1 vccd1 hold2145/X sky130_fd_sc_hd__buf_2
X_3389_ _3389_/A0 _5289_/Q _3396_/S vssd1 vssd1 vccd1 vccd1 _5289_/D sky130_fd_sc_hd__mux2_4
XFILLER_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5128_ _5128_/CLK _5128_/D vssd1 vssd1 vccd1 vccd1 _5128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2167 _4095_/X vssd1 vssd1 vccd1 vccd1 hold2167/X sky130_fd_sc_hd__buf_2
Xhold2156 _3860_/X vssd1 vssd1 vccd1 vccd1 hold2156/X sky130_fd_sc_hd__buf_2
Xhold1433 hold2095/X vssd1 vssd1 vccd1 vccd1 hold2096/A sky130_fd_sc_hd__buf_2
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2189 hold2189/A vssd1 vssd1 vccd1 vccd1 _5726_/D sky130_fd_sc_hd__buf_2
Xhold1477 hold2247/X vssd1 vssd1 vccd1 vccd1 hold2248/A sky130_fd_sc_hd__buf_2
Xhold1466 hold2238/X vssd1 vssd1 vccd1 vccd1 hold2239/A sky130_fd_sc_hd__buf_2
Xhold1444 hold2111/X vssd1 vssd1 vccd1 vccd1 hold2112/A sky130_fd_sc_hd__buf_2
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1455 hold1459/X vssd1 vssd1 vccd1 vccd1 hold1455/X sky130_fd_sc_hd__buf_2
X_5059_ _5059_/CLK _5059_/D vssd1 vssd1 vccd1 vccd1 _5059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1499 hold972/X vssd1 vssd1 vccd1 vccd1 _5093_/D sky130_fd_sc_hd__buf_2
Xhold1488 hold2256/X vssd1 vssd1 vccd1 vccd1 hold2257/A sky130_fd_sc_hd__buf_2
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4882__467/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xsplit5 split5/A vssd1 vssd1 vccd1 vccd1 split5/X sky130_fd_sc_hd__clkbuf_2
Xhold2690 hold291/X vssd1 vssd1 vccd1 vccd1 hold2690/X sky130_fd_sc_hd__buf_2
Xhold82 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__buf_2
Xhold71 hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__buf_2
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__buf_2
XFILLER_91_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__buf_2
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2760_ _3390_/A0 _5471_/Q _2766_/S vssd1 vssd1 vccd1 vccd1 _5471_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2691_ _3605_/A1 _5532_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5532_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _3145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4361_ _4361_/A _4361_/B vssd1 vssd1 vccd1 vccd1 _4361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4292_ _4258_/B _4308_/A2 _4308_/B1 _2452_/Y vssd1 vssd1 vccd1 vccd1 _4292_/X sky130_fd_sc_hd__o22a_1
Xfanout509 _2490_/X vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__buf_4
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _5481_/Q _5489_/Q _3312_/S vssd1 vssd1 vccd1 vccd1 _3312_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3336_/A1 _3223_/X _3226_/X _3242_/X _3136_/X vssd1 vssd1 vccd1 vccd1 _3243_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3174_ _5629_/Q _5519_/Q _5288_/Q _5471_/Q _3219_/S0 _3299_/S vssd1 vssd1 vccd1 vccd1
+ _3174_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4905__490 _4905__490/A vssd1 vssd1 vccd1 vccd1 _5626_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2958_ _3041_/B1 _2956_/X _2957_/X vssd1 vssd1 vccd1 vccd1 _2981_/B sky130_fd_sc_hd__o21a_1
X_5746_ _5747_/CLK _5746_/D vssd1 vssd1 vccd1 vccd1 _5746_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5677_ _5677_/CLK _5677_/D vssd1 vssd1 vccd1 vccd1 _5677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2889_ _5129_/Q _5161_/Q _5317_/Q _5362_/Q _2942_/S1 _3072_/S vssd1 vssd1 vccd1 vccd1
+ _2889_/X sky130_fd_sc_hd__mux4_2
XFILLER_144_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold552 hold578/X vssd1 vssd1 vccd1 vccd1 hold579/A sky130_fd_sc_hd__buf_2
Xhold541 hold541/A vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__buf_2
XFILLER_131_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold585 hold585/A vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__buf_2
Xhold596 _4243_/X vssd1 vssd1 vccd1 vccd1 _5565_/D sky130_fd_sc_hd__buf_2
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1241 hold1952/X vssd1 vssd1 vccd1 vccd1 hold1953/A sky130_fd_sc_hd__buf_2
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4954__539 _4956__541/A vssd1 vssd1 vccd1 vccd1 _5712_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4848__433 _5106_/CLK vssd1 vssd1 vccd1 vccd1 _5569_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput161 input161/A vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__buf_4
Xinput172 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__clkbuf_8
Xinput150 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _2495_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput194 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__buf_6
Xinput183 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _3652_/A sky130_fd_sc_hd__buf_4
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _3930_/A split1/A _3930_/C vssd1 vssd1 vccd1 vccd1 _3930_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3861_ _5754_/Q _3998_/A1 _3882_/A3 _3887_/A vssd1 vssd1 vccd1 vccd1 _3861_/X sky130_fd_sc_hd__a31o_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5600_ _5600_/CLK _5600_/D vssd1 vssd1 vccd1 vccd1 _5600_/Q sky130_fd_sc_hd__dfxtp_1
X_2812_ _2848_/A1 _5428_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5428_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3792_ hold137/X _5243_/Q _3796_/A3 _3795_/B1 _4992_/Q vssd1 vssd1 vccd1 vccd1 _3792_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_20_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5531_ _5531_/CLK _5531_/D vssd1 vssd1 vccd1 vccd1 _5531_/Q sky130_fd_sc_hd__dfxtp_1
X_2743_ _2743_/A0 _5486_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5486_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2674_ _2779_/A _3508_/A vssd1 vssd1 vccd1 vccd1 _2682_/S sky130_fd_sc_hd__or2_4
X_5462_ _5462_/CLK _5462_/D vssd1 vssd1 vccd1 vccd1 _5462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5393_ _5393_/CLK _5393_/D vssd1 vssd1 vccd1 vccd1 _5393_/Q sky130_fd_sc_hd__dfxtp_1
X_4413_ _4351_/A _4351_/B split4/A _4415_/A3 hold453/X vssd1 vssd1 vccd1 vccd1 _4413_/X
+ sky130_fd_sc_hd__a41o_1
X_4344_ _5689_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4344_/X sky130_fd_sc_hd__or2_1
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4275_ _4042_/B _4275_/B _4275_/C vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__and3b_1
X_3226_ _3357_/B _3224_/X _3225_/X vssd1 vssd1 vccd1 vccd1 _3226_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4485__70 _4485__70/A vssd1 vssd1 vccd1 vccd1 _5127_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3157_ _5345_/Q _4360_/B vssd1 vssd1 vccd1 vccd1 _3159_/B sky130_fd_sc_hd__nand2_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3088_ _3453_/C _3091_/A _2778_/A vssd1 vssd1 vccd1 vccd1 _3089_/B sky130_fd_sc_hd__o21ai_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4641__226 _4921__506/A vssd1 vssd1 vccd1 vccd1 _5327_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5729_ _5730_/CLK _5729_/D vssd1 vssd1 vccd1 vccd1 _5729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold371 _3782_/X vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__buf_2
XFILLER_2_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4535__120 _4478__63/A vssd1 vssd1 vccd1 vccd1 _5177_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold393 hold402/X vssd1 vssd1 vccd1 vccd1 hold403/A sky130_fd_sc_hd__buf_2
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1060 hold1964/X vssd1 vssd1 vccd1 vccd1 hold1965/A sky130_fd_sc_hd__buf_2
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1093 hold2321/X vssd1 vssd1 vccd1 vccd1 hold2322/A sky130_fd_sc_hd__buf_2
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4469__54/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4060_ _4259_/B _4259_/C _5753_/Q vssd1 vssd1 vccd1 vccd1 _4060_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3011_ _3008_/X _3010_/X _2919_/B _3007_/X vssd1 vssd1 vccd1 vccd1 _3011_/X sky130_fd_sc_hd__a211o_1
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3913_ _5080_/Q _2490_/X _3923_/B1 _3912_/X _3921_/C1 vssd1 vssd1 vccd1 vccd1 _5080_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3844_ _3844_/A _3955_/A _4399_/D vssd1 vssd1 vccd1 vccd1 _3888_/C sky130_fd_sc_hd__or3_4
XFILLER_60_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3775_ _5088_/Q _3931_/B vssd1 vssd1 vccd1 vccd1 _3775_/X sky130_fd_sc_hd__or2_1
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2726_ _3218_/A1 _5501_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5501_/D sky130_fd_sc_hd__mux2_1
X_5514_ _5514_/CLK _5514_/D vssd1 vssd1 vccd1 vccd1 _5514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2657_ _3600_/A1 _5589_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5589_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4519__104 _5262_/CLK vssd1 vssd1 vccd1 vccd1 _5161_/CLK sky130_fd_sc_hd__inv_2
X_5445_ _5445_/CLK _5445_/D vssd1 vssd1 vccd1 vccd1 _5445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5376_ _5376_/CLK _5376_/D vssd1 vssd1 vccd1 vccd1 _5376_/Q sky130_fd_sc_hd__dfxtp_1
X_2588_ _3390_/A0 _5629_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5629_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4327_ _5681_/Q _4325_/Y _4326_/X _4319_/B vssd1 vssd1 vccd1 vccd1 _5681_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4258_ _5753_/Q _4258_/B vssd1 vssd1 vccd1 vccd1 _4260_/C sky130_fd_sc_hd__xnor2_1
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3209_ _5501_/Q _5493_/Q _5485_/Q _5509_/Q _3281_/S _3130_/B vssd1 vssd1 vccd1 vccd1
+ _3209_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4189_ _5541_/Q _4187_/B1 _4210_/C _4141_/Y vssd1 vssd1 vccd1 vccd1 _4190_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold190 hold298/X vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__buf_2
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4810__395 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5501_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3560_ _5059_/Q _3605_/A1 _3561_/S vssd1 vssd1 vccd1 vccd1 _5059_/D sky130_fd_sc_hd__mux2_1
X_2511_ _3888_/A _4399_/C _3852_/A vssd1 vssd1 vccd1 vccd1 _2511_/Y sky130_fd_sc_hd__nor3_2
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3491_ _3590_/A1 _5169_/Q _3498_/S vssd1 vssd1 vccd1 vccd1 _5169_/D sky130_fd_sc_hd__mux2_1
X_5230_ _5230_/CLK _5230_/D vssd1 vssd1 vccd1 vccd1 _5230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2442_ _5676_/Q vssd1 vssd1 vccd1 vccd1 _2442_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5161_ _5161_/CLK _5161_/D vssd1 vssd1 vccd1 vccd1 _5161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1807 hold2536/X vssd1 vssd1 vccd1 vccd1 hold2537/A sky130_fd_sc_hd__buf_2
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4112_ _4114_/B _4114_/C vssd1 vssd1 vccd1 vccd1 _4112_/Y sky130_fd_sc_hd__nand2_1
X_5092_ _5751_/CLK _5092_/D vssd1 vssd1 vccd1 vccd1 _5092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4043_ _4065_/B _4008_/B _5671_/Q vssd1 vssd1 vccd1 vccd1 _4046_/C sky130_fd_sc_hd__a21o_1
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4455__40 _4455__40/A vssd1 vssd1 vccd1 vccd1 _5049_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3827_ _5024_/Q _5023_/Q _3827_/C vssd1 vssd1 vccd1 vccd1 _3827_/X sky130_fd_sc_hd__or3_1
X_3758_ _5006_/Q _3750_/B _3774_/B1 _3757_/X _3774_/C1 vssd1 vssd1 vccd1 vccd1 _3758_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2709_ _3394_/A0 _5515_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5515_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3689_ _5066_/Q input3/X _3931_/B vssd1 vssd1 vccd1 vccd1 _3689_/X sky130_fd_sc_hd__mux2_4
X_4753__338 _4786__371/A vssd1 vssd1 vccd1 vccd1 _5444_/CLK sky130_fd_sc_hd__inv_2
Xoutput251 _3652_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__clkbuf_2
Xoutput240 _3642_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput262 _3633_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__clkbuf_2
X_5428_ _5428_/CLK _5428_/D vssd1 vssd1 vccd1 vccd1 _5428_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput273 _3624_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__clkbuf_2
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5359_ _5359_/CLK _5359_/D vssd1 vssd1 vccd1 vccd1 _5359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput295 _5866_/X vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_12
Xoutput284 _5856_/X vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_12
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4647__232 _5248_/CLK vssd1 vssd1 vccd1 vccd1 _5333_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ _5228_/Q _2870_/B _2990_/X _3041_/B1 vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__o22a_1
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3612_ _4970_/Q _3612_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4970_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3543_ _3543_/A0 _5122_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5122_/D sky130_fd_sc_hd__mux2_1
X_3474_ _3609_/A1 _5184_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5184_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold959 hold959/A vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__buf_2
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5213_ _5213_/CLK _5213_/D vssd1 vssd1 vccd1 vccd1 _5213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5144_ _5144_/CLK _5144_/D vssd1 vssd1 vccd1 vccd1 _5144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2316 _4353_/X vssd1 vssd1 vccd1 vccd1 hold2316/X sky130_fd_sc_hd__buf_2
Xhold2327 hold2327/A vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__buf_2
Xhold2305 hold2305/A vssd1 vssd1 vccd1 vccd1 hold2305/X sky130_fd_sc_hd__buf_2
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1604 _3944_/X vssd1 vssd1 vccd1 vccd1 hold1604/X sky130_fd_sc_hd__buf_2
Xhold1615 hold1615/A vssd1 vssd1 vccd1 vccd1 _3943_/A0 sky130_fd_sc_hd__buf_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5075_ _5747_/CLK _5075_/D vssd1 vssd1 vccd1 vccd1 _5075_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1648 _4414_/X vssd1 vssd1 vccd1 vccd1 hold1648/X sky130_fd_sc_hd__buf_2
Xhold1659 hold2307/X vssd1 vssd1 vccd1 vccd1 hold2308/A sky130_fd_sc_hd__buf_2
X_4026_ _4026_/A _4274_/A _4026_/C vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__or3_1
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_108_wb_clk_i _5743_/CLK vssd1 vssd1 vccd1 vccd1 _5551_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2850 _4085_/X vssd1 vssd1 vccd1 vccd1 hold2850/X sky130_fd_sc_hd__buf_2
XFILLER_48_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2883 _4351_/X vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__buf_2
Xhold2894 hold2908/X vssd1 vssd1 vccd1 vccd1 hold2900/A sky130_fd_sc_hd__buf_2
X_4881__466 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5602_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4775__360 _4937__522/A vssd1 vssd1 vccd1 vccd1 _5466_/CLK sky130_fd_sc_hd__inv_2
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3190_ _3320_/C1 _3189_/X _3336_/A1 vssd1 vssd1 vccd1 vccd1 _3190_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5900_/A vssd1 vssd1 vccd1 vccd1 _5900_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4425__10 _4425__10/A vssd1 vssd1 vccd1 vccd1 _4976_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2974_ _5396_/Q _5404_/Q _3069_/S vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5733_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5693_ _5734_/CLK _5693_/D vssd1 vssd1 vccd1 vccd1 _5693_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold701 hold734/X vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__buf_2
X_3526_ _3526_/A _3526_/B vssd1 vssd1 vccd1 vccd1 _3534_/S sky130_fd_sc_hd__nor2_8
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold734 hold734/A vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__buf_2
Xhold723 hold723/A vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__buf_2
X_3457_ _3610_/A1 _5199_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5199_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2102 _3783_/X vssd1 vssd1 vccd1 vccd1 hold2102/X sky130_fd_sc_hd__buf_2
Xhold2135 hold2135/A vssd1 vssd1 vccd1 vccd1 hold521/A sky130_fd_sc_hd__buf_2
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3388_ _3397_/A _3388_/B vssd1 vssd1 vccd1 vccd1 _3396_/S sky130_fd_sc_hd__or2_4
XFILLER_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5127_ _5127_/CLK _5127_/D vssd1 vssd1 vccd1 vccd1 _5127_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2168 hold2168/A vssd1 vssd1 vccd1 vccd1 hold954/A sky130_fd_sc_hd__buf_2
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2157 hold2157/A vssd1 vssd1 vccd1 vccd1 hold561/A sky130_fd_sc_hd__buf_2
Xhold2146 hold2146/A vssd1 vssd1 vccd1 vccd1 _3885_/B1 sky130_fd_sc_hd__buf_2
Xhold1423 hold2081/X vssd1 vssd1 vccd1 vccd1 hold2082/A sky130_fd_sc_hd__buf_2
Xhold1434 hold2097/X vssd1 vssd1 vccd1 vccd1 hold2098/A sky130_fd_sc_hd__buf_2
X_5058_ _5058_/CLK _5058_/D vssd1 vssd1 vccd1 vccd1 _5058_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1456 hold1456/A vssd1 vssd1 vccd1 vccd1 hold452/A sky130_fd_sc_hd__buf_2
Xhold1467 hold2240/X vssd1 vssd1 vccd1 vccd1 hold2241/A sky130_fd_sc_hd__buf_2
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4009_ _5672_/Q _5671_/Q _5670_/Q _5669_/Q vssd1 vssd1 vccd1 vccd1 _4029_/C sky130_fd_sc_hd__and4_4
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1489 hold2258/X vssd1 vssd1 vccd1 vccd1 hold2259/A sky130_fd_sc_hd__buf_2
Xhold1478 hold2249/X vssd1 vssd1 vccd1 vccd1 hold2250/A sky130_fd_sc_hd__buf_2
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4759__344 _4883__468/A vssd1 vssd1 vccd1 vccd1 _5450_/CLK sky130_fd_sc_hd__inv_2
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_76_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5564_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__buf_2
Xhold2680 hold2680/A vssd1 vssd1 vccd1 vccd1 hold2680/X sky130_fd_sc_hd__buf_2
Xhold2691 hold2691/A vssd1 vssd1 vccd1 vccd1 hold2691/X sky130_fd_sc_hd__buf_2
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__buf_2
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__buf_2
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__buf_2
XFILLER_91_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2690_ _3604_/A1 _5533_/Q _2692_/S vssd1 vssd1 vccd1 vccd1 _5533_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _3219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4360_ _4360_/A _4360_/B vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3311_ _3328_/A _3309_/X _3310_/X _3171_/A vssd1 vssd1 vccd1 vccd1 _3311_/X sky130_fd_sc_hd__o211a_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4291_ _2453_/Y _4308_/A2 _4290_/X vssd1 vssd1 vccd1 vccd1 _5665_/D sky130_fd_sc_hd__a21oi_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4552__137 _4882__467/A vssd1 vssd1 vccd1 vccd1 _5194_/CLK sky130_fd_sc_hd__inv_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3353_/B _3242_/B _3242_/C vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__or3_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3240_/S _3172_/X _3333_/C1 vssd1 vssd1 vccd1 vccd1 _3173_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2957_ _2867_/A _5133_/Q _3041_/A2 _5141_/Q _3064_/C1 vssd1 vssd1 vccd1 vccd1 _2957_/X
+ sky130_fd_sc_hd__o221a_1
X_5745_ _5747_/CLK _5745_/D vssd1 vssd1 vccd1 vccd1 _5745_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2888_ _3029_/B1 _2886_/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__a21o_1
X_5676_ _5738_/CLK _5676_/D vssd1 vssd1 vccd1 vccd1 _5676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold553 hold580/X vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__buf_2
Xhold542 hold542/A vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__buf_2
XFILLER_1_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3509_ _3590_/A1 _5153_/Q _3516_/S vssd1 vssd1 vccd1 vccd1 _5153_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 hold1954/X vssd1 vssd1 vccd1 vccd1 hold1955/A sky130_fd_sc_hd__buf_2
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1220 hold1886/X vssd1 vssd1 vccd1 vccd1 hold1887/A sky130_fd_sc_hd__buf_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1275 hold2524/X vssd1 vssd1 vccd1 vccd1 hold2525/A sky130_fd_sc_hd__buf_2
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput162 input162/A vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__buf_4
XFILLER_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput140 input140/A vssd1 vssd1 vccd1 vccd1 _3675_/A sky130_fd_sc_hd__buf_4
Xinput151 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _2495_/D sky130_fd_sc_hd__clkbuf_2
X_4887__472 _4901__486/A vssd1 vssd1 vccd1 vccd1 _5608_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput195 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__buf_6
Xinput173 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__clkbuf_8
Xinput184 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _3653_/A sky130_fd_sc_hd__buf_4
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _5066_/Q _3959_/A _3860_/B1 vssd1 vssd1 vccd1 vccd1 _3860_/X sky130_fd_sc_hd__a21o_1
X_2811_ _3584_/A0 _5429_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5429_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3791_ hold137/X _5242_/Q _3796_/A3 _3795_/B1 _4991_/Q vssd1 vssd1 vccd1 vccd1 _3791_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5530_ _5557_/CLK _5530_/D vssd1 vssd1 vccd1 vccd1 _5530_/Q sky130_fd_sc_hd__dfxtp_4
X_2742_ _2790_/A0 _5487_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5487_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5461_ _5461_/CLK _5461_/D vssd1 vssd1 vccd1 vccd1 _5461_/Q sky130_fd_sc_hd__dfxtp_1
X_2673_ _5369_/Q _2673_/B _5370_/Q vssd1 vssd1 vccd1 vccd1 _3508_/A sky130_fd_sc_hd__or3b_4
X_4412_ _5753_/Q _4401_/Y _4411_/X vssd1 vssd1 vccd1 vccd1 _4412_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5392_ _5392_/CLK _5392_/D vssd1 vssd1 vccd1 vccd1 _5392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4343_ _5689_/Q _4324_/X _4342_/X _4082_/A vssd1 vssd1 vccd1 vccd1 _5688_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4274_ _4274_/A _4274_/B _4273_/X vssd1 vssd1 vccd1 vccd1 _4277_/C sky130_fd_sc_hd__or3b_1
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3225_ _5618_/Q _2464_/A _3128_/B _5610_/Q _3316_/C1 vssd1 vssd1 vccd1 vccd1 _3225_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3156_ _5345_/Q _4360_/B vssd1 vssd1 vccd1 vccd1 _3156_/X sky130_fd_sc_hd__and2_4
X_3087_ _3087_/A _3087_/B vssd1 vssd1 vccd1 vccd1 _5372_/D sky130_fd_sc_hd__nor2_1
XFILLER_94_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680__265 _5383_/CLK vssd1 vssd1 vccd1 vccd1 _5369_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ _3989_/A _3989_/B vssd1 vssd1 vccd1 vccd1 _3989_/X sky130_fd_sc_hd__and2_4
XFILLER_139_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5728_ _5734_/CLK _5728_/D vssd1 vssd1 vccd1 vccd1 _5728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5659_ _5659_/CLK _5659_/D vssd1 vssd1 vccd1 vccd1 _5659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold394 hold404/X vssd1 vssd1 vccd1 vccd1 _3970_/B sky130_fd_sc_hd__buf_2
Xhold372 hold372/A vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__buf_2
Xhold383 hold383/A vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__buf_2
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1050 hold150/X vssd1 vssd1 vccd1 vccd1 _3829_/C sky130_fd_sc_hd__buf_2
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1061 hold1966/X vssd1 vssd1 vccd1 vccd1 hold1967/A sky130_fd_sc_hd__buf_2
Xhold1072 hold2740/X vssd1 vssd1 vccd1 vccd1 hold1831/A sky130_fd_sc_hd__buf_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4921__506 _4921__506/A vssd1 vssd1 vccd1 vccd1 _5642_/CLK sky130_fd_sc_hd__inv_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4815__400 _4819__404/A vssd1 vssd1 vccd1 vccd1 _5506_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_91_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4892__477/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_20_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4438__23/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3010_ _5028_/Q _3041_/A2 _3041_/B1 _3009_/X vssd1 vssd1 vccd1 vccd1 _3010_/X sky130_fd_sc_hd__o22a_1
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664__249 _4477__62/A vssd1 vssd1 vccd1 vccd1 _5352_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3912_ _5741_/Q _3924_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3912_/X sky130_fd_sc_hd__and3_1
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3843_ _5090_/Q _3850_/B _3850_/C vssd1 vssd1 vccd1 vccd1 _4399_/D sky130_fd_sc_hd__or3_2
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3774_ _5014_/Q _3774_/A2 _3774_/B1 _3773_/X _3774_/C1 vssd1 vssd1 vccd1 vccd1 _3774_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2725_ _2743_/A0 _5502_/Q _2730_/S vssd1 vssd1 vccd1 vccd1 _5502_/D sky130_fd_sc_hd__mux2_1
X_5513_ _5513_/CLK _5513_/D vssd1 vssd1 vccd1 vccd1 _5513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4558__143 _4421__6/A vssd1 vssd1 vccd1 vccd1 _5200_/CLK sky130_fd_sc_hd__inv_2
X_2656_ _3599_/A1 _5590_/Q _2663_/S vssd1 vssd1 vccd1 vccd1 _5590_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput400 _3706_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__clkbuf_2
X_5444_ _5444_/CLK _5444_/D vssd1 vssd1 vccd1 vccd1 _5444_/Q sky130_fd_sc_hd__dfxtp_1
X_5375_ _5375_/CLK _5375_/D vssd1 vssd1 vccd1 vccd1 _5375_/Q sky130_fd_sc_hd__dfxtp_1
X_2587_ _3389_/A0 _5630_/Q _2594_/S vssd1 vssd1 vccd1 vccd1 _5630_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4326_ _2438_/Y _5664_/Q _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__a211o_1
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4257_ _4259_/B _4259_/C _5752_/Q vssd1 vssd1 vccd1 vccd1 _4260_/B sky130_fd_sc_hd__a21boi_1
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4188_ _4217_/A _4188_/B vssd1 vssd1 vccd1 vccd1 _5540_/D sky130_fd_sc_hd__nor2_1
X_3208_ _5627_/Q _5517_/Q _5286_/Q _5469_/Q _3219_/S0 _3330_/S vssd1 vssd1 vccd1 vccd1
+ _3208_/X sky130_fd_sc_hd__mux4_2
XFILLER_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3139_ _3140_/A _3140_/B vssd1 vssd1 vccd1 vccd1 _3139_/Y sky130_fd_sc_hd__nor2_2
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__buf_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold191 _3824_/X vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__buf_2
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3490_ _3607_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3498_/S sky130_fd_sc_hd__or2_4
X_2510_ _5090_/Q _3850_/B _2510_/C vssd1 vssd1 vccd1 vccd1 _3852_/A sky130_fd_sc_hd__or3_4
X_2441_ _5677_/Q vssd1 vssd1 vccd1 vccd1 _4027_/A sky130_fd_sc_hd__inv_2
XFILLER_111_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ _5160_/CLK _5160_/D vssd1 vssd1 vccd1 vccd1 _5160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1808 hold2538/X vssd1 vssd1 vccd1 vccd1 hold2539/A sky130_fd_sc_hd__buf_2
X_4111_ _4108_/B _4119_/C _4108_/D _5549_/Q vssd1 vssd1 vccd1 vccd1 _4114_/C sky130_fd_sc_hd__a31o_1
X_5091_ _5697_/CLK _5091_/D vssd1 vssd1 vccd1 vccd1 _5091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4042_ _4042_/A _4042_/B _4041_/Y vssd1 vssd1 vccd1 vccd1 _4042_/X sky130_fd_sc_hd__or3b_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470__55 _4470__55/A vssd1 vssd1 vccd1 vccd1 _5064_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3826_ _5024_/Q _5023_/Q vssd1 vssd1 vccd1 vccd1 _3828_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ _3757_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3757_/X sky130_fd_sc_hd__and2_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2708_ _3393_/A0 _5516_/Q _2711_/S vssd1 vssd1 vccd1 vccd1 _5516_/D sky130_fd_sc_hd__mux2_1
X_3688_ _5261_/Q _3688_/B vssd1 vssd1 vccd1 vccd1 _3688_/X sky130_fd_sc_hd__and2_1
XFILLER_118_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4792__377 _4816__401/A vssd1 vssd1 vccd1 vccd1 _5483_/CLK sky130_fd_sc_hd__inv_2
Xoutput252 _3653_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput241 _3643_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput230 _3666_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__clkbuf_2
X_2639_ _5604_/Q _3601_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _5604_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5427_ _5427_/CLK _5427_/D vssd1 vssd1 vccd1 vccd1 _5427_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput263 _3634_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5358_ _5358_/CLK _5358_/D vssd1 vssd1 vccd1 vccd1 _5358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput285 _5838_/X vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_12
Xoutput274 _5837_/X vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_12
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4309_ _4308_/X _4309_/B vssd1 vssd1 vccd1 vccd1 _5674_/D sky130_fd_sc_hd__and2b_1
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput296 _5839_/X vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_12
XFILLER_101_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5289_ _5289_/CLK _5289_/D vssd1 vssd1 vccd1 vccd1 _5289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4686__271 _4693__278/A vssd1 vssd1 vccd1 vccd1 _5375_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout490 hold364/A vssd1 vssd1 vccd1 vccd1 _3795_/B1 sky130_fd_sc_hd__clkbuf_8
X_4927__512 _4451__36/A vssd1 vssd1 vccd1 vccd1 _5648_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2990_ _5164_/Q _5349_/Q _3040_/S vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3611_ _4971_/Q _3611_/A1 _3615_/S vssd1 vssd1 vccd1 vccd1 _4971_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3542_ _3605_/A1 _5123_/Q _3543_/S vssd1 vssd1 vccd1 vccd1 _5123_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3473_ _3608_/A1 _5185_/Q _3480_/S vssd1 vssd1 vccd1 vccd1 _5185_/D sky130_fd_sc_hd__mux2_1
X_5212_ _5212_/CLK _5212_/D vssd1 vssd1 vccd1 vccd1 _5212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5143_ _5143_/CLK _5143_/D vssd1 vssd1 vccd1 vccd1 _5143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2306 hold2306/A vssd1 vssd1 vccd1 vccd1 hold717/A sky130_fd_sc_hd__buf_2
Xhold2328 hold36/X vssd1 vssd1 vccd1 vccd1 hold2328/X sky130_fd_sc_hd__buf_2
Xhold2317 hold2317/A vssd1 vssd1 vccd1 vccd1 hold2317/X sky130_fd_sc_hd__buf_2
XFILLER_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1605 hold1605/A vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__buf_2
Xhold1616 _3943_/X vssd1 vssd1 vccd1 vccd1 hold1616/X sky130_fd_sc_hd__buf_2
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2339 _4354_/X vssd1 vssd1 vccd1 vccd1 hold2339/X sky130_fd_sc_hd__buf_2
X_5074_ _5291_/CLK _5074_/D vssd1 vssd1 vccd1 vccd1 _5074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1649 hold1649/A vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__buf_2
XFILLER_38_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4025_ _4026_/A _4026_/C vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__or2_1
XFILLER_80_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4720__305 _4941__526/A vssd1 vssd1 vccd1 vccd1 _5411_/CLK sky130_fd_sc_hd__inv_2
X_3809_ _5260_/Q hold358/X _3810_/A3 hold349/X _5009_/Q vssd1 vssd1 vccd1 vccd1 _3809_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2862 _4086_/X vssd1 vssd1 vccd1 vccd1 hold2862/X sky130_fd_sc_hd__buf_2
XFILLER_85_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2884 hold184/X vssd1 vssd1 vccd1 vccd1 hold2884/X sky130_fd_sc_hd__buf_2
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440__25 _4424__9/A vssd1 vssd1 vccd1 vccd1 _5034_/CLK sky130_fd_sc_hd__inv_2
X_2973_ _5029_/Q _3041_/A2 _3041_/B1 _2972_/X vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5692_ _5734_/CLK _5692_/D vssd1 vssd1 vccd1 vccd1 _5692_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 hold702/A vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__buf_2
X_3525_ _5138_/Q _3615_/A1 _3525_/S vssd1 vssd1 vccd1 vccd1 _5138_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3456_ _3609_/A1 _5200_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _5200_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2103 hold2103/A vssd1 vssd1 vccd1 vccd1 hold463/A sky130_fd_sc_hd__buf_2
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2125 _3864_/X vssd1 vssd1 vccd1 vccd1 hold2125/X sky130_fd_sc_hd__buf_2
Xhold2136 hold521/X vssd1 vssd1 vccd1 vccd1 hold2136/X sky130_fd_sc_hd__buf_2
X_3387_ _5293_/Q _3387_/A1 _3387_/S vssd1 vssd1 vccd1 vccd1 _5293_/D sky130_fd_sc_hd__mux2_1
X_5126_ _5126_/CLK _5126_/D vssd1 vssd1 vccd1 vccd1 _5126_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1402 hold2163/X vssd1 vssd1 vccd1 vccd1 hold2164/A sky130_fd_sc_hd__buf_2
XFILLER_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2147 _3885_/X vssd1 vssd1 vccd1 vccd1 hold2147/X sky130_fd_sc_hd__buf_2
Xhold1413 hold2707/X vssd1 vssd1 vccd1 vccd1 hold2708/A sky130_fd_sc_hd__buf_2
Xhold1424 hold2083/X vssd1 vssd1 vccd1 vccd1 hold2084/A sky130_fd_sc_hd__buf_2
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5057_ _5057_/CLK _5057_/D vssd1 vssd1 vccd1 vccd1 _5057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1468 hold2242/X vssd1 vssd1 vccd1 vccd1 hold2243/A sky130_fd_sc_hd__buf_2
X_4008_ _4065_/B _4008_/B vssd1 vssd1 vccd1 vccd1 _4254_/B sky130_fd_sc_hd__nand2_2
Xhold1479 hold2251/X vssd1 vssd1 vccd1 vccd1 hold2252/A sky130_fd_sc_hd__buf_2
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4798__383 _4897__482/A vssd1 vssd1 vccd1 vccd1 _5489_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__buf_2
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2670 _3790_/X vssd1 vssd1 vccd1 vccd1 hold2670/X sky130_fd_sc_hd__buf_2
Xhold2681 hold2681/A vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__buf_2
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__buf_2
Xhold62 hold82/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__buf_2
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__buf_2
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__buf_2
XFILLER_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__buf_2
XFILLER_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_wb_clk_i clkbuf_4_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5677_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _3778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3310_ _5465_/Q _3331_/A2 _3237_/B _5623_/Q vssd1 vssd1 vccd1 vccd1 _3310_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4290_ _5665_/Q _4308_/B1 _4309_/B vssd1 vssd1 vccd1 vccd1 _4290_/X sky130_fd_sc_hd__a21bo_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4591__176 _4438__23/A vssd1 vssd1 vccd1 vccd1 _5241_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3334_/A1 _3240_/X _3239_/X _3169_/B vssd1 vssd1 vccd1 vccd1 _3241_/X sky130_fd_sc_hd__o211a_1
XFILLER_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ _5415_/Q _5391_/Q _5661_/Q _5423_/Q _3327_/S _3184_/S1 vssd1 vssd1 vccd1 vccd1
+ _3172_/X sky130_fd_sc_hd__mux4_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2956_ _5213_/Q _5149_/Q _3063_/S vssd1 vssd1 vccd1 vccd1 _2956_/X sky130_fd_sc_hd__mux2_1
X_5744_ _5747_/CLK _5744_/D vssd1 vssd1 vccd1 vccd1 _5744_/Q sky130_fd_sc_hd__dfxtp_4
X_2887_ _3073_/C1 _2885_/X _3043_/A vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5675_ _5738_/CLK _5675_/D vssd1 vssd1 vccd1 vccd1 _5675_/Q sky130_fd_sc_hd__dfxtp_2
Xhold554 hold554/A vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__buf_2
Xhold521 hold521/A vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__buf_2
X_4832__417 _4456__41/A vssd1 vssd1 vccd1 vccd1 _5523_/CLK sky130_fd_sc_hd__inv_2
XFILLER_131_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3508_ _3508_/A _3526_/B vssd1 vssd1 vccd1 vccd1 _3516_/S sky130_fd_sc_hd__or2_4
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold576 hold599/X vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__buf_2
X_3439_ _5221_/Q _3594_/A1 _3442_/S vssd1 vssd1 vccd1 vccd1 _5221_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5256_/CLK _5109_/D vssd1 vssd1 vccd1 vccd1 _5109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1232 hold1937/X vssd1 vssd1 vccd1 vccd1 hold1938/A sky130_fd_sc_hd__buf_2
Xhold1221 hold1888/X vssd1 vssd1 vccd1 vccd1 hold1889/A sky130_fd_sc_hd__buf_2
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1254 hold2472/X vssd1 vssd1 vccd1 vccd1 hold2473/A sky130_fd_sc_hd__buf_2
Xhold1276 hold2528/X vssd1 vssd1 vccd1 vccd1 hold2529/A sky130_fd_sc_hd__buf_2
XFILLER_58_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1298 hold2584/X vssd1 vssd1 vccd1 vccd1 hold2585/A sky130_fd_sc_hd__buf_2
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4726__311 _4941__526/A vssd1 vssd1 vccd1 vccd1 _5417_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput130 probe_out[95] vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput163 input163/A vssd1 vssd1 vccd1 vccd1 _3667_/A sky130_fd_sc_hd__buf_4
Xinput141 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _3732_/B sky130_fd_sc_hd__buf_6
Xinput152 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _2495_/C sky130_fd_sc_hd__clkbuf_2
Xinput196 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__buf_6
Xinput174 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__clkbuf_8
Xinput185 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__buf_4
XFILLER_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2810_ _3601_/A1 _5430_/Q _2815_/S vssd1 vssd1 vccd1 vccd1 _5430_/D sky130_fd_sc_hd__mux2_1
X_3790_ hold137/X _5022_/Q _3829_/A _3796_/B1 _4990_/Q vssd1 vssd1 vccd1 vccd1 _3790_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_20_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2741_ _2853_/A1 _5488_/Q _2748_/S vssd1 vssd1 vccd1 vccd1 _5488_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5460_ _5460_/CLK _5460_/D vssd1 vssd1 vccd1 vccd1 _5460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4411_ _4352_/A split5/A _4415_/A3 hold453/X vssd1 vssd1 vccd1 vccd1 _4411_/X sky130_fd_sc_hd__a31o_1
X_2672_ _5575_/Q _3387_/A1 _2672_/S vssd1 vssd1 vccd1 vccd1 _5575_/D sky130_fd_sc_hd__mux2_1
X_5391_ _5391_/CLK _5391_/D vssd1 vssd1 vccd1 vccd1 _5391_/Q sky130_fd_sc_hd__dfxtp_1
X_4342_ _5688_/Q _4348_/B vssd1 vssd1 vccd1 vccd1 _4342_/X sky130_fd_sc_hd__or2_1
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4273_ _5743_/Q _4266_/B _4049_/Y _4050_/X _4041_/Y vssd1 vssd1 vccd1 vccd1 _4273_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3224_ _5578_/Q _5594_/Q _3318_/S vssd1 vssd1 vccd1 vccd1 _3224_/X sky130_fd_sc_hd__mux2_1
.ends

